magic
tech sky130A
magscale 1 2
timestamp 1731114203
<< viali >>
rect 7113 31977 7147 32011
rect 10149 31977 10183 32011
rect 17877 31977 17911 32011
rect 18797 31977 18831 32011
rect 31677 31977 31711 32011
rect 5641 31909 5675 31943
rect 8677 31909 8711 31943
rect 12541 31909 12575 31943
rect 14381 31909 14415 31943
rect 3065 31841 3099 31875
rect 3893 31841 3927 31875
rect 6653 31841 6687 31875
rect 6929 31841 6963 31875
rect 9689 31841 9723 31875
rect 9965 31841 9999 31875
rect 11805 31841 11839 31875
rect 15393 31841 15427 31875
rect 16405 31841 16439 31875
rect 17693 31841 17727 31875
rect 18981 31841 19015 31875
rect 20913 31841 20947 31875
rect 22569 31841 22603 31875
rect 24041 31841 24075 31875
rect 25513 31841 25547 31875
rect 25605 31841 25639 31875
rect 25697 31841 25731 31875
rect 26249 31841 26283 31875
rect 26525 31841 26559 31875
rect 28641 31841 28675 31875
rect 30113 31841 30147 31875
rect 30389 31841 30423 31875
rect 31861 31841 31895 31875
rect 4353 31773 4387 31807
rect 14105 31773 14139 31807
rect 16681 31773 16715 31807
rect 21373 31773 21407 31807
rect 24409 31773 24443 31807
rect 26985 31773 27019 31807
rect 29101 31773 29135 31807
rect 26065 31705 26099 31739
rect 3249 31637 3283 31671
rect 22385 31637 22419 31671
rect 25789 31637 25823 31671
rect 11713 31365 11747 31399
rect 27537 31365 27571 31399
rect 3249 31297 3283 31331
rect 11069 31297 11103 31331
rect 12357 31297 12391 31331
rect 13461 31297 13495 31331
rect 14565 31297 14599 31331
rect 26065 31297 26099 31331
rect 30113 31297 30147 31331
rect 4261 31229 4295 31263
rect 11345 31229 11379 31263
rect 13001 31229 13035 31263
rect 15393 31229 15427 31263
rect 16589 31229 16623 31263
rect 18061 31229 18095 31263
rect 21281 31229 21315 31263
rect 23489 31229 23523 31263
rect 23765 31229 23799 31263
rect 24133 31229 24167 31263
rect 24593 31229 24627 31263
rect 24869 31229 24903 31263
rect 25053 31229 25087 31263
rect 25237 31229 25271 31263
rect 25395 31229 25429 31263
rect 25697 31229 25731 31263
rect 26203 31229 26237 31263
rect 26341 31229 26375 31263
rect 26433 31229 26467 31263
rect 26525 31229 26559 31263
rect 26893 31229 26927 31263
rect 27445 31229 27479 31263
rect 27721 31229 27755 31263
rect 28181 31229 28215 31263
rect 29653 31229 29687 31263
rect 24291 31161 24325 31195
rect 24409 31161 24443 31195
rect 24501 31161 24535 31195
rect 24961 31161 24995 31195
rect 25513 31161 25547 31195
rect 25605 31161 25639 31195
rect 29377 31161 29411 31195
rect 10793 31093 10827 31127
rect 11253 31093 11287 31127
rect 11805 31093 11839 31127
rect 15117 31093 15151 31127
rect 15301 31093 15335 31127
rect 16037 31093 16071 31127
rect 17509 31093 17543 31127
rect 18521 31093 18555 31127
rect 21373 31093 21407 31127
rect 23581 31093 23615 31127
rect 23949 31093 23983 31127
rect 24777 31093 24811 31127
rect 25881 31093 25915 31127
rect 26709 31093 26743 31127
rect 24041 30889 24075 30923
rect 26433 30889 26467 30923
rect 28273 30889 28307 30923
rect 10885 30821 10919 30855
rect 12541 30821 12575 30855
rect 15945 30821 15979 30855
rect 26247 30821 26281 30855
rect 30205 30821 30239 30855
rect 31585 30821 31619 30855
rect 4445 30753 4479 30787
rect 4537 30753 4571 30787
rect 12633 30753 12667 30787
rect 12817 30753 12851 30787
rect 18613 30753 18647 30787
rect 19349 30753 19383 30787
rect 19487 30753 19521 30787
rect 23857 30753 23891 30787
rect 25145 30753 25179 30787
rect 25329 30753 25363 30787
rect 26065 30753 26099 30787
rect 28825 30753 28859 30787
rect 29009 30753 29043 30787
rect 30481 30753 30515 30787
rect 3249 30685 3283 30719
rect 4813 30685 4847 30719
rect 10609 30685 10643 30719
rect 12357 30685 12391 30719
rect 13277 30685 13311 30719
rect 13553 30685 13587 30719
rect 15669 30685 15703 30719
rect 18429 30685 18463 30719
rect 19625 30685 19659 30719
rect 20361 30685 20395 30719
rect 20637 30685 20671 30719
rect 22109 30685 22143 30719
rect 22937 30685 22971 30719
rect 26525 30685 26559 30719
rect 26801 30685 26835 30719
rect 15025 30617 15059 30651
rect 17417 30617 17451 30651
rect 18153 30617 18187 30651
rect 19073 30617 19107 30651
rect 25513 30617 25547 30651
rect 12909 30549 12943 30583
rect 15485 30549 15519 30583
rect 20269 30549 20303 30583
rect 22293 30549 22327 30583
rect 24593 30549 24627 30583
rect 28733 30549 28767 30583
rect 14657 30345 14691 30379
rect 16957 30345 16991 30379
rect 23489 30345 23523 30379
rect 25329 30345 25363 30379
rect 12357 30277 12391 30311
rect 16037 30277 16071 30311
rect 18981 30277 19015 30311
rect 20913 30277 20947 30311
rect 25421 30277 25455 30311
rect 26065 30277 26099 30311
rect 28549 30277 28583 30311
rect 28733 30277 28767 30311
rect 30941 30277 30975 30311
rect 3249 30209 3283 30243
rect 9689 30209 9723 30243
rect 10609 30209 10643 30243
rect 12817 30209 12851 30243
rect 14565 30209 14599 30243
rect 15209 30209 15243 30243
rect 16589 30209 16623 30243
rect 17509 30209 17543 30243
rect 21465 30209 21499 30243
rect 21741 30209 21775 30243
rect 23581 30209 23615 30243
rect 23857 30209 23891 30243
rect 27537 30209 27571 30243
rect 27813 30209 27847 30243
rect 4445 30141 4479 30175
rect 8217 30141 8251 30175
rect 15025 30141 15059 30175
rect 16405 30141 16439 30175
rect 16865 30141 16899 30175
rect 17233 30141 17267 30175
rect 19257 30141 19291 30175
rect 20269 30141 20303 30175
rect 20453 30141 20487 30175
rect 25605 30141 25639 30175
rect 25789 30141 25823 30175
rect 25881 30141 25915 30175
rect 27905 30141 27939 30175
rect 28641 30141 28675 30175
rect 29160 30141 29194 30175
rect 29929 30141 29963 30175
rect 30665 30141 30699 30175
rect 31033 30141 31067 30175
rect 31401 30141 31435 30175
rect 31861 30141 31895 30175
rect 10885 30073 10919 30107
rect 14289 30073 14323 30107
rect 16497 30073 16531 30107
rect 19165 30073 19199 30107
rect 19625 30073 19659 30107
rect 21281 30073 21315 30107
rect 22017 30073 22051 30107
rect 8309 30005 8343 30039
rect 9137 30005 9171 30039
rect 15117 30005 15151 30039
rect 19717 30005 19751 30039
rect 20545 30005 20579 30039
rect 21373 30005 21407 30039
rect 29101 30005 29135 30039
rect 29285 30005 29319 30039
rect 29377 30005 29411 30039
rect 30113 30005 30147 30039
rect 31309 30005 31343 30039
rect 31677 30005 31711 30039
rect 4537 29801 4571 29835
rect 9781 29801 9815 29835
rect 10333 29801 10367 29835
rect 11989 29801 12023 29835
rect 13001 29801 13035 29835
rect 13921 29801 13955 29835
rect 15577 29801 15611 29835
rect 17233 29801 17267 29835
rect 21189 29801 21223 29835
rect 22753 29801 22787 29835
rect 25145 29801 25179 29835
rect 25789 29801 25823 29835
rect 27629 29801 27663 29835
rect 28825 29801 28859 29835
rect 29009 29801 29043 29835
rect 30205 29801 30239 29835
rect 11437 29733 11471 29767
rect 16865 29733 16899 29767
rect 19717 29733 19751 29767
rect 23489 29733 23523 29767
rect 31677 29733 31711 29767
rect 3157 29665 3191 29699
rect 4721 29665 4755 29699
rect 12081 29665 12115 29699
rect 14657 29665 14691 29699
rect 14933 29665 14967 29699
rect 16405 29665 16439 29699
rect 17693 29665 17727 29699
rect 19257 29665 19291 29699
rect 19441 29665 19475 29699
rect 22661 29665 22695 29699
rect 23029 29665 23063 29699
rect 23213 29665 23247 29699
rect 23305 29665 23339 29699
rect 24409 29665 24443 29699
rect 24501 29665 24535 29699
rect 24593 29665 24627 29699
rect 24711 29665 24745 29699
rect 25237 29665 25271 29699
rect 25329 29665 25363 29699
rect 25605 29665 25639 29699
rect 25789 29665 25823 29699
rect 28950 29665 28984 29699
rect 29469 29665 29503 29699
rect 30297 29665 30331 29699
rect 30481 29665 30515 29699
rect 3525 29597 3559 29631
rect 8033 29597 8067 29631
rect 8309 29597 8343 29631
rect 10977 29597 11011 29631
rect 11529 29597 11563 29631
rect 11621 29597 11655 29631
rect 12449 29597 12483 29631
rect 14013 29597 14047 29631
rect 14105 29597 14139 29631
rect 14565 29597 14599 29631
rect 15025 29597 15059 29631
rect 15761 29597 15795 29631
rect 16589 29597 16623 29631
rect 16773 29597 16807 29631
rect 17417 29597 17451 29631
rect 17601 29597 17635 29631
rect 18889 29597 18923 29631
rect 24133 29597 24167 29631
rect 24225 29597 24259 29631
rect 24869 29597 24903 29631
rect 24961 29597 24995 29631
rect 25881 29597 25915 29631
rect 26157 29597 26191 29631
rect 27721 29597 27755 29631
rect 28365 29597 28399 29631
rect 11069 29529 11103 29563
rect 13553 29529 13587 29563
rect 18061 29529 18095 29563
rect 23305 29529 23339 29563
rect 5089 29461 5123 29495
rect 13461 29461 13495 29495
rect 14381 29461 14415 29495
rect 18337 29461 18371 29495
rect 19165 29461 19199 29495
rect 21557 29461 21591 29495
rect 25513 29461 25547 29495
rect 29377 29461 29411 29495
rect 30021 29461 30055 29495
rect 3525 29257 3559 29291
rect 8033 29257 8067 29291
rect 19717 29257 19751 29291
rect 22004 29257 22038 29291
rect 23581 29257 23615 29291
rect 26341 29257 26375 29291
rect 26893 29257 26927 29291
rect 28273 29257 28307 29291
rect 29180 29257 29214 29291
rect 30665 29257 30699 29291
rect 7757 29189 7791 29223
rect 19533 29189 19567 29223
rect 28365 29189 28399 29223
rect 5549 29121 5583 29155
rect 8585 29121 8619 29155
rect 9781 29121 9815 29155
rect 10885 29121 10919 29155
rect 11897 29121 11931 29155
rect 13185 29121 13219 29155
rect 15393 29121 15427 29155
rect 17325 29121 17359 29155
rect 18797 29121 18831 29155
rect 20269 29121 20303 29155
rect 21741 29121 21775 29155
rect 23489 29121 23523 29155
rect 24225 29121 24259 29155
rect 25237 29121 25271 29155
rect 27445 29121 27479 29155
rect 27905 29121 27939 29155
rect 5273 29053 5307 29087
rect 5641 29053 5675 29087
rect 7665 29053 7699 29087
rect 8401 29053 8435 29087
rect 8861 29053 8895 29087
rect 11805 29053 11839 29087
rect 12541 29053 12575 29087
rect 13369 29053 13403 29087
rect 14657 29053 14691 29087
rect 15945 29053 15979 29087
rect 16221 29053 16255 29087
rect 17049 29053 17083 29087
rect 24961 29053 24995 29087
rect 25053 29053 25087 29087
rect 26249 29053 26283 29087
rect 26617 29053 26651 29087
rect 26709 29053 26743 29087
rect 27813 29053 27847 29087
rect 27997 29053 28031 29087
rect 28089 29053 28123 29087
rect 28733 29053 28767 29087
rect 28917 29053 28951 29087
rect 30941 29053 30975 29087
rect 31677 29053 31711 29087
rect 4997 28985 5031 29019
rect 9505 28985 9539 29019
rect 11161 28985 11195 29019
rect 14013 28985 14047 29019
rect 16865 28985 16899 29019
rect 20085 28985 20119 29019
rect 24041 28985 24075 29019
rect 28549 28985 28583 29019
rect 31401 28985 31435 29019
rect 8493 28917 8527 28951
rect 14105 28917 14139 28951
rect 14841 28917 14875 28951
rect 15853 28917 15887 28951
rect 20177 28917 20211 28951
rect 23949 28917 23983 28951
rect 26065 28917 26099 28951
rect 30849 28917 30883 28951
rect 8033 28713 8067 28747
rect 12633 28713 12667 28747
rect 15761 28713 15795 28747
rect 22661 28713 22695 28747
rect 23581 28713 23615 28747
rect 24593 28713 24627 28747
rect 26985 28713 27019 28747
rect 28641 28713 28675 28747
rect 29009 28713 29043 28747
rect 31033 28713 31067 28747
rect 12817 28645 12851 28679
rect 14289 28645 14323 28679
rect 24409 28645 24443 28679
rect 27169 28645 27203 28679
rect 27353 28645 27387 28679
rect 28917 28645 28951 28679
rect 29193 28645 29227 28679
rect 31677 28645 31711 28679
rect 6469 28577 6503 28611
rect 10885 28577 10919 28611
rect 12909 28577 12943 28611
rect 16037 28577 16071 28611
rect 16313 28577 16347 28611
rect 22569 28577 22603 28611
rect 23673 28577 23707 28611
rect 23765 28577 23799 28611
rect 24501 28577 24535 28611
rect 24685 28577 24719 28611
rect 27629 28577 27663 28611
rect 27813 28577 27847 28611
rect 27905 28577 27939 28611
rect 28089 28577 28123 28611
rect 28825 28577 28859 28611
rect 31401 28577 31435 28611
rect 3985 28509 4019 28543
rect 4261 28509 4295 28543
rect 5733 28509 5767 28543
rect 7205 28509 7239 28543
rect 9505 28509 9539 28543
rect 9781 28509 9815 28543
rect 10241 28509 10275 28543
rect 10793 28509 10827 28543
rect 11161 28509 11195 28543
rect 14013 28509 14047 28543
rect 17141 28509 17175 28543
rect 19809 28509 19843 28543
rect 29285 28509 29319 28543
rect 29561 28509 29595 28543
rect 31309 28509 31343 28543
rect 31769 28509 31803 28543
rect 27537 28441 27571 28475
rect 31125 28441 31159 28475
rect 5825 28373 5859 28407
rect 7849 28373 7883 28407
rect 13921 28373 13955 28407
rect 15945 28373 15979 28407
rect 16221 28373 16255 28407
rect 16589 28373 16623 28407
rect 17785 28373 17819 28407
rect 20453 28373 20487 28407
rect 27169 28373 27203 28407
rect 27997 28373 28031 28407
rect 5273 28169 5307 28203
rect 5457 28169 5491 28203
rect 9321 28169 9355 28203
rect 10701 28169 10735 28203
rect 13093 28169 13127 28203
rect 15577 28169 15611 28203
rect 19441 28169 19475 28203
rect 23949 28169 23983 28203
rect 26525 28169 26559 28203
rect 29837 28169 29871 28203
rect 30849 28169 30883 28203
rect 31033 28169 31067 28203
rect 28273 28101 28307 28135
rect 29193 28101 29227 28135
rect 3893 28033 3927 28067
rect 4721 28033 4755 28067
rect 6009 28033 6043 28067
rect 11345 28033 11379 28067
rect 14105 28033 14139 28067
rect 15853 28033 15887 28067
rect 17693 28033 17727 28067
rect 24685 28033 24719 28067
rect 24777 28033 24811 28067
rect 26065 28033 26099 28067
rect 26249 28033 26283 28067
rect 27537 28033 27571 28067
rect 28733 28033 28767 28067
rect 30389 28033 30423 28067
rect 5825 27965 5859 27999
rect 5917 27965 5951 27999
rect 7297 27965 7331 27999
rect 9873 27965 9907 27999
rect 10425 27965 10459 27999
rect 10885 27965 10919 27999
rect 10977 27965 11011 27999
rect 11253 27965 11287 27999
rect 13369 27965 13403 27999
rect 13829 27965 13863 27999
rect 19717 27965 19751 27999
rect 23305 27965 23339 27999
rect 23563 27965 23597 27999
rect 23673 27965 23707 27999
rect 24041 27965 24075 27999
rect 24501 27965 24535 27999
rect 24593 27965 24627 27999
rect 25053 27965 25087 27999
rect 25605 27965 25639 27999
rect 26157 27965 26191 27999
rect 26709 27965 26743 27999
rect 26893 27965 26927 27999
rect 28089 27965 28123 27999
rect 28457 27965 28491 27999
rect 28549 27965 28583 27999
rect 28641 27965 28675 27999
rect 29561 27965 29595 27999
rect 31217 27965 31251 27999
rect 4445 27897 4479 27931
rect 4905 27897 4939 27931
rect 6469 27897 6503 27931
rect 7573 27897 7607 27931
rect 11069 27897 11103 27931
rect 11621 27897 11655 27931
rect 13277 27897 13311 27931
rect 16681 27897 16715 27931
rect 17969 27897 18003 27931
rect 19625 27897 19659 27931
rect 26433 27897 26467 27931
rect 27169 27897 27203 27931
rect 27353 27897 27387 27931
rect 29469 27897 29503 27931
rect 30665 27897 30699 27931
rect 4813 27829 4847 27863
rect 7205 27829 7239 27863
rect 9045 27829 9079 27863
rect 10333 27829 10367 27863
rect 13737 27829 13771 27863
rect 17049 27829 17083 27863
rect 22753 27829 22787 27863
rect 24225 27829 24259 27863
rect 24317 27829 24351 27863
rect 26341 27829 26375 27863
rect 26985 27829 27019 27863
rect 29009 27829 29043 27863
rect 29653 27829 29687 27863
rect 30205 27829 30239 27863
rect 30297 27829 30331 27863
rect 30865 27829 30899 27863
rect 31861 27829 31895 27863
rect 6469 27625 6503 27659
rect 11897 27625 11931 27659
rect 17877 27625 17911 27659
rect 25329 27625 25363 27659
rect 30757 27625 30791 27659
rect 30920 27625 30954 27659
rect 5089 27557 5123 27591
rect 6745 27557 6779 27591
rect 8861 27557 8895 27591
rect 12449 27557 12483 27591
rect 13921 27557 13955 27591
rect 14657 27557 14691 27591
rect 17601 27557 17635 27591
rect 23029 27557 23063 27591
rect 25605 27557 25639 27591
rect 31125 27557 31159 27591
rect 4445 27489 4479 27523
rect 5181 27489 5215 27523
rect 6653 27489 6687 27523
rect 6837 27489 6871 27523
rect 7021 27489 7055 27523
rect 9413 27489 9447 27523
rect 9781 27489 9815 27523
rect 10057 27489 10091 27523
rect 12173 27489 12207 27523
rect 14289 27489 14323 27523
rect 17325 27489 17359 27523
rect 17509 27489 17543 27523
rect 17693 27489 17727 27523
rect 19165 27489 19199 27523
rect 21741 27489 21775 27523
rect 21925 27489 21959 27523
rect 22017 27489 22051 27523
rect 23213 27489 23247 27523
rect 23305 27489 23339 27523
rect 23489 27489 23523 27523
rect 25145 27489 25179 27523
rect 25237 27489 25271 27523
rect 25881 27489 25915 27523
rect 27721 27489 27755 27523
rect 28089 27489 28123 27523
rect 28273 27489 28307 27523
rect 28825 27489 28859 27523
rect 29285 27489 29319 27523
rect 29745 27489 29779 27523
rect 31217 27489 31251 27523
rect 3249 27421 3283 27455
rect 7113 27421 7147 27455
rect 8125 27421 8159 27455
rect 10333 27421 10367 27455
rect 12081 27421 12115 27455
rect 12541 27421 12575 27455
rect 12909 27421 12943 27455
rect 13553 27421 13587 27455
rect 14197 27421 14231 27455
rect 14565 27421 14599 27455
rect 14749 27421 14783 27455
rect 15025 27421 15059 27455
rect 16497 27421 16531 27455
rect 18521 27421 18555 27455
rect 19257 27421 19291 27455
rect 20545 27421 20579 27455
rect 22845 27421 22879 27455
rect 24869 27421 24903 27455
rect 25789 27421 25823 27455
rect 26893 27421 26927 27455
rect 27997 27421 28031 27455
rect 29469 27421 29503 27455
rect 30665 27421 30699 27455
rect 31401 27421 31435 27455
rect 9689 27353 9723 27387
rect 11805 27353 11839 27387
rect 21925 27353 21959 27387
rect 23029 27353 23063 27387
rect 24133 27353 24167 27387
rect 24961 27353 24995 27387
rect 29101 27353 29135 27387
rect 5549 27285 5583 27319
rect 7757 27285 7791 27319
rect 8769 27285 8803 27319
rect 14013 27285 14047 27319
rect 17141 27285 17175 27319
rect 19073 27285 19107 27319
rect 19901 27285 19935 27319
rect 19993 27285 20027 27319
rect 22109 27285 22143 27319
rect 22293 27285 22327 27319
rect 24225 27285 24259 27319
rect 25513 27285 25547 27319
rect 25605 27285 25639 27319
rect 26065 27285 26099 27319
rect 26341 27285 26375 27319
rect 28181 27285 28215 27319
rect 28733 27285 28767 27319
rect 29653 27285 29687 27319
rect 30021 27285 30055 27319
rect 30941 27285 30975 27319
rect 7021 27081 7055 27115
rect 9597 27081 9631 27115
rect 10701 27081 10735 27115
rect 14933 27081 14967 27115
rect 23121 27081 23155 27115
rect 26328 27081 26362 27115
rect 27813 27081 27847 27115
rect 31033 27081 31067 27115
rect 8861 27013 8895 27047
rect 14657 27013 14691 27047
rect 23213 27013 23247 27047
rect 25789 27013 25823 27047
rect 29653 27013 29687 27047
rect 30481 27013 30515 27047
rect 8493 26945 8527 26979
rect 10885 26945 10919 26979
rect 11253 26945 11287 26979
rect 11345 26945 11379 26979
rect 11713 26945 11747 26979
rect 15117 26945 15151 26979
rect 15485 26945 15519 26979
rect 19809 26945 19843 26979
rect 20085 26945 20119 26979
rect 21373 26945 21407 26979
rect 21649 26945 21683 26979
rect 23857 26945 23891 26979
rect 25605 26945 25639 26979
rect 29101 26945 29135 26979
rect 30297 26945 30331 26979
rect 6837 26877 6871 26911
rect 8769 26877 8803 26911
rect 9413 26877 9447 26911
rect 9781 26877 9815 26911
rect 9873 26877 9907 26911
rect 10149 26877 10183 26911
rect 10977 26877 11011 26911
rect 14105 26877 14139 26911
rect 15209 26877 15243 26911
rect 16313 26877 16347 26911
rect 17325 26877 17359 26911
rect 24409 26877 24443 26911
rect 24501 26877 24535 26911
rect 25421 26877 25455 26911
rect 25881 26877 25915 26911
rect 26065 26877 26099 26911
rect 28457 26877 28491 26911
rect 28641 26877 28675 26911
rect 28825 26877 28859 26911
rect 30849 26877 30883 26911
rect 31769 26877 31803 26911
rect 9965 26809 9999 26843
rect 12081 26809 12115 26843
rect 12449 26809 12483 26843
rect 15577 26809 15611 26843
rect 16037 26809 16071 26843
rect 23581 26809 23615 26843
rect 24225 26809 24259 26843
rect 24777 26809 24811 26843
rect 24869 26809 24903 26843
rect 30757 26809 30791 26843
rect 6745 26741 6779 26775
rect 13921 26741 13955 26775
rect 16681 26741 16715 26775
rect 18337 26741 18371 26775
rect 23673 26741 23707 26775
rect 24593 26741 24627 26775
rect 25605 26741 25639 26775
rect 27905 26741 27939 26775
rect 28733 26741 28767 26775
rect 29193 26741 29227 26775
rect 29285 26741 29319 26775
rect 29745 26741 29779 26775
rect 30665 26741 30699 26775
rect 31493 26741 31527 26775
rect 5641 26537 5675 26571
rect 7757 26537 7791 26571
rect 8033 26537 8067 26571
rect 8401 26537 8435 26571
rect 8493 26537 8527 26571
rect 8861 26537 8895 26571
rect 10517 26537 10551 26571
rect 12265 26537 12299 26571
rect 14933 26537 14967 26571
rect 18153 26537 18187 26571
rect 19349 26537 19383 26571
rect 19717 26537 19751 26571
rect 19809 26537 19843 26571
rect 20177 26537 20211 26571
rect 23305 26537 23339 26571
rect 25237 26537 25271 26571
rect 26249 26537 26283 26571
rect 27353 26537 27387 26571
rect 27537 26537 27571 26571
rect 27813 26537 27847 26571
rect 30665 26537 30699 26571
rect 7113 26469 7147 26503
rect 9137 26469 9171 26503
rect 9229 26469 9263 26503
rect 10701 26469 10735 26503
rect 11529 26469 11563 26503
rect 18429 26469 18463 26503
rect 21833 26469 21867 26503
rect 26525 26469 26559 26503
rect 26617 26469 26651 26503
rect 26755 26469 26789 26503
rect 27169 26469 27203 26503
rect 29193 26469 29227 26503
rect 30849 26469 30883 26503
rect 4445 26401 4479 26435
rect 4537 26401 4571 26435
rect 7849 26401 7883 26435
rect 9045 26401 9079 26435
rect 9413 26401 9447 26435
rect 10609 26401 10643 26435
rect 10793 26401 10827 26435
rect 11345 26401 11379 26435
rect 11621 26401 11655 26435
rect 11713 26401 11747 26435
rect 15209 26401 15243 26435
rect 15945 26401 15979 26435
rect 16405 26401 16439 26435
rect 18521 26401 18555 26435
rect 20269 26401 20303 26435
rect 21557 26401 21591 26435
rect 23489 26401 23523 26435
rect 25605 26401 25639 26435
rect 25973 26401 26007 26435
rect 26433 26401 26467 26435
rect 26893 26401 26927 26435
rect 27445 26401 27479 26435
rect 27997 26401 28031 26435
rect 28273 26401 28307 26435
rect 28457 26401 28491 26435
rect 28825 26401 28859 26435
rect 30941 26401 30975 26435
rect 3249 26333 3283 26367
rect 7389 26333 7423 26367
rect 8585 26333 8619 26367
rect 11161 26333 11195 26367
rect 13369 26333 13403 26367
rect 14289 26333 14323 26367
rect 16681 26333 16715 26367
rect 19073 26333 19107 26367
rect 19257 26333 19291 26367
rect 20361 26333 20395 26367
rect 21189 26333 21223 26367
rect 23765 26333 23799 26367
rect 25513 26333 25547 26367
rect 28917 26333 28951 26367
rect 10149 26265 10183 26299
rect 14013 26265 14047 26299
rect 15577 26265 15611 26299
rect 26157 26265 26191 26299
rect 27721 26265 27755 26299
rect 5181 26197 5215 26231
rect 9689 26197 9723 26231
rect 11897 26197 11931 26231
rect 15117 26197 15151 26231
rect 16037 26197 16071 26231
rect 18797 26197 18831 26231
rect 20637 26197 20671 26231
rect 25881 26197 25915 26231
rect 28733 26197 28767 26231
rect 3525 25993 3559 26027
rect 10333 25993 10367 26027
rect 10885 25993 10919 26027
rect 12173 25993 12207 26027
rect 17785 25993 17819 26027
rect 18797 25993 18831 26027
rect 25237 25993 25271 26027
rect 30113 25993 30147 26027
rect 20913 25925 20947 25959
rect 5273 25857 5307 25891
rect 6745 25857 6779 25891
rect 9873 25857 9907 25891
rect 12909 25857 12943 25891
rect 14657 25857 14691 25891
rect 15301 25857 15335 25891
rect 17049 25857 17083 25891
rect 22109 25857 22143 25891
rect 24777 25857 24811 25891
rect 27537 25857 27571 25891
rect 29285 25857 29319 25891
rect 8493 25789 8527 25823
rect 9229 25789 9263 25823
rect 10701 25789 10735 25823
rect 10885 25789 10919 25823
rect 10977 25789 11011 25823
rect 11621 25789 11655 25823
rect 12817 25789 12851 25823
rect 14749 25789 14783 25823
rect 16313 25789 16347 25823
rect 17233 25789 17267 25823
rect 17509 25789 17543 25823
rect 17601 25789 17635 25823
rect 20545 25789 20579 25823
rect 21465 25789 21499 25823
rect 21833 25789 21867 25823
rect 25145 25789 25179 25823
rect 25789 25789 25823 25823
rect 29377 25789 29411 25823
rect 30297 25789 30331 25823
rect 30389 25789 30423 25823
rect 4997 25721 5031 25755
rect 8217 25721 8251 25755
rect 13185 25721 13219 25755
rect 17417 25721 17451 25755
rect 20269 25721 20303 25755
rect 21741 25721 21775 25755
rect 22385 25721 22419 25755
rect 26157 25721 26191 25755
rect 27813 25721 27847 25755
rect 5641 25653 5675 25687
rect 6193 25653 6227 25687
rect 8585 25653 8619 25687
rect 9321 25653 9355 25687
rect 11897 25653 11931 25687
rect 15761 25653 15795 25687
rect 16497 25653 16531 25687
rect 18061 25653 18095 25687
rect 18521 25653 18555 25687
rect 23857 25653 23891 25687
rect 26249 25653 26283 25687
rect 29561 25653 29595 25687
rect 4721 25449 4755 25483
rect 5089 25449 5123 25483
rect 6285 25449 6319 25483
rect 7113 25449 7147 25483
rect 7757 25449 7791 25483
rect 8033 25449 8067 25483
rect 8401 25449 8435 25483
rect 10609 25449 10643 25483
rect 13001 25449 13035 25483
rect 13461 25449 13495 25483
rect 13829 25449 13863 25483
rect 16681 25449 16715 25483
rect 22661 25449 22695 25483
rect 24869 25449 24903 25483
rect 24961 25449 24995 25483
rect 25697 25449 25731 25483
rect 26617 25449 26651 25483
rect 5825 25381 5859 25415
rect 5917 25381 5951 25415
rect 11529 25381 11563 25415
rect 13277 25381 13311 25415
rect 15209 25381 15243 25415
rect 16957 25381 16991 25415
rect 21465 25381 21499 25415
rect 22477 25381 22511 25415
rect 5181 25313 5215 25347
rect 5733 25313 5767 25347
rect 6101 25313 6135 25347
rect 6377 25313 6411 25347
rect 7849 25313 7883 25347
rect 8493 25313 8527 25347
rect 9965 25313 9999 25347
rect 10241 25313 10275 25347
rect 10333 25313 10367 25347
rect 10517 25313 10551 25347
rect 11161 25313 11195 25347
rect 13369 25313 13403 25347
rect 13921 25313 13955 25347
rect 14289 25313 14323 25347
rect 17785 25313 17819 25347
rect 18705 25313 18739 25347
rect 21557 25313 21591 25347
rect 22385 25313 22419 25347
rect 23673 25313 23707 25347
rect 23949 25313 23983 25347
rect 24133 25313 24167 25347
rect 24225 25313 24259 25347
rect 25145 25313 25179 25347
rect 25237 25313 25271 25347
rect 25421 25313 25455 25347
rect 25605 25313 25639 25347
rect 26065 25313 26099 25347
rect 28457 25313 28491 25347
rect 29653 25313 29687 25347
rect 30481 25313 30515 25347
rect 3433 25245 3467 25279
rect 5365 25245 5399 25279
rect 8585 25245 8619 25279
rect 9321 25245 9355 25279
rect 10885 25245 10919 25279
rect 11253 25245 11287 25279
rect 14013 25245 14047 25279
rect 14565 25245 14599 25279
rect 14933 25245 14967 25279
rect 18981 25245 19015 25279
rect 21281 25245 21315 25279
rect 23305 25245 23339 25279
rect 23489 25245 23523 25279
rect 31677 25245 31711 25279
rect 9045 25177 9079 25211
rect 20453 25177 20487 25211
rect 25329 25177 25363 25211
rect 28181 25177 28215 25211
rect 4077 25109 4111 25143
rect 5549 25109 5583 25143
rect 6745 25109 6779 25143
rect 10149 25109 10183 25143
rect 10333 25109 10367 25143
rect 10885 25109 10919 25143
rect 14565 25109 14599 25143
rect 14841 25109 14875 25143
rect 18153 25109 18187 25143
rect 20637 25109 20671 25143
rect 27997 25109 28031 25143
rect 29009 25109 29043 25143
rect 5917 24905 5951 24939
rect 7836 24905 7870 24939
rect 9321 24905 9355 24939
rect 9413 24905 9447 24939
rect 11713 24905 11747 24939
rect 15577 24905 15611 24939
rect 15761 24905 15795 24939
rect 19533 24905 19567 24939
rect 28181 24905 28215 24939
rect 30021 24905 30055 24939
rect 10333 24837 10367 24871
rect 3525 24769 3559 24803
rect 7573 24769 7607 24803
rect 11989 24769 12023 24803
rect 12633 24769 12667 24803
rect 14381 24769 14415 24803
rect 15025 24769 15059 24803
rect 16313 24769 16347 24803
rect 17693 24769 17727 24803
rect 19993 24769 20027 24803
rect 20085 24769 20119 24803
rect 23305 24769 23339 24803
rect 27721 24769 27755 24803
rect 28273 24769 28307 24803
rect 28549 24769 28583 24803
rect 3249 24701 3283 24735
rect 5273 24701 5307 24735
rect 5825 24701 5859 24735
rect 6469 24701 6503 24735
rect 7297 24701 7331 24735
rect 9597 24701 9631 24735
rect 9689 24701 9723 24735
rect 9965 24701 9999 24735
rect 10241 24701 10275 24735
rect 10793 24701 10827 24735
rect 10977 24701 11011 24735
rect 11161 24701 11195 24735
rect 11529 24701 11563 24735
rect 11805 24701 11839 24735
rect 11897 24701 11931 24735
rect 12081 24701 12115 24735
rect 12357 24701 12391 24735
rect 12541 24701 12575 24735
rect 14473 24701 14507 24735
rect 16129 24701 16163 24735
rect 19901 24701 19935 24735
rect 22569 24701 22603 24735
rect 23397 24701 23431 24735
rect 27813 24701 27847 24735
rect 27905 24701 27939 24735
rect 27997 24701 28031 24735
rect 30297 24701 30331 24735
rect 9781 24633 9815 24667
rect 10885 24633 10919 24667
rect 12909 24633 12943 24667
rect 17969 24633 18003 24667
rect 30205 24633 30239 24667
rect 4629 24565 4663 24599
rect 5733 24565 5767 24599
rect 6653 24565 6687 24599
rect 10609 24565 10643 24599
rect 11253 24565 11287 24599
rect 12449 24565 12483 24599
rect 16221 24565 16255 24599
rect 16773 24565 16807 24599
rect 17141 24565 17175 24599
rect 17509 24565 17543 24599
rect 19441 24565 19475 24599
rect 23121 24565 23155 24599
rect 3433 24361 3467 24395
rect 3893 24361 3927 24395
rect 6009 24361 6043 24395
rect 8677 24361 8711 24395
rect 13001 24361 13035 24395
rect 21373 24361 21407 24395
rect 22661 24361 22695 24395
rect 4537 24293 4571 24327
rect 9137 24293 9171 24327
rect 10885 24293 10919 24327
rect 13553 24293 13587 24327
rect 14381 24293 14415 24327
rect 14749 24293 14783 24327
rect 18153 24293 18187 24327
rect 18705 24293 18739 24327
rect 19073 24293 19107 24327
rect 19901 24293 19935 24327
rect 26985 24293 27019 24327
rect 3801 24225 3835 24259
rect 4261 24225 4295 24259
rect 8953 24225 8987 24259
rect 9045 24225 9079 24259
rect 9321 24225 9355 24259
rect 11161 24225 11195 24259
rect 11621 24225 11655 24259
rect 12449 24225 12483 24259
rect 17049 24225 17083 24259
rect 18521 24225 18555 24259
rect 18613 24225 18647 24259
rect 18889 24225 18923 24259
rect 19165 24225 19199 24259
rect 21557 24225 21591 24259
rect 22293 24225 22327 24259
rect 25153 24225 25187 24259
rect 25421 24225 25455 24259
rect 25605 24225 25639 24259
rect 26249 24225 26283 24259
rect 26525 24225 26559 24259
rect 26617 24225 26651 24259
rect 26801 24225 26835 24259
rect 3341 24157 3375 24191
rect 4077 24157 4111 24191
rect 12725 24157 12759 24191
rect 14473 24157 14507 24191
rect 16221 24157 16255 24191
rect 16865 24157 16899 24191
rect 17233 24157 17267 24191
rect 22109 24157 22143 24191
rect 22201 24157 22235 24191
rect 24317 24157 24351 24191
rect 28641 24157 28675 24191
rect 29285 24157 29319 24191
rect 31585 24157 31619 24191
rect 31861 24157 31895 24191
rect 18337 24089 18371 24123
rect 25789 24089 25823 24123
rect 6653 24021 6687 24055
rect 8769 24021 8803 24055
rect 9413 24021 9447 24055
rect 11897 24021 11931 24055
rect 12265 24021 12299 24055
rect 12817 24021 12851 24055
rect 16313 24021 16347 24055
rect 19441 24021 19475 24055
rect 21649 24021 21683 24055
rect 24869 24021 24903 24055
rect 25053 24021 25087 24055
rect 3157 23817 3191 23851
rect 7665 23817 7699 23851
rect 13001 23817 13035 23851
rect 14013 23817 14047 23851
rect 16589 23817 16623 23851
rect 18337 23817 18371 23851
rect 18429 23817 18463 23851
rect 25789 23817 25823 23851
rect 27629 23817 27663 23851
rect 16129 23749 16163 23783
rect 26433 23749 26467 23783
rect 29193 23749 29227 23783
rect 4629 23681 4663 23715
rect 4905 23681 4939 23715
rect 7021 23681 7055 23715
rect 8401 23681 8435 23715
rect 8677 23681 8711 23715
rect 12909 23681 12943 23715
rect 22569 23681 22603 23715
rect 25329 23681 25363 23715
rect 5181 23613 5215 23647
rect 6377 23613 6411 23647
rect 7941 23613 7975 23647
rect 8309 23613 8343 23647
rect 10425 23613 10459 23647
rect 13553 23613 13587 23647
rect 14105 23613 14139 23647
rect 14289 23613 14323 23647
rect 15301 23613 15335 23647
rect 15485 23613 15519 23647
rect 16313 23613 16347 23647
rect 16681 23613 16715 23647
rect 17601 23613 17635 23647
rect 18613 23613 18647 23647
rect 18705 23613 18739 23647
rect 19717 23613 19751 23647
rect 20453 23613 20487 23647
rect 21557 23613 21591 23647
rect 21833 23613 21867 23647
rect 23029 23613 23063 23647
rect 25605 23613 25639 23647
rect 25881 23613 25915 23647
rect 26065 23613 26099 23647
rect 26249 23613 26283 23647
rect 26341 23613 26375 23647
rect 26433 23613 26467 23647
rect 26617 23623 26651 23657
rect 26709 23613 26743 23647
rect 26893 23613 26927 23647
rect 27720 23613 27754 23647
rect 27813 23613 27847 23647
rect 5089 23545 5123 23579
rect 8033 23545 8067 23579
rect 8125 23545 8159 23579
rect 10333 23545 10367 23579
rect 15117 23545 15151 23579
rect 25053 23545 25087 23579
rect 28917 23545 28951 23579
rect 5733 23477 5767 23511
rect 6469 23477 6503 23511
rect 7757 23477 7791 23511
rect 10149 23477 10183 23511
rect 12541 23477 12575 23511
rect 15393 23477 15427 23511
rect 15945 23477 15979 23511
rect 16957 23477 16991 23511
rect 17969 23477 18003 23511
rect 18889 23477 18923 23511
rect 19073 23477 19107 23511
rect 20361 23477 20395 23511
rect 21005 23477 21039 23511
rect 23121 23477 23155 23511
rect 23581 23477 23615 23511
rect 25421 23477 25455 23511
rect 27077 23477 27111 23511
rect 29377 23477 29411 23511
rect 3985 23273 4019 23307
rect 6193 23273 6227 23307
rect 6561 23273 6595 23307
rect 12909 23273 12943 23307
rect 13185 23273 13219 23307
rect 15025 23273 15059 23307
rect 17601 23273 17635 23307
rect 18521 23273 18555 23307
rect 25237 23273 25271 23307
rect 30389 23273 30423 23307
rect 5457 23205 5491 23239
rect 7021 23205 7055 23239
rect 8769 23205 8803 23239
rect 10701 23205 10735 23239
rect 10977 23205 11011 23239
rect 11345 23205 11379 23239
rect 13469 23205 13503 23239
rect 14657 23205 14691 23239
rect 19257 23205 19291 23239
rect 21005 23205 21039 23239
rect 5733 23137 5767 23171
rect 7757 23137 7791 23171
rect 9505 23137 9539 23171
rect 13323 23137 13357 23171
rect 13553 23137 13587 23171
rect 13737 23137 13771 23171
rect 14401 23137 14435 23171
rect 14565 23137 14599 23171
rect 14749 23137 14783 23171
rect 17693 23137 17727 23171
rect 24225 23137 24259 23171
rect 24409 23137 24443 23171
rect 24685 23137 24719 23171
rect 25053 23137 25087 23171
rect 25727 23137 25761 23171
rect 25835 23137 25869 23171
rect 26341 23137 26375 23171
rect 26709 23137 26743 23171
rect 26801 23137 26835 23171
rect 27261 23137 27295 23171
rect 27445 23137 27479 23171
rect 28641 23137 28675 23171
rect 31309 23137 31343 23171
rect 5917 23069 5951 23103
rect 6101 23069 6135 23103
rect 8677 23069 8711 23103
rect 9965 23069 9999 23103
rect 12265 23069 12299 23103
rect 12633 23069 12667 23103
rect 15577 23069 15611 23103
rect 15853 23069 15887 23103
rect 16129 23069 16163 23103
rect 17969 23069 18003 23103
rect 19073 23069 19107 23103
rect 21281 23069 21315 23103
rect 22845 23069 22879 23103
rect 23121 23069 23155 23103
rect 24041 23069 24075 23103
rect 24593 23069 24627 23103
rect 25329 23069 25363 23103
rect 27629 23069 27663 23103
rect 28917 23069 28951 23103
rect 30665 23069 30699 23103
rect 14933 23001 14967 23035
rect 25881 23001 25915 23035
rect 26249 23001 26283 23035
rect 7205 22933 7239 22967
rect 8033 22933 8067 22967
rect 14013 22933 14047 22967
rect 21373 22933 21407 22967
rect 23489 22933 23523 22967
rect 24409 22933 24443 22967
rect 25053 22933 25087 22967
rect 5089 22729 5123 22763
rect 7646 22729 7680 22763
rect 9137 22729 9171 22763
rect 14289 22729 14323 22763
rect 14473 22729 14507 22763
rect 14749 22729 14783 22763
rect 16681 22729 16715 22763
rect 20913 22729 20947 22763
rect 22385 22729 22419 22763
rect 22832 22729 22866 22763
rect 24317 22729 24351 22763
rect 27629 22729 27663 22763
rect 28733 22729 28767 22763
rect 29101 22729 29135 22763
rect 29837 22729 29871 22763
rect 15577 22661 15611 22695
rect 15853 22661 15887 22695
rect 18889 22661 18923 22695
rect 29469 22661 29503 22695
rect 7113 22593 7147 22627
rect 12541 22593 12575 22627
rect 16037 22593 16071 22627
rect 16957 22593 16991 22627
rect 17233 22593 17267 22627
rect 19349 22593 19383 22627
rect 19441 22593 19475 22627
rect 21465 22593 21499 22627
rect 28181 22593 28215 22627
rect 29193 22593 29227 22627
rect 4445 22525 4479 22559
rect 5181 22525 5215 22559
rect 6101 22525 6135 22559
rect 6377 22525 6411 22559
rect 7389 22525 7423 22559
rect 9781 22525 9815 22559
rect 10149 22525 10183 22559
rect 10701 22525 10735 22559
rect 11621 22525 11655 22559
rect 12817 22525 12851 22559
rect 14105 22525 14139 22559
rect 14473 22525 14507 22559
rect 14657 22525 14691 22559
rect 14749 22525 14783 22559
rect 14933 22525 14967 22559
rect 15025 22525 15059 22559
rect 15301 22525 15335 22559
rect 15393 22525 15427 22559
rect 15761 22525 15795 22559
rect 19257 22525 19291 22559
rect 19901 22525 19935 22559
rect 20729 22525 20763 22559
rect 21741 22525 21775 22559
rect 22569 22525 22603 22559
rect 24409 22525 24443 22559
rect 25416 22525 25450 22559
rect 25513 22525 25547 22559
rect 25788 22525 25822 22559
rect 25881 22525 25915 22559
rect 26065 22525 26099 22559
rect 26801 22525 26835 22559
rect 27077 22525 27111 22559
rect 27445 22525 27479 22559
rect 27629 22525 27663 22559
rect 27721 22525 27755 22559
rect 27905 22525 27939 22559
rect 28917 22525 28951 22559
rect 29285 22525 29319 22559
rect 29929 22525 29963 22559
rect 3249 22457 3283 22491
rect 6929 22457 6963 22491
rect 10057 22457 10091 22491
rect 12449 22457 12483 22491
rect 13553 22457 13587 22491
rect 15209 22457 15243 22491
rect 21281 22457 21315 22491
rect 25053 22457 25087 22491
rect 25605 22457 25639 22491
rect 5457 22389 5491 22423
rect 6285 22389 6319 22423
rect 6561 22389 6595 22423
rect 7021 22389 7055 22423
rect 9229 22389 9263 22423
rect 10793 22389 10827 22423
rect 11069 22389 11103 22423
rect 11989 22389 12023 22423
rect 12357 22389 12391 22423
rect 13461 22389 13495 22423
rect 18705 22389 18739 22423
rect 19809 22389 19843 22423
rect 20085 22389 20119 22423
rect 21373 22389 21407 22423
rect 25237 22389 25271 22423
rect 27261 22389 27295 22423
rect 27813 22389 27847 22423
rect 7849 22185 7883 22219
rect 10517 22185 10551 22219
rect 12725 22185 12759 22219
rect 13461 22185 13495 22219
rect 13553 22185 13587 22219
rect 17969 22185 18003 22219
rect 21649 22185 21683 22219
rect 23673 22185 23707 22219
rect 24317 22185 24351 22219
rect 25053 22185 25087 22219
rect 27261 22185 27295 22219
rect 4537 22117 4571 22151
rect 6377 22117 6411 22151
rect 11253 22117 11287 22151
rect 20269 22117 20303 22151
rect 21741 22117 21775 22151
rect 22937 22117 22971 22151
rect 25303 22117 25337 22151
rect 25513 22117 25547 22151
rect 26801 22117 26835 22151
rect 27353 22117 27387 22151
rect 8677 22049 8711 22083
rect 9045 22049 9079 22083
rect 10057 22049 10091 22083
rect 10609 22049 10643 22083
rect 13001 22049 13035 22083
rect 15025 22049 15059 22083
rect 15301 22049 15335 22083
rect 15853 22049 15887 22083
rect 18061 22049 18095 22083
rect 23121 22049 23155 22083
rect 23949 22049 23983 22083
rect 25420 22049 25454 22083
rect 25605 22049 25639 22083
rect 27721 22049 27755 22083
rect 27997 22049 28031 22083
rect 28181 22049 28215 22083
rect 30481 22049 30515 22083
rect 31677 22049 31711 22083
rect 3525 21981 3559 22015
rect 4261 21981 4295 22015
rect 6101 21981 6135 22015
rect 8309 21981 8343 22015
rect 10793 21981 10827 22015
rect 10977 21981 11011 22015
rect 13369 21981 13403 22015
rect 14565 21981 14599 22015
rect 16129 21981 16163 22015
rect 20545 21981 20579 22015
rect 21189 21981 21223 22015
rect 22477 21981 22511 22015
rect 23857 21981 23891 22015
rect 24501 21981 24535 22015
rect 25145 21981 25179 22015
rect 26065 21981 26099 22015
rect 27445 21981 27479 22015
rect 13921 21913 13955 21947
rect 18705 21913 18739 21947
rect 4169 21845 4203 21879
rect 6009 21845 6043 21879
rect 9965 21845 9999 21879
rect 10149 21845 10183 21879
rect 12909 21845 12943 21879
rect 14013 21845 14047 21879
rect 14749 21845 14783 21879
rect 14933 21845 14967 21879
rect 15577 21845 15611 21879
rect 17601 21845 17635 21879
rect 18797 21845 18831 21879
rect 20637 21845 20671 21879
rect 23213 21845 23247 21879
rect 25789 21845 25823 21879
rect 26893 21845 26927 21879
rect 27813 21845 27847 21879
rect 3157 21641 3191 21675
rect 6745 21641 6779 21675
rect 7481 21641 7515 21675
rect 7941 21641 7975 21675
rect 8309 21641 8343 21675
rect 11805 21641 11839 21675
rect 11989 21641 12023 21675
rect 13479 21641 13513 21675
rect 15209 21641 15243 21675
rect 16313 21641 16347 21675
rect 18245 21641 18279 21675
rect 20361 21641 20395 21675
rect 20913 21641 20947 21675
rect 25513 21641 25547 21675
rect 26249 21641 26283 21675
rect 14657 21573 14691 21607
rect 24593 21573 24627 21607
rect 5089 21505 5123 21539
rect 6009 21505 6043 21539
rect 6653 21505 6687 21539
rect 8677 21505 8711 21539
rect 13737 21505 13771 21539
rect 14289 21505 14323 21539
rect 15025 21505 15059 21539
rect 19809 21505 19843 21539
rect 22385 21505 22419 21539
rect 22753 21505 22787 21539
rect 26433 21505 26467 21539
rect 26709 21505 26743 21539
rect 28641 21505 28675 21539
rect 4905 21437 4939 21471
rect 5181 21437 5215 21471
rect 5733 21437 5767 21471
rect 6929 21437 6963 21471
rect 7021 21437 7055 21471
rect 7113 21437 7147 21471
rect 7297 21437 7331 21471
rect 7573 21437 7607 21471
rect 11437 21437 11471 21471
rect 11713 21437 11747 21471
rect 14473 21437 14507 21471
rect 14565 21437 14599 21471
rect 14841 21437 14875 21471
rect 15301 21437 15335 21471
rect 15761 21437 15795 21471
rect 16129 21437 16163 21471
rect 16957 21437 16991 21471
rect 17877 21437 17911 21471
rect 18153 21437 18187 21471
rect 19993 21437 20027 21471
rect 20545 21437 20579 21471
rect 22661 21437 22695 21471
rect 23305 21437 23339 21471
rect 24133 21437 24167 21471
rect 24225 21437 24259 21471
rect 24409 21437 24443 21471
rect 24685 21437 24719 21471
rect 25329 21437 25363 21471
rect 28457 21437 28491 21471
rect 28733 21437 28767 21471
rect 4629 21369 4663 21403
rect 8953 21369 8987 21403
rect 10885 21369 10919 21403
rect 14105 21369 14139 21403
rect 15945 21369 15979 21403
rect 16037 21369 16071 21403
rect 16497 21369 16531 21403
rect 17141 21369 17175 21403
rect 20637 21369 20671 21403
rect 25697 21369 25731 21403
rect 25881 21369 25915 21403
rect 28365 21369 28399 21403
rect 5825 21301 5859 21335
rect 10425 21301 10459 21335
rect 14565 21301 14599 21335
rect 16589 21301 16623 21335
rect 19901 21301 19935 21335
rect 23489 21301 23523 21335
rect 24777 21301 24811 21335
rect 28181 21301 28215 21335
rect 4537 21097 4571 21131
rect 4905 21097 4939 21131
rect 11529 21097 11563 21131
rect 14289 21097 14323 21131
rect 15853 21097 15887 21131
rect 22017 21097 22051 21131
rect 22477 21097 22511 21131
rect 23765 21097 23799 21131
rect 25329 21097 25363 21131
rect 10057 21029 10091 21063
rect 12173 21029 12207 21063
rect 12725 21029 12759 21063
rect 13921 21029 13955 21063
rect 16497 21029 16531 21063
rect 20085 21029 20119 21063
rect 20453 21029 20487 21063
rect 21557 21029 21591 21063
rect 22109 21029 22143 21063
rect 25145 21029 25179 21063
rect 3341 20961 3375 20995
rect 4445 20961 4479 20995
rect 6193 20961 6227 20995
rect 9781 20961 9815 20995
rect 13461 20961 13495 20995
rect 14038 20961 14072 20995
rect 14841 20961 14875 20995
rect 15485 20961 15519 20995
rect 23673 20961 23707 20995
rect 24133 20961 24167 20995
rect 24317 20961 24351 20995
rect 24409 20961 24443 20995
rect 24593 20961 24627 20995
rect 24777 20961 24811 20995
rect 25053 20961 25087 20995
rect 25421 20961 25455 20995
rect 28181 20961 28215 20995
rect 31861 20961 31895 20995
rect 3065 20893 3099 20927
rect 4261 20893 4295 20927
rect 5825 20893 5859 20927
rect 6745 20893 6779 20927
rect 12265 20893 12299 20927
rect 13553 20893 13587 20927
rect 13829 20893 13863 20927
rect 15209 20893 15243 20927
rect 15301 20893 15335 20927
rect 15393 20893 15427 20927
rect 18337 20893 18371 20927
rect 20361 20893 20395 20927
rect 21005 20893 21039 20927
rect 21925 20893 21959 20927
rect 25513 20893 25547 20927
rect 25789 20893 25823 20927
rect 26065 20893 26099 20927
rect 27537 20893 27571 20927
rect 29193 20893 29227 20927
rect 29469 20893 29503 20927
rect 30665 20893 30699 20927
rect 12725 20825 12759 20859
rect 14197 20825 14231 20859
rect 24225 20825 24259 20859
rect 31677 20825 31711 20859
rect 5273 20757 5307 20791
rect 11989 20757 12023 20791
rect 15025 20757 15059 20791
rect 16865 20757 16899 20791
rect 23949 20757 23983 20791
rect 24869 20757 24903 20791
rect 25697 20757 25731 20791
rect 27629 20757 27663 20791
rect 28641 20757 28675 20791
rect 30021 20757 30055 20791
rect 30113 20757 30147 20791
rect 4813 20553 4847 20587
rect 5457 20553 5491 20587
rect 10425 20553 10459 20587
rect 11621 20553 11655 20587
rect 14197 20553 14231 20587
rect 15945 20553 15979 20587
rect 18889 20553 18923 20587
rect 19165 20553 19199 20587
rect 20085 20553 20119 20587
rect 24409 20553 24443 20587
rect 24777 20553 24811 20587
rect 25145 20553 25179 20587
rect 25605 20553 25639 20587
rect 26690 20553 26724 20587
rect 28181 20553 28215 20587
rect 30573 20553 30607 20587
rect 10609 20485 10643 20519
rect 26157 20485 26191 20519
rect 6101 20417 6135 20451
rect 7849 20417 7883 20451
rect 7941 20417 7975 20451
rect 8677 20417 8711 20451
rect 11161 20417 11195 20451
rect 11989 20417 12023 20451
rect 12474 20417 12508 20451
rect 15485 20417 15519 20451
rect 19533 20417 19567 20451
rect 22845 20417 22879 20451
rect 23581 20417 23615 20451
rect 24041 20417 24075 20451
rect 24685 20417 24719 20451
rect 25513 20417 25547 20451
rect 26433 20417 26467 20451
rect 30297 20417 30331 20451
rect 5641 20349 5675 20383
rect 5733 20349 5767 20383
rect 6009 20349 6043 20383
rect 10977 20349 11011 20383
rect 12357 20349 12391 20383
rect 14013 20349 14047 20383
rect 14105 20349 14139 20383
rect 15025 20349 15059 20383
rect 19073 20349 19107 20383
rect 19625 20349 19659 20383
rect 23305 20349 23339 20383
rect 23397 20349 23431 20383
rect 23489 20349 23523 20383
rect 23857 20349 23891 20383
rect 23949 20349 23983 20383
rect 24133 20349 24167 20383
rect 24961 20349 24995 20383
rect 25421 20349 25455 20383
rect 25697 20349 25731 20383
rect 25881 20349 25915 20383
rect 26065 20349 26099 20383
rect 28273 20349 28307 20383
rect 5825 20281 5859 20315
rect 6377 20281 6411 20315
rect 8953 20281 8987 20315
rect 11069 20281 11103 20315
rect 22569 20281 22603 20315
rect 30021 20281 30055 20315
rect 5273 20213 5307 20247
rect 8585 20213 8619 20247
rect 12265 20213 12299 20247
rect 12633 20213 12667 20247
rect 13645 20213 13679 20247
rect 13921 20213 13955 20247
rect 14657 20213 14691 20247
rect 19717 20213 19751 20247
rect 21097 20213 21131 20247
rect 23121 20213 23155 20247
rect 24317 20213 24351 20247
rect 30941 20213 30975 20247
rect 31401 20213 31435 20247
rect 6469 20009 6503 20043
rect 7113 20009 7147 20043
rect 8033 20009 8067 20043
rect 9413 20009 9447 20043
rect 10149 20009 10183 20043
rect 14381 20009 14415 20043
rect 14841 20009 14875 20043
rect 15209 20009 15243 20043
rect 19257 20009 19291 20043
rect 20453 20009 20487 20043
rect 22109 20009 22143 20043
rect 23673 20009 23707 20043
rect 26341 20009 26375 20043
rect 29009 20009 29043 20043
rect 29377 20009 29411 20043
rect 4997 19941 5031 19975
rect 8309 19941 8343 19975
rect 8401 19941 8435 19975
rect 14565 19941 14599 19975
rect 15025 19941 15059 19975
rect 16221 19941 16255 19975
rect 22753 19941 22787 19975
rect 28917 19941 28951 19975
rect 7021 19873 7055 19907
rect 8217 19873 8251 19907
rect 8585 19873 8619 19907
rect 9597 19873 9631 19907
rect 9689 19873 9723 19907
rect 9781 19873 9815 19907
rect 9965 19873 9999 19907
rect 10241 19873 10275 19907
rect 10793 19873 10827 19907
rect 11437 19873 11471 19907
rect 13553 19873 13587 19907
rect 14197 19873 14231 19907
rect 14749 19873 14783 19907
rect 15117 19873 15151 19907
rect 15579 19873 15613 19907
rect 17969 19873 18003 19907
rect 18521 19873 18555 19907
rect 21097 19873 21131 19907
rect 22201 19873 22235 19907
rect 22477 19873 22511 19907
rect 22661 19873 22695 19907
rect 22937 19873 22971 19907
rect 23029 19873 23063 19907
rect 23213 19873 23247 19907
rect 24041 19873 24075 19907
rect 24501 19873 24535 19907
rect 26065 19873 26099 19907
rect 26525 19873 26559 19907
rect 27537 19873 27571 19907
rect 27813 19873 27847 19907
rect 27905 19873 27939 19907
rect 28089 19873 28123 19907
rect 29653 19873 29687 19907
rect 30665 19873 30699 19907
rect 30824 19873 30858 19907
rect 30941 19873 30975 19907
rect 31861 19873 31895 19907
rect 4721 19805 4755 19839
rect 6837 19805 6871 19839
rect 13277 19805 13311 19839
rect 13369 19805 13403 19839
rect 13461 19805 13495 19839
rect 13737 19805 13771 19839
rect 14289 19805 14323 19839
rect 14657 19805 14691 19839
rect 15945 19805 15979 19839
rect 21741 19805 21775 19839
rect 24133 19805 24167 19839
rect 24593 19805 24627 19839
rect 25789 19805 25823 19839
rect 28825 19805 28859 19839
rect 31677 19805 31711 19839
rect 15025 19737 15059 19771
rect 15393 19737 15427 19771
rect 22661 19737 22695 19771
rect 23121 19737 23155 19771
rect 27997 19737 28031 19771
rect 31217 19737 31251 19771
rect 9229 19669 9263 19703
rect 10609 19669 10643 19703
rect 14013 19669 14047 19703
rect 17877 19669 17911 19703
rect 18429 19669 18463 19703
rect 21189 19669 21223 19703
rect 24869 19669 24903 19703
rect 25145 19669 25179 19703
rect 25973 19669 26007 19703
rect 27261 19669 27295 19703
rect 28273 19669 28307 19703
rect 29561 19669 29595 19703
rect 30021 19669 30055 19703
rect 21649 19465 21683 19499
rect 23949 19465 23983 19499
rect 24133 19465 24167 19499
rect 26249 19465 26283 19499
rect 27537 19465 27571 19499
rect 28549 19465 28583 19499
rect 28917 19465 28951 19499
rect 14289 19397 14323 19431
rect 19993 19397 20027 19431
rect 8493 19329 8527 19363
rect 9413 19329 9447 19363
rect 20545 19329 20579 19363
rect 23121 19329 23155 19363
rect 24041 19329 24075 19363
rect 26341 19329 26375 19363
rect 27721 19329 27755 19363
rect 27813 19329 27847 19363
rect 27905 19329 27939 19363
rect 27997 19329 28031 19363
rect 3065 19261 3099 19295
rect 7849 19261 7883 19295
rect 9137 19261 9171 19295
rect 10701 19261 10735 19295
rect 11805 19261 11839 19295
rect 12541 19261 12575 19295
rect 14657 19261 14691 19295
rect 15393 19261 15427 19295
rect 15577 19261 15611 19295
rect 16773 19261 16807 19295
rect 17041 19263 17075 19297
rect 17130 19261 17164 19295
rect 19901 19261 19935 19295
rect 20361 19261 20395 19295
rect 23397 19261 23431 19295
rect 23857 19261 23891 19295
rect 24317 19261 24351 19295
rect 24961 19261 24995 19295
rect 25145 19261 25179 19295
rect 26617 19261 26651 19295
rect 27445 19261 27479 19295
rect 28181 19261 28215 19295
rect 28365 19261 28399 19295
rect 28641 19261 28675 19295
rect 29285 19261 29319 19295
rect 31769 19261 31803 19295
rect 12817 19193 12851 19227
rect 17417 19193 17451 19227
rect 19165 19193 19199 19227
rect 21097 19193 21131 19227
rect 21465 19193 21499 19227
rect 29561 19193 29595 19227
rect 3249 19125 3283 19159
rect 8769 19125 8803 19159
rect 9229 19125 9263 19159
rect 10057 19125 10091 19159
rect 11345 19125 11379 19159
rect 11989 19125 12023 19159
rect 14841 19125 14875 19159
rect 15301 19125 15335 19159
rect 15577 19125 15611 19159
rect 16129 19125 16163 19159
rect 16957 19125 16991 19159
rect 19257 19125 19291 19159
rect 20453 19125 20487 19159
rect 21373 19125 21407 19159
rect 23581 19125 23615 19159
rect 24409 19125 24443 19159
rect 25789 19125 25823 19159
rect 26065 19125 26099 19159
rect 27261 19125 27295 19159
rect 28181 19125 28215 19159
rect 31033 19125 31067 19159
rect 31217 19125 31251 19159
rect 7849 18921 7883 18955
rect 8493 18921 8527 18955
rect 9781 18921 9815 18955
rect 13185 18921 13219 18955
rect 13645 18921 13679 18955
rect 14473 18921 14507 18955
rect 17325 18921 17359 18955
rect 22661 18921 22695 18955
rect 23213 18921 23247 18955
rect 24685 18921 24719 18955
rect 29377 18921 29411 18955
rect 30297 18921 30331 18955
rect 9045 18853 9079 18887
rect 19625 18853 19659 18887
rect 25145 18853 25179 18887
rect 29745 18853 29779 18887
rect 31677 18853 31711 18887
rect 8585 18785 8619 18819
rect 9597 18785 9631 18819
rect 10885 18785 10919 18819
rect 12081 18785 12115 18819
rect 13553 18785 13587 18819
rect 14105 18785 14139 18819
rect 15025 18785 15059 18819
rect 15209 18785 15243 18819
rect 17693 18785 17727 18819
rect 18429 18785 18463 18819
rect 21649 18785 21683 18819
rect 22753 18785 22787 18819
rect 23121 18785 23155 18819
rect 23305 18785 23339 18819
rect 24593 18785 24627 18819
rect 24777 18785 24811 18819
rect 24869 18785 24903 18819
rect 28365 18785 28399 18819
rect 30205 18785 30239 18819
rect 30665 18785 30699 18819
rect 4721 18717 4755 18751
rect 4997 18717 5031 18751
rect 7113 18717 7147 18751
rect 8769 18717 8803 18751
rect 9505 18717 9539 18751
rect 9873 18717 9907 18751
rect 12541 18717 12575 18751
rect 12633 18717 12667 18751
rect 13001 18717 13035 18751
rect 13737 18717 13771 18751
rect 14381 18717 14415 18751
rect 15485 18717 15519 18751
rect 17785 18717 17819 18751
rect 17877 18717 17911 18751
rect 19073 18717 19107 18751
rect 19349 18717 19383 18751
rect 21097 18717 21131 18751
rect 24501 18717 24535 18751
rect 26617 18717 26651 18751
rect 26893 18717 26927 18751
rect 27813 18717 27847 18751
rect 29837 18717 29871 18751
rect 29929 18717 29963 18751
rect 6561 18649 6595 18683
rect 9045 18649 9079 18683
rect 12173 18649 12207 18683
rect 14197 18649 14231 18683
rect 27537 18649 27571 18683
rect 6469 18581 6503 18615
rect 8125 18581 8159 18615
rect 10517 18581 10551 18615
rect 12357 18581 12391 18615
rect 14105 18581 14139 18615
rect 16957 18581 16991 18615
rect 21557 18581 21591 18615
rect 23857 18581 23891 18615
rect 28273 18581 28307 18615
rect 29009 18581 29043 18615
rect 5457 18377 5491 18411
rect 6377 18377 6411 18411
rect 6745 18377 6779 18411
rect 8388 18377 8422 18411
rect 9873 18377 9907 18411
rect 11897 18377 11931 18411
rect 12173 18377 12207 18411
rect 14105 18377 14139 18411
rect 15761 18377 15795 18411
rect 20177 18377 20211 18411
rect 23489 18377 23523 18411
rect 24593 18377 24627 18411
rect 25053 18377 25087 18411
rect 25881 18377 25915 18411
rect 26433 18377 26467 18411
rect 28273 18377 28307 18411
rect 10609 18309 10643 18343
rect 18981 18309 19015 18343
rect 19073 18309 19107 18343
rect 21741 18309 21775 18343
rect 27353 18309 27387 18343
rect 6009 18241 6043 18275
rect 7941 18241 7975 18275
rect 18889 18241 18923 18275
rect 21097 18241 21131 18275
rect 22385 18241 22419 18275
rect 23673 18241 23707 18275
rect 23949 18241 23983 18275
rect 26801 18241 26835 18275
rect 26893 18241 26927 18275
rect 27445 18241 27479 18275
rect 29193 18241 29227 18275
rect 5825 18173 5859 18207
rect 6469 18173 6503 18207
rect 8125 18173 8159 18207
rect 10149 18173 10183 18207
rect 10425 18173 10459 18207
rect 11161 18173 11195 18207
rect 12081 18173 12115 18207
rect 12265 18173 12299 18207
rect 12357 18173 12391 18207
rect 14289 18173 14323 18207
rect 14933 18173 14967 18207
rect 15945 18173 15979 18207
rect 16037 18173 16071 18207
rect 16497 18173 16531 18207
rect 16589 18173 16623 18207
rect 16773 18173 16807 18207
rect 16865 18173 16899 18207
rect 17141 18173 17175 18207
rect 19717 18173 19751 18207
rect 19993 18173 20027 18207
rect 20085 18173 20119 18207
rect 20269 18173 20303 18207
rect 20545 18173 20579 18207
rect 22569 18173 22603 18207
rect 23765 18173 23799 18207
rect 23857 18173 23891 18207
rect 24409 18173 24443 18207
rect 24593 18173 24627 18207
rect 24961 18173 24995 18207
rect 25329 18173 25363 18207
rect 26249 18173 26283 18207
rect 26433 18173 26467 18207
rect 26985 18173 27019 18207
rect 28917 18173 28951 18207
rect 29929 18173 29963 18207
rect 30849 18173 30883 18207
rect 31401 18173 31435 18207
rect 12633 18105 12667 18139
rect 19441 18105 19475 18139
rect 19625 18105 19659 18139
rect 21373 18105 21407 18139
rect 30205 18105 30239 18139
rect 31769 18105 31803 18139
rect 5917 18037 5951 18071
rect 7297 18037 7331 18071
rect 7665 18037 7699 18071
rect 7757 18037 7791 18071
rect 11529 18037 11563 18071
rect 14841 18037 14875 18071
rect 15577 18037 15611 18071
rect 16405 18037 16439 18071
rect 17049 18037 17083 18071
rect 19901 18037 19935 18071
rect 21281 18037 21315 18071
rect 21833 18037 21867 18071
rect 23213 18037 23247 18071
rect 28089 18037 28123 18071
rect 10241 17833 10275 17867
rect 10609 17833 10643 17867
rect 11345 17833 11379 17867
rect 12449 17833 12483 17867
rect 13385 17833 13419 17867
rect 13737 17833 13771 17867
rect 16865 17833 16899 17867
rect 22385 17833 22419 17867
rect 22845 17833 22879 17867
rect 25513 17833 25547 17867
rect 25973 17833 26007 17867
rect 28825 17833 28859 17867
rect 30021 17833 30055 17867
rect 10149 17765 10183 17799
rect 10358 17765 10392 17799
rect 13185 17765 13219 17799
rect 14013 17765 14047 17799
rect 16773 17765 16807 17799
rect 17937 17765 17971 17799
rect 18153 17765 18187 17799
rect 21741 17765 21775 17799
rect 22753 17765 22787 17799
rect 24041 17765 24075 17799
rect 25881 17765 25915 17799
rect 28181 17765 28215 17799
rect 29193 17765 29227 17799
rect 6101 17697 6135 17731
rect 8033 17697 8067 17731
rect 9873 17697 9907 17731
rect 11897 17697 11931 17731
rect 12633 17697 12667 17731
rect 12817 17697 12851 17731
rect 12909 17697 12943 17731
rect 13829 17697 13863 17731
rect 14289 17697 14323 17731
rect 14565 17697 14599 17731
rect 15761 17697 15795 17731
rect 15853 17697 15887 17731
rect 16313 17697 16347 17731
rect 16957 17697 16991 17731
rect 17601 17697 17635 17731
rect 19074 17719 19108 17753
rect 26433 17697 26467 17731
rect 29929 17697 29963 17731
rect 30665 17697 30699 17731
rect 6377 17629 6411 17663
rect 8309 17629 8343 17663
rect 11161 17629 11195 17663
rect 11621 17629 11655 17663
rect 12725 17629 12759 17663
rect 14381 17629 14415 17663
rect 15117 17629 15151 17663
rect 15301 17629 15335 17663
rect 15393 17629 15427 17663
rect 16405 17629 16439 17663
rect 17141 17629 17175 17663
rect 18889 17629 18923 17663
rect 19165 17629 19199 17663
rect 19349 17629 19383 17663
rect 19533 17629 19567 17663
rect 20269 17629 20303 17663
rect 22017 17629 22051 17663
rect 23029 17629 23063 17663
rect 23765 17629 23799 17663
rect 25789 17629 25823 17663
rect 28457 17629 28491 17663
rect 30113 17629 30147 17663
rect 31677 17629 31711 17663
rect 7849 17561 7883 17595
rect 9781 17561 9815 17595
rect 19257 17561 19291 17595
rect 10517 17493 10551 17527
rect 11805 17493 11839 17527
rect 12357 17493 12391 17527
rect 13369 17493 13403 17527
rect 13553 17493 13587 17527
rect 14013 17493 14047 17527
rect 14197 17493 14231 17527
rect 17509 17493 17543 17527
rect 17785 17493 17819 17527
rect 17969 17493 18003 17527
rect 18337 17493 18371 17527
rect 20085 17493 20119 17527
rect 26341 17493 26375 17527
rect 29561 17493 29595 17527
rect 9321 17289 9355 17323
rect 11897 17289 11931 17323
rect 13093 17289 13127 17323
rect 13277 17289 13311 17323
rect 13921 17289 13955 17323
rect 14197 17289 14231 17323
rect 16313 17289 16347 17323
rect 18889 17289 18923 17323
rect 21005 17289 21039 17323
rect 24869 17289 24903 17323
rect 28825 17289 28859 17323
rect 29239 17289 29273 17323
rect 31217 17289 31251 17323
rect 9229 17221 9263 17255
rect 16865 17221 16899 17255
rect 7757 17153 7791 17187
rect 9781 17153 9815 17187
rect 9965 17153 9999 17187
rect 20637 17153 20671 17187
rect 23029 17153 23063 17187
rect 28181 17153 28215 17187
rect 31033 17153 31067 17187
rect 7481 17085 7515 17119
rect 10977 17085 11011 17119
rect 11989 17085 12023 17119
rect 12265 17085 12299 17119
rect 12358 17085 12392 17119
rect 12909 17085 12943 17119
rect 13369 17085 13403 17119
rect 13461 17085 13495 17119
rect 13553 17085 13587 17119
rect 14453 17085 14487 17119
rect 14565 17082 14599 17116
rect 14657 17082 14691 17116
rect 14835 17085 14869 17119
rect 14933 17085 14967 17119
rect 16037 17085 16071 17119
rect 16221 17085 16255 17119
rect 16773 17085 16807 17119
rect 17233 17085 17267 17119
rect 17509 17085 17543 17119
rect 17601 17085 17635 17119
rect 18705 17085 18739 17119
rect 21097 17085 21131 17119
rect 23305 17085 23339 17119
rect 24961 17085 24995 17119
rect 28917 17085 28951 17119
rect 30665 17085 30699 17119
rect 31769 17085 31803 17119
rect 11345 17017 11379 17051
rect 11437 17017 11471 17051
rect 12173 17017 12207 17051
rect 17049 17017 17083 17051
rect 17141 17017 17175 17051
rect 18061 17017 18095 17051
rect 20361 17017 20395 17051
rect 22753 17017 22787 17051
rect 23213 17017 23247 17051
rect 27905 17017 27939 17051
rect 29009 17017 29043 17051
rect 9689 16949 9723 16983
rect 10333 16949 10367 16983
rect 12633 16949 12667 16983
rect 12817 16949 12851 16983
rect 13921 16949 13955 16983
rect 14105 16949 14139 16983
rect 15117 16949 15151 16983
rect 15853 16949 15887 16983
rect 16589 16949 16623 16983
rect 17417 16949 17451 16983
rect 18153 16949 18187 16983
rect 21281 16949 21315 16983
rect 25421 16949 25455 16983
rect 26433 16949 26467 16983
rect 8217 16745 8251 16779
rect 8585 16745 8619 16779
rect 8861 16745 8895 16779
rect 9137 16745 9171 16779
rect 11805 16745 11839 16779
rect 14105 16745 14139 16779
rect 15025 16745 15059 16779
rect 15853 16745 15887 16779
rect 16037 16745 16071 16779
rect 17233 16745 17267 16779
rect 18797 16745 18831 16779
rect 22845 16745 22879 16779
rect 27077 16745 27111 16779
rect 27353 16745 27387 16779
rect 31217 16745 31251 16779
rect 14381 16677 14415 16711
rect 20269 16677 20303 16711
rect 29653 16677 29687 16711
rect 5917 16609 5951 16643
rect 8309 16609 8343 16643
rect 8493 16609 8527 16643
rect 8769 16609 8803 16643
rect 9045 16609 9079 16643
rect 10241 16609 10275 16643
rect 10425 16609 10459 16643
rect 10977 16609 11011 16643
rect 11345 16609 11379 16643
rect 12081 16609 12115 16643
rect 12633 16609 12667 16643
rect 13277 16609 13311 16643
rect 13461 16609 13495 16643
rect 13553 16609 13587 16643
rect 13737 16609 13771 16643
rect 14933 16609 14967 16643
rect 15117 16609 15151 16643
rect 15393 16609 15427 16643
rect 15978 16609 16012 16643
rect 16405 16609 16439 16643
rect 16681 16609 16715 16643
rect 17417 16609 17451 16643
rect 17509 16609 17543 16643
rect 18705 16609 18739 16643
rect 19349 16609 19383 16643
rect 20085 16609 20119 16643
rect 22201 16609 22235 16643
rect 26433 16609 26467 16643
rect 27445 16609 27479 16643
rect 10333 16541 10367 16575
rect 11437 16541 11471 16575
rect 12265 16541 12299 16575
rect 12541 16541 12575 16575
rect 15761 16541 15795 16575
rect 16497 16541 16531 16575
rect 18889 16541 18923 16575
rect 19993 16541 20027 16575
rect 29377 16541 29411 16575
rect 31861 16541 31895 16575
rect 6745 16473 6779 16507
rect 13369 16473 13403 16507
rect 14749 16473 14783 16507
rect 17785 16473 17819 16507
rect 5273 16405 5307 16439
rect 14841 16405 14875 16439
rect 17417 16405 17451 16439
rect 18337 16405 18371 16439
rect 31125 16405 31159 16439
rect 11805 16201 11839 16235
rect 13093 16201 13127 16235
rect 13645 16201 13679 16235
rect 14197 16201 14231 16235
rect 15301 16201 15335 16235
rect 15485 16201 15519 16235
rect 17601 16201 17635 16235
rect 19901 16201 19935 16235
rect 22937 16201 22971 16235
rect 31861 16201 31895 16235
rect 8309 16133 8343 16167
rect 12541 16133 12575 16167
rect 13829 16133 13863 16167
rect 14381 16133 14415 16167
rect 17141 16133 17175 16167
rect 22569 16133 22603 16167
rect 6193 16065 6227 16099
rect 8217 16065 8251 16099
rect 9137 16065 9171 16099
rect 12265 16065 12299 16099
rect 14657 16065 14691 16099
rect 18429 16065 18463 16099
rect 23397 16065 23431 16099
rect 24041 16065 24075 16099
rect 29101 16065 29135 16099
rect 4261 15997 4295 16031
rect 4629 15997 4663 16031
rect 6469 15997 6503 16031
rect 6837 15997 6871 16031
rect 7297 15997 7331 16031
rect 8493 15997 8527 16031
rect 8861 15997 8895 16031
rect 11345 15997 11379 16031
rect 11713 15997 11747 16031
rect 11989 15997 12023 16031
rect 12541 15997 12575 16031
rect 12725 15997 12759 16031
rect 15945 15997 15979 16031
rect 16129 15997 16163 16031
rect 16957 15997 16991 16031
rect 17877 15997 17911 16031
rect 18153 15997 18187 16031
rect 24133 15997 24167 16031
rect 26893 15997 26927 16031
rect 29469 15997 29503 16031
rect 30895 15997 30929 16031
rect 31217 15997 31251 16031
rect 3249 15929 3283 15963
rect 5273 15929 5307 15963
rect 8585 15929 8619 15963
rect 8677 15929 8711 15963
rect 14105 15929 14139 15963
rect 14933 15929 14967 15963
rect 15310 15929 15344 15963
rect 17233 15929 17267 15963
rect 17647 15929 17681 15963
rect 6745 15861 6779 15895
rect 7205 15861 7239 15895
rect 7573 15861 7607 15895
rect 11161 15861 11195 15895
rect 11529 15861 11563 15895
rect 22937 15861 22971 15895
rect 23121 15861 23155 15895
rect 24777 15861 24811 15895
rect 26341 15861 26375 15895
rect 3433 15657 3467 15691
rect 12081 15657 12115 15691
rect 17785 15657 17819 15691
rect 19257 15657 19291 15691
rect 19993 15657 20027 15691
rect 23305 15657 23339 15691
rect 30205 15657 30239 15691
rect 4905 15589 4939 15623
rect 6745 15589 6779 15623
rect 7113 15589 7147 15623
rect 13277 15589 13311 15623
rect 13921 15589 13955 15623
rect 19809 15589 19843 15623
rect 21281 15589 21315 15623
rect 31677 15589 31711 15623
rect 11069 15521 11103 15555
rect 11161 15521 11195 15555
rect 11345 15521 11379 15555
rect 12633 15521 12667 15555
rect 12817 15521 12851 15555
rect 12909 15521 12943 15555
rect 13185 15521 13219 15555
rect 13369 15521 13403 15555
rect 14013 15521 14047 15555
rect 14197 15521 14231 15555
rect 14289 15521 14323 15555
rect 14565 15521 14599 15555
rect 14657 15521 14691 15555
rect 15025 15521 15059 15555
rect 15393 15521 15427 15555
rect 15577 15521 15611 15555
rect 15945 15521 15979 15555
rect 16681 15521 16715 15555
rect 17141 15521 17175 15555
rect 19165 15521 19199 15555
rect 21097 15521 21131 15555
rect 21373 15521 21407 15555
rect 24409 15521 24443 15555
rect 24593 15521 24627 15555
rect 24685 15521 24719 15555
rect 25881 15521 25915 15555
rect 27721 15521 27755 15555
rect 30297 15521 30331 15555
rect 30481 15521 30515 15555
rect 5181 15453 5215 15487
rect 7021 15453 7055 15487
rect 7665 15453 7699 15487
rect 9045 15453 9079 15487
rect 11529 15453 11563 15487
rect 17029 15453 17063 15487
rect 17417 15453 17451 15487
rect 17509 15453 17543 15487
rect 20729 15453 20763 15487
rect 20913 15453 20947 15487
rect 21557 15453 21591 15487
rect 21833 15453 21867 15487
rect 23489 15453 23523 15487
rect 24133 15453 24167 15487
rect 24225 15453 24259 15487
rect 26157 15453 26191 15487
rect 14841 15385 14875 15419
rect 19441 15385 19475 15419
rect 27629 15385 27663 15419
rect 5273 15317 5307 15351
rect 8493 15317 8527 15351
rect 10885 15317 10919 15351
rect 11345 15317 11379 15351
rect 12449 15317 12483 15351
rect 14013 15317 14047 15351
rect 16865 15317 16899 15351
rect 19809 15317 19843 15351
rect 20085 15317 20119 15351
rect 27905 15317 27939 15351
rect 6193 15113 6227 15147
rect 8769 15113 8803 15147
rect 11069 15113 11103 15147
rect 12265 15113 12299 15147
rect 15393 15113 15427 15147
rect 16865 15113 16899 15147
rect 17049 15113 17083 15147
rect 23765 15113 23799 15147
rect 27905 15113 27939 15147
rect 31309 15113 31343 15147
rect 11897 15045 11931 15079
rect 12633 15045 12667 15079
rect 29561 15045 29595 15079
rect 4905 14977 4939 15011
rect 5089 14977 5123 15011
rect 5641 14977 5675 15011
rect 6285 14977 6319 15011
rect 7021 14977 7055 15011
rect 10977 14977 11011 15011
rect 17417 14977 17451 15011
rect 18981 14977 19015 15011
rect 19257 14977 19291 15011
rect 20729 14977 20763 15011
rect 21005 14977 21039 15011
rect 22385 14977 22419 15011
rect 23581 14977 23615 15011
rect 26341 14977 26375 15011
rect 27813 14977 27847 15011
rect 29193 14977 29227 15011
rect 30481 14977 30515 15011
rect 3801 14909 3835 14943
rect 5825 14909 5859 14943
rect 11253 14909 11287 14943
rect 11529 14909 11563 14943
rect 11621 14909 11655 14943
rect 11989 14909 12023 14943
rect 13139 14909 13173 14943
rect 13369 14909 13403 14943
rect 14013 14909 14047 14943
rect 14657 14909 14691 14943
rect 14841 14909 14875 14943
rect 15117 14909 15151 14943
rect 15577 14909 15611 14943
rect 15945 14909 15979 14943
rect 16129 14909 16163 14943
rect 16313 14909 16347 14943
rect 16773 14909 16807 14943
rect 17877 14909 17911 14943
rect 18705 14909 18739 14943
rect 21925 14909 21959 14943
rect 22477 14909 22511 14943
rect 22569 14909 22603 14943
rect 24317 14909 24351 14943
rect 25697 14909 25731 14943
rect 26065 14909 26099 14943
rect 28457 14909 28491 14943
rect 29837 14909 29871 14943
rect 30665 14909 30699 14943
rect 31217 14909 31251 14943
rect 4353 14841 4387 14875
rect 4813 14841 4847 14875
rect 7297 14841 7331 14875
rect 12265 14841 12299 14875
rect 17693 14841 17727 14875
rect 21833 14841 21867 14875
rect 25789 14841 25823 14875
rect 30113 14841 30147 14875
rect 4445 14773 4479 14807
rect 5733 14773 5767 14807
rect 6929 14773 6963 14807
rect 9321 14773 9355 14807
rect 11345 14773 11379 14807
rect 12081 14773 12115 14807
rect 13001 14773 13035 14807
rect 17049 14773 17083 14807
rect 17601 14773 17635 14807
rect 17969 14773 18003 14807
rect 18153 14773 18187 14807
rect 21649 14773 21683 14807
rect 22937 14773 22971 14807
rect 23029 14773 23063 14807
rect 24777 14773 24811 14807
rect 28641 14773 28675 14807
rect 29745 14773 29779 14807
rect 29929 14773 29963 14807
rect 6101 14569 6135 14603
rect 6837 14569 6871 14603
rect 8125 14569 8159 14603
rect 8953 14569 8987 14603
rect 10701 14569 10735 14603
rect 11713 14569 11747 14603
rect 15393 14569 15427 14603
rect 17417 14569 17451 14603
rect 18153 14569 18187 14603
rect 20453 14569 20487 14603
rect 23581 14569 23615 14603
rect 27629 14569 27663 14603
rect 28089 14569 28123 14603
rect 31677 14569 31711 14603
rect 5457 14501 5491 14535
rect 7389 14501 7423 14535
rect 11345 14501 11379 14535
rect 20177 14501 20211 14535
rect 21005 14501 21039 14535
rect 21649 14501 21683 14535
rect 23857 14501 23891 14535
rect 28273 14501 28307 14535
rect 28809 14501 28843 14535
rect 29009 14501 29043 14535
rect 30297 14501 30331 14535
rect 5549 14433 5583 14467
rect 6285 14433 6319 14467
rect 6469 14433 6503 14467
rect 6561 14433 6595 14467
rect 6653 14433 6687 14467
rect 8033 14433 8067 14467
rect 8861 14433 8895 14467
rect 9321 14433 9355 14467
rect 10977 14433 11011 14467
rect 11253 14433 11287 14467
rect 11529 14433 11563 14467
rect 11619 14433 11653 14467
rect 11897 14433 11931 14467
rect 11989 14433 12023 14467
rect 12357 14433 12391 14467
rect 12725 14433 12759 14467
rect 13185 14433 13219 14467
rect 13277 14433 13311 14467
rect 13461 14433 13495 14467
rect 14657 14433 14691 14467
rect 14749 14433 14783 14467
rect 15209 14433 15243 14467
rect 15669 14433 15703 14467
rect 16865 14433 16899 14467
rect 17049 14433 17083 14467
rect 17141 14433 17175 14467
rect 17233 14433 17267 14467
rect 18613 14433 18647 14467
rect 20545 14433 20579 14467
rect 20729 14433 20763 14467
rect 21189 14433 21223 14467
rect 23673 14433 23707 14467
rect 23949 14433 23983 14467
rect 24041 14433 24075 14467
rect 25513 14433 25547 14467
rect 27721 14433 27755 14467
rect 28365 14433 28399 14467
rect 30665 14433 30699 14467
rect 31861 14433 31895 14467
rect 4997 14365 5031 14399
rect 5273 14365 5307 14399
rect 9045 14365 9079 14399
rect 9873 14365 9907 14399
rect 12081 14365 12115 14399
rect 12173 14365 12207 14399
rect 13921 14365 13955 14399
rect 15025 14365 15059 14399
rect 15853 14365 15887 14399
rect 15945 14365 15979 14399
rect 17509 14365 17543 14399
rect 19441 14365 19475 14399
rect 21373 14365 21407 14399
rect 25789 14365 25823 14399
rect 27445 14365 27479 14399
rect 29285 14365 29319 14399
rect 31309 14365 31343 14399
rect 7757 14297 7791 14331
rect 15485 14297 15519 14331
rect 18889 14297 18923 14331
rect 23121 14297 23155 14331
rect 27261 14297 27295 14331
rect 30481 14297 30515 14331
rect 3525 14229 3559 14263
rect 8493 14229 8527 14263
rect 10517 14229 10551 14263
rect 10885 14229 10919 14263
rect 11621 14229 11655 14263
rect 13645 14229 13679 14263
rect 14841 14229 14875 14263
rect 16589 14229 16623 14263
rect 18705 14229 18739 14263
rect 20085 14229 20119 14263
rect 24225 14229 24259 14263
rect 25421 14229 25455 14263
rect 28641 14229 28675 14263
rect 28825 14229 28859 14263
rect 29929 14229 29963 14263
rect 30757 14229 30791 14263
rect 5641 14025 5675 14059
rect 6285 14025 6319 14059
rect 6916 14025 6950 14059
rect 11161 14025 11195 14059
rect 13369 14025 13403 14059
rect 14197 14025 14231 14059
rect 14749 14025 14783 14059
rect 15209 14025 15243 14059
rect 17509 14025 17543 14059
rect 19441 14025 19475 14059
rect 25237 14025 25271 14059
rect 26341 14025 26375 14059
rect 27905 14025 27939 14059
rect 29193 14025 29227 14059
rect 31033 14025 31067 14059
rect 8401 13957 8435 13991
rect 10701 13957 10735 13991
rect 13461 13957 13495 13991
rect 15025 13957 15059 13991
rect 20637 13957 20671 13991
rect 26249 13957 26283 13991
rect 28457 13957 28491 13991
rect 3249 13889 3283 13923
rect 6653 13889 6687 13923
rect 8861 13889 8895 13923
rect 10885 13889 10919 13923
rect 11621 13889 11655 13923
rect 15761 13889 15795 13923
rect 16037 13889 16071 13923
rect 17693 13889 17727 13923
rect 17969 13889 18003 13923
rect 22661 13889 22695 13923
rect 26801 13889 26835 13923
rect 26985 13889 27019 13923
rect 27813 13889 27847 13923
rect 28273 13889 28307 13923
rect 29285 13889 29319 13923
rect 29561 13889 29595 13923
rect 4261 13821 4295 13855
rect 9597 13821 9631 13855
rect 9873 13821 9907 13855
rect 10333 13821 10367 13855
rect 10609 13821 10643 13855
rect 11253 13821 11287 13855
rect 14013 13821 14047 13855
rect 14322 13821 14356 13855
rect 14841 13821 14875 13855
rect 15577 13821 15611 13855
rect 20085 13821 20119 13855
rect 20453 13821 20487 13855
rect 20729 13821 20763 13855
rect 21465 13821 21499 13855
rect 22201 13821 22235 13855
rect 22845 13821 22879 13855
rect 23581 13821 23615 13855
rect 25881 13821 25915 13855
rect 26065 13821 26099 13855
rect 26249 13821 26283 13855
rect 26709 13821 26743 13855
rect 28089 13821 28123 13855
rect 28549 13821 28583 13855
rect 28733 13821 28767 13855
rect 28825 13821 28859 13855
rect 29009 13821 29043 13855
rect 31769 13821 31803 13855
rect 11897 13753 11931 13787
rect 15163 13753 15197 13787
rect 24133 13753 24167 13787
rect 24869 13753 24903 13787
rect 31217 13753 31251 13787
rect 9781 13685 9815 13719
rect 11069 13685 11103 13719
rect 11161 13685 11195 13719
rect 14381 13685 14415 13719
rect 19533 13685 19567 13719
rect 20913 13685 20947 13719
rect 21649 13685 21683 13719
rect 23489 13685 23523 13719
rect 27169 13685 27203 13719
rect 7665 13481 7699 13515
rect 10425 13481 10459 13515
rect 14565 13481 14599 13515
rect 15853 13481 15887 13515
rect 16681 13481 16715 13515
rect 18981 13481 19015 13515
rect 21373 13481 21407 13515
rect 23259 13481 23293 13515
rect 24777 13481 24811 13515
rect 24961 13481 24995 13515
rect 25973 13481 26007 13515
rect 26341 13481 26375 13515
rect 31217 13481 31251 13515
rect 31585 13481 31619 13515
rect 12817 13413 12851 13447
rect 14197 13413 14231 13447
rect 15025 13413 15059 13447
rect 19073 13413 19107 13447
rect 19901 13413 19935 13447
rect 31125 13413 31159 13447
rect 4445 13345 4479 13379
rect 7573 13345 7607 13379
rect 10057 13345 10091 13379
rect 10609 13345 10643 13379
rect 12909 13345 12943 13379
rect 13461 13345 13495 13379
rect 14473 13345 14507 13379
rect 14749 13345 14783 13379
rect 16037 13345 16071 13379
rect 16129 13345 16163 13379
rect 16313 13345 16347 13379
rect 16865 13345 16899 13379
rect 23673 13345 23707 13379
rect 24777 13345 24811 13379
rect 25605 13345 25639 13379
rect 27905 13345 27939 13379
rect 28273 13345 28307 13379
rect 28733 13345 28767 13379
rect 29009 13345 29043 13379
rect 31677 13345 31711 13379
rect 3249 13277 3283 13311
rect 9781 13277 9815 13311
rect 10885 13277 10919 13311
rect 12633 13277 12667 13311
rect 16221 13277 16255 13311
rect 17233 13277 17267 13311
rect 19165 13277 19199 13311
rect 19625 13277 19659 13311
rect 21465 13277 21499 13311
rect 21833 13277 21867 13311
rect 26433 13277 26467 13311
rect 26617 13277 26651 13311
rect 27353 13277 27387 13311
rect 27813 13277 27847 13311
rect 29285 13277 29319 13311
rect 30941 13277 30975 13311
rect 31769 13277 31803 13311
rect 14933 13209 14967 13243
rect 15301 13209 15335 13243
rect 8309 13141 8343 13175
rect 15485 13141 15519 13175
rect 18613 13141 18647 13175
rect 26801 13141 26835 13175
rect 28273 13141 28307 13175
rect 28457 13141 28491 13175
rect 28825 13141 28859 13175
rect 30757 13141 30791 13175
rect 6653 12937 6687 12971
rect 7389 12937 7423 12971
rect 10241 12937 10275 12971
rect 11989 12937 12023 12971
rect 12173 12937 12207 12971
rect 15301 12937 15335 12971
rect 16773 12937 16807 12971
rect 17693 12937 17727 12971
rect 20913 12937 20947 12971
rect 21833 12937 21867 12971
rect 24317 12937 24351 12971
rect 26328 12937 26362 12971
rect 27905 12937 27939 12971
rect 29009 12937 29043 12971
rect 30849 12937 30883 12971
rect 12541 12869 12575 12903
rect 17969 12869 18003 12903
rect 8677 12801 8711 12835
rect 10885 12801 10919 12835
rect 13001 12801 13035 12835
rect 15025 12801 15059 12835
rect 18245 12801 18279 12835
rect 21465 12801 21499 12835
rect 22569 12801 22603 12835
rect 26065 12801 26099 12835
rect 28089 12801 28123 12835
rect 28181 12801 28215 12835
rect 29101 12801 29135 12835
rect 31769 12801 31803 12835
rect 6193 12733 6227 12767
rect 7849 12733 7883 12767
rect 7941 12733 7975 12767
rect 9873 12733 9907 12767
rect 17049 12733 17083 12767
rect 17233 12733 17267 12767
rect 17417 12733 17451 12767
rect 18153 12733 18187 12767
rect 21281 12733 21315 12767
rect 22385 12733 22419 12767
rect 25697 12733 25731 12767
rect 28273 12733 28307 12767
rect 28365 12733 28399 12767
rect 28636 12733 28670 12767
rect 9045 12665 9079 12699
rect 12173 12665 12207 12699
rect 12909 12665 12943 12699
rect 14749 12665 14783 12699
rect 17141 12665 17175 12699
rect 18521 12665 18555 12699
rect 21373 12665 21407 12699
rect 22845 12665 22879 12699
rect 28733 12665 28767 12699
rect 28825 12665 28859 12699
rect 29009 12665 29043 12699
rect 29377 12665 29411 12699
rect 5641 12597 5675 12631
rect 7021 12597 7055 12631
rect 8125 12597 8159 12631
rect 16037 12597 16071 12631
rect 16405 12597 16439 12631
rect 16865 12597 16899 12631
rect 19993 12597 20027 12631
rect 25789 12597 25823 12631
rect 27813 12597 27847 12631
rect 31217 12597 31251 12631
rect 5733 12393 5767 12427
rect 6193 12393 6227 12427
rect 9873 12393 9907 12427
rect 13001 12393 13035 12427
rect 18613 12393 18647 12427
rect 20177 12393 20211 12427
rect 22017 12393 22051 12427
rect 22661 12393 22695 12427
rect 22937 12393 22971 12427
rect 24041 12393 24075 12427
rect 24869 12393 24903 12427
rect 26065 12393 26099 12427
rect 27629 12393 27663 12427
rect 5365 12325 5399 12359
rect 6929 12325 6963 12359
rect 10425 12325 10459 12359
rect 11161 12325 11195 12359
rect 12265 12325 12299 12359
rect 14105 12325 14139 12359
rect 14289 12325 14323 12359
rect 16037 12325 16071 12359
rect 21833 12325 21867 12359
rect 23857 12325 23891 12359
rect 25237 12325 25271 12359
rect 25789 12325 25823 12359
rect 26341 12325 26375 12359
rect 6101 12257 6135 12291
rect 6745 12257 6779 12291
rect 6837 12257 6871 12291
rect 7113 12257 7147 12291
rect 8033 12257 8067 12291
rect 10149 12257 10183 12291
rect 16865 12257 16899 12291
rect 19165 12257 19199 12291
rect 20269 12257 20303 12291
rect 22201 12257 22235 12291
rect 22385 12257 22419 12291
rect 22477 12257 22511 12291
rect 22753 12257 22787 12291
rect 22845 12257 22879 12291
rect 23029 12257 23063 12291
rect 23673 12257 23707 12291
rect 24133 12257 24167 12291
rect 25145 12257 25179 12291
rect 25559 12257 25593 12291
rect 25697 12257 25731 12291
rect 25881 12257 25915 12291
rect 27077 12257 27111 12291
rect 27353 12257 27387 12291
rect 27813 12257 27847 12291
rect 29193 12257 29227 12291
rect 29469 12257 29503 12291
rect 29653 12257 29687 12291
rect 29837 12257 29871 12291
rect 30205 12257 30239 12291
rect 30481 12257 30515 12291
rect 31677 12257 31711 12291
rect 3893 12189 3927 12223
rect 5641 12189 5675 12223
rect 6377 12189 6411 12223
rect 7297 12189 7331 12223
rect 7849 12189 7883 12223
rect 8309 12189 8343 12223
rect 10057 12189 10091 12223
rect 10517 12189 10551 12223
rect 10793 12189 10827 12223
rect 13277 12189 13311 12223
rect 16313 12189 16347 12223
rect 17509 12189 17543 12223
rect 19441 12189 19475 12223
rect 25421 12189 25455 12223
rect 29101 12189 29135 12223
rect 6561 12053 6595 12087
rect 9781 12053 9815 12087
rect 12633 12053 12667 12087
rect 16681 12053 16715 12087
rect 17417 12053 17451 12087
rect 18153 12053 18187 12087
rect 19993 12053 20027 12087
rect 23489 12053 23523 12087
rect 29009 12053 29043 12087
rect 4445 11849 4479 11883
rect 6009 11849 6043 11883
rect 8953 11849 8987 11883
rect 14473 11849 14507 11883
rect 14841 11849 14875 11883
rect 20637 11849 20671 11883
rect 27629 11849 27663 11883
rect 30665 11849 30699 11883
rect 31217 11849 31251 11883
rect 11345 11781 11379 11815
rect 15393 11781 15427 11815
rect 16957 11781 16991 11815
rect 19533 11781 19567 11815
rect 24501 11781 24535 11815
rect 30849 11781 30883 11815
rect 4721 11713 4755 11747
rect 8493 11713 8527 11747
rect 9781 11713 9815 11747
rect 11253 11713 11287 11747
rect 18429 11713 18463 11747
rect 18981 11713 19015 11747
rect 19073 11713 19107 11747
rect 21649 11713 21683 11747
rect 27169 11713 27203 11747
rect 28457 11713 28491 11747
rect 29745 11713 29779 11747
rect 31769 11713 31803 11747
rect 4537 11645 4571 11679
rect 5641 11645 5675 11679
rect 5733 11645 5767 11679
rect 6653 11645 6687 11679
rect 10333 11645 10367 11679
rect 11529 11645 11563 11679
rect 11621 11645 11655 11679
rect 11897 11645 11931 11679
rect 12173 11645 12207 11679
rect 12265 11645 12299 11679
rect 13553 11645 13587 11679
rect 14105 11645 14139 11679
rect 14197 11645 14231 11679
rect 15485 11645 15519 11679
rect 15761 11645 15795 11679
rect 18705 11645 18739 11679
rect 20361 11645 20395 11679
rect 20913 11645 20947 11679
rect 24225 11645 24259 11679
rect 24685 11645 24719 11679
rect 24961 11645 24995 11679
rect 25145 11645 25179 11679
rect 25421 11645 25455 11679
rect 25881 11645 25915 11679
rect 26982 11645 27016 11679
rect 27261 11645 27295 11679
rect 27629 11645 27663 11679
rect 28089 11645 28123 11679
rect 28181 11645 28215 11679
rect 28641 11645 28675 11679
rect 8217 11577 8251 11611
rect 11713 11577 11747 11611
rect 25513 11577 25547 11611
rect 25605 11577 25639 11611
rect 25743 11577 25777 11611
rect 26249 11577 26283 11611
rect 27905 11577 27939 11611
rect 28273 11577 28307 11611
rect 30481 11577 30515 11611
rect 30681 11577 30715 11611
rect 5273 11509 5307 11543
rect 5549 11509 5583 11543
rect 5825 11509 5859 11543
rect 6745 11509 6779 11543
rect 9137 11509 9171 11543
rect 10609 11509 10643 11543
rect 12081 11509 12115 11543
rect 12909 11509 12943 11543
rect 13001 11509 13035 11543
rect 16405 11509 16439 11543
rect 16773 11509 16807 11543
rect 19165 11509 19199 11543
rect 19717 11509 19751 11543
rect 25145 11509 25179 11543
rect 25237 11509 25271 11543
rect 27813 11509 27847 11543
rect 29285 11509 29319 11543
rect 30389 11509 30423 11543
rect 6745 11305 6779 11339
rect 7757 11305 7791 11339
rect 8401 11305 8435 11339
rect 8493 11305 8527 11339
rect 11989 11305 12023 11339
rect 12357 11305 12391 11339
rect 12817 11305 12851 11339
rect 17969 11305 18003 11339
rect 21741 11305 21775 11339
rect 28809 11305 28843 11339
rect 30757 11305 30791 11339
rect 30941 11305 30975 11339
rect 31585 11305 31619 11339
rect 5273 11237 5307 11271
rect 10517 11237 10551 11271
rect 13645 11237 13679 11271
rect 17785 11237 17819 11271
rect 19901 11237 19935 11271
rect 29009 11237 29043 11271
rect 29101 11237 29135 11271
rect 4445 11169 4479 11203
rect 4997 11169 5031 11203
rect 7481 11169 7515 11203
rect 7665 11169 7699 11203
rect 9045 11169 9079 11203
rect 9137 11169 9171 11203
rect 9229 11169 9263 11203
rect 9413 11169 9447 11203
rect 9873 11169 9907 11203
rect 10241 11169 10275 11203
rect 12449 11169 12483 11203
rect 13921 11169 13955 11203
rect 14013 11169 14047 11203
rect 14289 11169 14323 11203
rect 16405 11169 16439 11203
rect 18061 11169 18095 11203
rect 20177 11169 20211 11203
rect 21649 11169 21683 11203
rect 22109 11169 22143 11203
rect 22293 11169 22327 11203
rect 24869 11169 24903 11203
rect 26985 11169 27019 11203
rect 29285 11169 29319 11203
rect 30021 11169 30055 11203
rect 30113 11169 30147 11203
rect 30297 11169 30331 11203
rect 30849 11169 30883 11203
rect 31033 11169 31067 11203
rect 31401 11169 31435 11203
rect 31677 11169 31711 11203
rect 3249 11101 3283 11135
rect 8585 11101 8619 11135
rect 9505 11101 9539 11135
rect 9597 11101 9631 11135
rect 9965 11101 9999 11135
rect 12265 11101 12299 11135
rect 14381 11101 14415 11135
rect 15577 11101 15611 11135
rect 17325 11101 17359 11135
rect 21833 11101 21867 11135
rect 22201 11101 22235 11135
rect 25145 11101 25179 11135
rect 26617 11101 26651 11135
rect 26709 11101 26743 11135
rect 28181 11101 28215 11135
rect 13737 11033 13771 11067
rect 14749 11033 14783 11067
rect 18429 11033 18463 11067
rect 21281 11033 21315 11067
rect 29469 11033 29503 11067
rect 30297 11033 30331 11067
rect 8033 10965 8067 10999
rect 8861 10965 8895 10999
rect 10149 10965 10183 10999
rect 16773 10965 16807 10999
rect 27629 10965 27663 10999
rect 28641 10965 28675 10999
rect 28825 10965 28859 10999
rect 31217 10965 31251 10999
rect 8585 10761 8619 10795
rect 18981 10761 19015 10795
rect 20729 10761 20763 10795
rect 23581 10761 23615 10795
rect 23765 10761 23799 10795
rect 25237 10761 25271 10795
rect 26065 10761 26099 10795
rect 29285 10761 29319 10795
rect 30297 10761 30331 10795
rect 6193 10693 6227 10727
rect 14841 10693 14875 10727
rect 18797 10693 18831 10727
rect 23121 10693 23155 10727
rect 29101 10693 29135 10727
rect 5641 10625 5675 10659
rect 5733 10625 5767 10659
rect 6837 10625 6871 10659
rect 8033 10625 8067 10659
rect 10149 10625 10183 10659
rect 10425 10625 10459 10659
rect 12173 10625 12207 10659
rect 12449 10625 12483 10659
rect 13369 10625 13403 10659
rect 16313 10625 16347 10659
rect 16589 10625 16623 10659
rect 18061 10625 18095 10659
rect 18153 10625 18187 10659
rect 25789 10625 25823 10659
rect 27813 10625 27847 10659
rect 4629 10557 4663 10591
rect 12725 10557 12759 10591
rect 13093 10557 13127 10591
rect 15209 10557 15243 10591
rect 15485 10557 15519 10591
rect 18889 10557 18923 10591
rect 21005 10557 21039 10591
rect 22201 10557 22235 10591
rect 22293 10557 22327 10591
rect 23765 10557 23799 10591
rect 23949 10557 23983 10591
rect 24041 10557 24075 10591
rect 24225 10557 24259 10591
rect 28549 10557 28583 10591
rect 29561 10557 29595 10591
rect 30941 10557 30975 10591
rect 31217 10557 31251 10591
rect 5273 10489 5307 10523
rect 5825 10489 5859 10523
rect 21465 10489 21499 10523
rect 23489 10489 23523 10523
rect 27537 10489 27571 10523
rect 27905 10489 27939 10523
rect 29469 10489 29503 10523
rect 31493 10489 31527 10523
rect 6285 10421 6319 10455
rect 8677 10421 8711 10455
rect 10701 10421 10735 10455
rect 12633 10421 12667 10455
rect 15025 10421 15059 10455
rect 15393 10421 15427 10455
rect 21097 10421 21131 10455
rect 22477 10421 22511 10455
rect 23029 10421 23063 10455
rect 24133 10421 24167 10455
rect 29269 10421 29303 10455
rect 30205 10421 30239 10455
rect 6377 10217 6411 10251
rect 9505 10217 9539 10251
rect 10149 10217 10183 10251
rect 10517 10217 10551 10251
rect 12909 10217 12943 10251
rect 14105 10217 14139 10251
rect 14565 10217 14599 10251
rect 16865 10217 16899 10251
rect 18429 10217 18463 10251
rect 18797 10217 18831 10251
rect 20545 10217 20579 10251
rect 22753 10217 22787 10251
rect 24225 10217 24259 10251
rect 25789 10217 25823 10251
rect 26433 10217 26467 10251
rect 27261 10217 27295 10251
rect 29285 10217 29319 10251
rect 31125 10217 31159 10251
rect 5825 10149 5859 10183
rect 9873 10149 9907 10183
rect 16589 10149 16623 10183
rect 17233 10149 17267 10183
rect 22017 10149 22051 10183
rect 23489 10149 23523 10183
rect 24393 10149 24427 10183
rect 24593 10149 24627 10183
rect 27997 10149 28031 10183
rect 29653 10149 29687 10183
rect 31309 10149 31343 10183
rect 3065 10081 3099 10115
rect 10241 10081 10275 10115
rect 14013 10081 14047 10115
rect 16681 10081 16715 10115
rect 18521 10081 18555 10115
rect 19809 10081 19843 10115
rect 25697 10081 25731 10115
rect 26341 10081 26375 10115
rect 26893 10081 26927 10115
rect 26985 10081 27019 10115
rect 27077 10081 27111 10115
rect 27537 10081 27571 10115
rect 28273 10081 28307 10115
rect 28733 10081 28767 10115
rect 28917 10081 28951 10115
rect 29009 10081 29043 10115
rect 29101 10081 29135 10115
rect 31401 10081 31435 10115
rect 31493 10081 31527 10115
rect 31677 10081 31711 10115
rect 6101 10013 6135 10047
rect 14657 10013 14691 10047
rect 14933 10013 14967 10047
rect 16405 10013 16439 10047
rect 17325 10013 17359 10047
rect 17509 10013 17543 10047
rect 22293 10013 22327 10047
rect 22477 10013 22511 10047
rect 22661 10013 22695 10047
rect 24041 10013 24075 10047
rect 26801 10013 26835 10047
rect 27721 10013 27755 10047
rect 28089 10013 28123 10047
rect 29377 10013 29411 10047
rect 23121 9945 23155 9979
rect 3249 9877 3283 9911
rect 4353 9877 4387 9911
rect 17969 9877 18003 9911
rect 19901 9877 19935 9911
rect 24409 9877 24443 9911
rect 27353 9877 27387 9911
rect 28273 9877 28307 9911
rect 28457 9877 28491 9911
rect 31493 9877 31527 9911
rect 14565 9673 14599 9707
rect 14933 9673 14967 9707
rect 15945 9673 15979 9707
rect 21649 9673 21683 9707
rect 25145 9673 25179 9707
rect 27537 9673 27571 9707
rect 28181 9673 28215 9707
rect 29745 9673 29779 9707
rect 14749 9605 14783 9639
rect 21097 9605 21131 9639
rect 22017 9605 22051 9639
rect 22661 9605 22695 9639
rect 25237 9605 25271 9639
rect 28365 9605 28399 9639
rect 29561 9605 29595 9639
rect 8769 9537 8803 9571
rect 15485 9537 15519 9571
rect 16589 9537 16623 9571
rect 20269 9537 20303 9571
rect 20729 9537 20763 9571
rect 25329 9537 25363 9571
rect 27721 9537 27755 9571
rect 27905 9537 27939 9571
rect 29120 9537 29154 9571
rect 14197 9469 14231 9503
rect 16681 9469 16715 9503
rect 18061 9469 18095 9503
rect 19993 9469 20027 9503
rect 20085 9469 20119 9503
rect 20361 9469 20395 9503
rect 21281 9469 21315 9503
rect 21925 9469 21959 9503
rect 22201 9469 22235 9503
rect 22385 9469 22419 9503
rect 23765 9469 23799 9503
rect 24777 9469 24811 9503
rect 25053 9469 25087 9503
rect 25421 9469 25455 9503
rect 25605 9469 25639 9503
rect 25697 9469 25731 9503
rect 25881 9469 25915 9503
rect 26617 9469 26651 9503
rect 26801 9469 26835 9503
rect 27291 9469 27325 9503
rect 27445 9469 27479 9503
rect 27537 9469 27571 9503
rect 27813 9469 27847 9503
rect 28457 9469 28491 9503
rect 28641 9469 28675 9503
rect 28917 9469 28951 9503
rect 29009 9469 29043 9503
rect 29745 9469 29779 9503
rect 30113 9469 30147 9503
rect 30205 9469 30239 9503
rect 30941 9469 30975 9503
rect 31217 9469 31251 9503
rect 18613 9401 18647 9435
rect 21465 9401 21499 9435
rect 22937 9401 22971 9435
rect 23949 9401 23983 9435
rect 24593 9401 24627 9435
rect 25789 9401 25823 9435
rect 26249 9401 26283 9435
rect 26433 9401 26467 9435
rect 26985 9401 27019 9435
rect 27997 9401 28031 9435
rect 29189 9401 29223 9435
rect 8217 9333 8251 9367
rect 14013 9333 14047 9367
rect 14565 9333 14599 9367
rect 17325 9333 17359 9367
rect 18981 9333 19015 9367
rect 19349 9333 19383 9367
rect 21665 9333 21699 9367
rect 21833 9333 21867 9367
rect 22293 9333 22327 9367
rect 24041 9333 24075 9367
rect 24409 9333 24443 9367
rect 24961 9333 24995 9367
rect 25421 9333 25455 9367
rect 26065 9333 26099 9367
rect 27077 9333 27111 9367
rect 28197 9333 28231 9367
rect 28825 9333 28859 9367
rect 30389 9333 30423 9367
rect 31861 9333 31895 9367
rect 6377 9129 6411 9163
rect 10517 9129 10551 9163
rect 12541 9129 12575 9163
rect 16405 9129 16439 9163
rect 17601 9129 17635 9163
rect 23213 9129 23247 9163
rect 25053 9129 25087 9163
rect 26617 9129 26651 9163
rect 27353 9129 27387 9163
rect 27445 9129 27479 9163
rect 27537 9129 27571 9163
rect 27813 9129 27847 9163
rect 31309 9129 31343 9163
rect 13553 9061 13587 9095
rect 14381 9061 14415 9095
rect 19717 9061 19751 9095
rect 28917 9061 28951 9095
rect 29837 9061 29871 9095
rect 10701 8993 10735 9027
rect 10885 8993 10919 9027
rect 14013 8993 14047 9027
rect 18521 8993 18555 9027
rect 19441 8993 19475 9027
rect 21465 8993 21499 9027
rect 24501 8993 24535 9027
rect 24777 8993 24811 9027
rect 25145 8993 25179 9027
rect 25697 8993 25731 9027
rect 25789 8993 25823 9027
rect 25973 8993 26007 9027
rect 26433 8993 26467 9027
rect 27997 8993 28031 9027
rect 29126 8993 29160 9027
rect 31585 8993 31619 9027
rect 31861 8993 31895 9027
rect 11621 8925 11655 8959
rect 11738 8925 11772 8959
rect 11897 8925 11931 8959
rect 14657 8925 14691 8959
rect 14933 8925 14967 8959
rect 17049 8925 17083 8959
rect 17693 8925 17727 8959
rect 17877 8925 17911 8959
rect 19257 8925 19291 8959
rect 21189 8925 21223 8959
rect 21741 8925 21775 8959
rect 23489 8925 23523 8959
rect 24133 8925 24167 8959
rect 24409 8925 24443 8959
rect 24869 8925 24903 8959
rect 25881 8925 25915 8959
rect 28181 8925 28215 8959
rect 28641 8925 28675 8959
rect 29009 8925 29043 8959
rect 29561 8925 29595 8959
rect 11345 8857 11379 8891
rect 24225 8857 24259 8891
rect 27169 8857 27203 8891
rect 31677 8857 31711 8891
rect 12909 8789 12943 8823
rect 13921 8789 13955 8823
rect 14381 8789 14415 8823
rect 14565 8789 14599 8823
rect 16497 8789 16531 8823
rect 17233 8789 17267 8823
rect 18429 8789 18463 8823
rect 18705 8789 18739 8823
rect 26157 8789 26191 8823
rect 27721 8789 27755 8823
rect 29285 8789 29319 8823
rect 31493 8789 31527 8823
rect 12909 8585 12943 8619
rect 14933 8585 14967 8619
rect 17049 8585 17083 8619
rect 18889 8585 18923 8619
rect 21833 8585 21867 8619
rect 27445 8585 27479 8619
rect 27905 8585 27939 8619
rect 28365 8585 28399 8619
rect 29101 8585 29135 8619
rect 30481 8585 30515 8619
rect 31309 8585 31343 8619
rect 6193 8517 6227 8551
rect 14105 8517 14139 8551
rect 21649 8517 21683 8551
rect 24317 8517 24351 8551
rect 29653 8517 29687 8551
rect 30941 8517 30975 8551
rect 5641 8449 5675 8483
rect 6837 8449 6871 8483
rect 13691 8449 13725 8483
rect 14749 8449 14783 8483
rect 16957 8449 16991 8483
rect 18521 8449 18555 8483
rect 19349 8449 19383 8483
rect 19533 8449 19567 8483
rect 22845 8449 22879 8483
rect 23673 8449 23707 8483
rect 26157 8449 26191 8483
rect 27077 8449 27111 8483
rect 27261 8449 27295 8483
rect 29929 8449 29963 8483
rect 5733 8381 5767 8415
rect 13553 8381 13587 8415
rect 13829 8381 13863 8415
rect 14565 8381 14599 8415
rect 15485 8381 15519 8415
rect 15945 8381 15979 8415
rect 16129 8381 16163 8415
rect 16221 8381 16255 8415
rect 18797 8381 18831 8415
rect 21005 8381 21039 8415
rect 21163 8381 21197 8415
rect 21465 8381 21499 8415
rect 21741 8381 21775 8415
rect 21925 8381 21959 8415
rect 22661 8381 22695 8415
rect 23305 8381 23339 8415
rect 23397 8381 23431 8415
rect 24501 8381 24535 8415
rect 25329 8381 25363 8415
rect 25881 8381 25915 8415
rect 26985 8381 27019 8415
rect 27169 8381 27203 8415
rect 27445 8381 27479 8415
rect 27629 8381 27663 8415
rect 27721 8381 27755 8415
rect 28089 8381 28123 8415
rect 28181 8381 28215 8415
rect 28825 8381 28859 8415
rect 29009 8381 29043 8415
rect 29377 8381 29411 8415
rect 30113 8381 30147 8415
rect 30573 8381 30607 8415
rect 30665 8381 30699 8415
rect 30757 8381 30791 8415
rect 30849 8381 30883 8415
rect 31033 8381 31067 8415
rect 31401 8381 31435 8415
rect 5825 8313 5859 8347
rect 16313 8313 16347 8347
rect 21281 8313 21315 8347
rect 21373 8313 21407 8347
rect 23765 8313 23799 8347
rect 24685 8313 24719 8347
rect 28917 8313 28951 8347
rect 6285 8245 6319 8279
rect 12725 8245 12759 8279
rect 15761 8245 15795 8279
rect 19257 8245 19291 8279
rect 19993 8245 20027 8279
rect 22293 8245 22327 8279
rect 22753 8245 22787 8279
rect 23121 8245 23155 8279
rect 25789 8245 25823 8279
rect 26709 8245 26743 8279
rect 26801 8245 26835 8279
rect 28733 8245 28767 8279
rect 29285 8245 29319 8279
rect 29469 8245 29503 8279
rect 30021 8245 30055 8279
rect 31677 8245 31711 8279
rect 18153 8041 18187 8075
rect 18981 8041 19015 8075
rect 22201 8041 22235 8075
rect 22845 8041 22879 8075
rect 25053 8041 25087 8075
rect 28273 8041 28307 8075
rect 31033 8041 31067 8075
rect 6193 7973 6227 8007
rect 16681 7973 16715 8007
rect 21005 7973 21039 8007
rect 21833 7973 21867 8007
rect 21925 7973 21959 8007
rect 26525 7973 26559 8007
rect 3065 7905 3099 7939
rect 6285 7905 6319 7939
rect 14222 7905 14256 7939
rect 15853 7905 15887 7939
rect 16221 7905 16255 7939
rect 18337 7905 18371 7939
rect 19165 7905 19199 7939
rect 20202 7905 20236 7939
rect 20361 7905 20395 7939
rect 21649 7905 21683 7939
rect 22017 7905 22051 7939
rect 22569 7905 22603 7939
rect 22661 7905 22695 7939
rect 22753 7905 22787 7939
rect 22937 7905 22971 7939
rect 23673 7905 23707 7939
rect 24409 7905 24443 7939
rect 28825 7905 28859 7939
rect 28917 7905 28951 7939
rect 29101 7905 29135 7939
rect 29653 7905 29687 7939
rect 30849 7905 30883 7939
rect 31861 7905 31895 7939
rect 5733 7837 5767 7871
rect 6009 7837 6043 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 14105 7837 14139 7871
rect 14381 7837 14415 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 19349 7837 19383 7871
rect 20085 7837 20119 7871
rect 26801 7837 26835 7871
rect 27445 7837 27479 7871
rect 27721 7837 27755 7871
rect 29009 7837 29043 7871
rect 29469 7837 29503 7871
rect 29561 7837 29595 7871
rect 30665 7837 30699 7871
rect 3249 7769 3283 7803
rect 13829 7769 13863 7803
rect 15025 7769 15059 7803
rect 19809 7769 19843 7803
rect 22293 7769 22327 7803
rect 30021 7769 30055 7803
rect 4261 7701 4295 7735
rect 15301 7701 15335 7735
rect 22477 7701 22511 7735
rect 24317 7701 24351 7735
rect 24501 7701 24535 7735
rect 26893 7701 26927 7735
rect 28733 7701 28767 7735
rect 30113 7701 30147 7735
rect 31677 7701 31711 7735
rect 7665 7497 7699 7531
rect 13277 7497 13311 7531
rect 14092 7497 14126 7531
rect 15761 7497 15795 7531
rect 16589 7497 16623 7531
rect 18153 7497 18187 7531
rect 18429 7497 18463 7531
rect 23397 7497 23431 7531
rect 27813 7497 27847 7531
rect 28825 7497 28859 7531
rect 29364 7497 29398 7531
rect 30849 7497 30883 7531
rect 13829 7361 13863 7395
rect 15577 7361 15611 7395
rect 17509 7361 17543 7395
rect 21649 7361 21683 7395
rect 23765 7361 23799 7395
rect 26065 7361 26099 7395
rect 16313 7293 16347 7327
rect 16681 7293 16715 7327
rect 17325 7293 17359 7327
rect 18521 7293 18555 7327
rect 24133 7293 24167 7327
rect 28457 7293 28491 7327
rect 29101 7293 29135 7327
rect 21925 7225 21959 7259
rect 26341 7225 26375 7259
rect 28641 7225 28675 7259
rect 13737 7157 13771 7191
rect 16773 7157 16807 7191
rect 20637 7157 20671 7191
rect 25559 7157 25593 7191
rect 27905 7157 27939 7191
rect 28841 7157 28875 7191
rect 29009 7157 29043 7191
rect 16129 6953 16163 6987
rect 16313 6953 16347 6987
rect 20177 6953 20211 6987
rect 20637 6953 20671 6987
rect 22753 6953 22787 6987
rect 23489 6953 23523 6987
rect 26525 6953 26559 6987
rect 27629 6953 27663 6987
rect 27997 6953 28031 6987
rect 7297 6885 7331 6919
rect 8309 6885 8343 6919
rect 15393 6885 15427 6919
rect 16681 6885 16715 6919
rect 27537 6885 27571 6919
rect 28457 6885 28491 6919
rect 7113 6817 7147 6851
rect 7205 6817 7239 6851
rect 7481 6817 7515 6851
rect 13369 6817 13403 6851
rect 13461 6817 13495 6851
rect 13553 6817 13587 6851
rect 13737 6817 13771 6851
rect 14473 6817 14507 6851
rect 14565 6817 14599 6851
rect 14749 6817 14783 6851
rect 14933 6817 14967 6851
rect 15025 6817 15059 6851
rect 16405 6817 16439 6851
rect 18981 6817 19015 6851
rect 20269 6817 20303 6851
rect 22661 6817 22695 6851
rect 23857 6817 23891 6851
rect 23949 6817 23983 6851
rect 24317 6817 24351 6851
rect 24501 6817 24535 6851
rect 26249 6817 26283 6851
rect 28181 6817 28215 6851
rect 28273 6817 28307 6851
rect 29929 6817 29963 6851
rect 31493 6817 31527 6851
rect 12541 6749 12575 6783
rect 18153 6749 18187 6783
rect 18337 6749 18371 6783
rect 19717 6749 19751 6783
rect 20453 6749 20487 6783
rect 21189 6749 21223 6783
rect 24041 6749 24075 6783
rect 26065 6749 26099 6783
rect 26433 6749 26467 6783
rect 27077 6749 27111 6783
rect 27445 6749 27479 6783
rect 28641 6749 28675 6783
rect 30665 6749 30699 6783
rect 15577 6681 15611 6715
rect 15761 6681 15795 6715
rect 19809 6681 19843 6715
rect 28457 6681 28491 6715
rect 29377 6681 29411 6715
rect 31309 6681 31343 6715
rect 6929 6613 6963 6647
rect 7757 6613 7791 6647
rect 12909 6613 12943 6647
rect 13185 6613 13219 6647
rect 14381 6613 14415 6647
rect 15393 6613 15427 6647
rect 16129 6613 16163 6647
rect 19073 6613 19107 6647
rect 24685 6613 24719 6647
rect 24961 6613 24995 6647
rect 29285 6613 29319 6647
rect 30113 6613 30147 6647
rect 17233 6409 17267 6443
rect 18429 6409 18463 6443
rect 20729 6409 20763 6443
rect 28457 6409 28491 6443
rect 28812 6409 28846 6443
rect 30481 6409 30515 6443
rect 30297 6341 30331 6375
rect 31677 6341 31711 6375
rect 7205 6273 7239 6307
rect 13461 6273 13495 6307
rect 17877 6273 17911 6307
rect 19257 6273 19291 6307
rect 22201 6273 22235 6307
rect 22477 6273 22511 6307
rect 24041 6273 24075 6307
rect 25329 6273 25363 6307
rect 26709 6273 26743 6307
rect 28549 6273 28583 6307
rect 3065 6205 3099 6239
rect 8125 6205 8159 6239
rect 9781 6205 9815 6239
rect 14381 6205 14415 6239
rect 15209 6205 15243 6239
rect 16405 6205 16439 6239
rect 17141 6205 17175 6239
rect 17601 6205 17635 6239
rect 18521 6205 18555 6239
rect 18981 6205 19015 6239
rect 21097 6205 21131 6239
rect 24593 6205 24627 6239
rect 30573 6205 30607 6239
rect 31861 6205 31895 6239
rect 15577 6137 15611 6171
rect 16497 6137 16531 6171
rect 17693 6137 17727 6171
rect 21005 6137 21039 6171
rect 26985 6137 27019 6171
rect 3249 6069 3283 6103
rect 6653 6069 6687 6103
rect 7573 6069 7607 6103
rect 9229 6069 9263 6103
rect 12817 6069 12851 6103
rect 12909 6069 12943 6103
rect 13829 6069 13863 6103
rect 14565 6069 14599 6103
rect 15761 6069 15795 6103
rect 18889 6069 18923 6103
rect 23949 6069 23983 6103
rect 24777 6069 24811 6103
rect 7849 5865 7883 5899
rect 9413 5865 9447 5899
rect 9873 5865 9907 5899
rect 13001 5865 13035 5899
rect 15485 5865 15519 5899
rect 17325 5865 17359 5899
rect 17693 5865 17727 5899
rect 18613 5865 18647 5899
rect 20637 5865 20671 5899
rect 22385 5865 22419 5899
rect 23765 5865 23799 5899
rect 23857 5865 23891 5899
rect 24225 5865 24259 5899
rect 25053 5865 25087 5899
rect 27813 5865 27847 5899
rect 28917 5865 28951 5899
rect 29561 5865 29595 5899
rect 6377 5797 6411 5831
rect 8125 5797 8159 5831
rect 12633 5797 12667 5831
rect 15853 5797 15887 5831
rect 21465 5797 21499 5831
rect 22753 5797 22787 5831
rect 26065 5797 26099 5831
rect 28641 5797 28675 5831
rect 8217 5729 8251 5763
rect 9781 5729 9815 5763
rect 13829 5729 13863 5763
rect 14841 5729 14875 5763
rect 21557 5729 21591 5763
rect 22201 5729 22235 5763
rect 22477 5729 22511 5763
rect 23121 5729 23155 5763
rect 24869 5729 24903 5763
rect 27721 5729 27755 5763
rect 28917 5729 28951 5763
rect 29469 5729 29503 5763
rect 5365 5661 5399 5695
rect 6101 5661 6135 5695
rect 9965 5661 9999 5695
rect 13645 5661 13679 5695
rect 14289 5661 14323 5695
rect 14565 5661 14599 5695
rect 14703 5661 14737 5695
rect 15577 5661 15611 5695
rect 18797 5661 18831 5695
rect 19073 5661 19107 5695
rect 20545 5661 20579 5695
rect 21189 5661 21223 5695
rect 23673 5661 23707 5695
rect 24317 5661 24351 5695
rect 25605 5661 25639 5695
rect 28825 5661 28859 5695
rect 13553 5593 13587 5627
rect 6009 5525 6043 5559
rect 9229 5525 9263 5559
rect 18061 5525 18095 5559
rect 22017 5525 22051 5559
rect 22569 5525 22603 5559
rect 22753 5525 22787 5559
rect 29285 5525 29319 5559
rect 6929 5321 6963 5355
rect 14289 5321 14323 5355
rect 16497 5321 16531 5355
rect 17141 5321 17175 5355
rect 19533 5321 19567 5355
rect 21097 5321 21131 5355
rect 24317 5321 24351 5355
rect 20913 5253 20947 5287
rect 21465 5253 21499 5287
rect 5825 5185 5859 5219
rect 5917 5185 5951 5219
rect 8677 5185 8711 5219
rect 8953 5185 8987 5219
rect 12357 5185 12391 5219
rect 12541 5185 12575 5219
rect 12817 5185 12851 5219
rect 14841 5185 14875 5219
rect 15025 5185 15059 5219
rect 15577 5185 15611 5219
rect 18613 5185 18647 5219
rect 19073 5185 19107 5219
rect 19257 5185 19291 5219
rect 22569 5185 22603 5219
rect 22845 5185 22879 5219
rect 4353 5117 4387 5151
rect 6009 5117 6043 5151
rect 6469 5117 6503 5151
rect 7665 5117 7699 5151
rect 16313 5117 16347 5151
rect 16681 5117 16715 5151
rect 16865 5117 16899 5151
rect 16957 5117 16991 5151
rect 17233 5117 17267 5151
rect 18061 5117 18095 5151
rect 18199 5117 18233 5151
rect 18337 5117 18371 5151
rect 20177 5117 20211 5151
rect 20269 5117 20303 5151
rect 20453 5117 20487 5151
rect 20637 5117 20671 5151
rect 20729 5117 20763 5151
rect 21833 5117 21867 5151
rect 22385 5117 22419 5151
rect 24961 5117 24995 5151
rect 25145 5117 25179 5151
rect 30021 5117 30055 5151
rect 3249 5049 3283 5083
rect 7113 5049 7147 5083
rect 14749 5049 14783 5083
rect 15761 5049 15795 5083
rect 21097 5049 21131 5083
rect 25237 5049 25271 5083
rect 6377 4981 6411 5015
rect 6561 4981 6595 5015
rect 10425 4981 10459 5015
rect 14381 4981 14415 5015
rect 17417 4981 17451 5015
rect 24409 4981 24443 5015
rect 28549 4981 28583 5015
rect 29469 4981 29503 5015
rect 4629 4777 4663 4811
rect 6837 4777 6871 4811
rect 6929 4777 6963 4811
rect 9781 4777 9815 4811
rect 12265 4777 12299 4811
rect 12541 4777 12575 4811
rect 13001 4777 13035 4811
rect 13553 4777 13587 4811
rect 14289 4777 14323 4811
rect 14657 4777 14691 4811
rect 17417 4777 17451 4811
rect 23305 4777 23339 4811
rect 23581 4777 23615 4811
rect 29009 4777 29043 4811
rect 30021 4777 30055 4811
rect 7389 4709 7423 4743
rect 7849 4709 7883 4743
rect 14197 4709 14231 4743
rect 15485 4709 15519 4743
rect 18521 4709 18555 4743
rect 21281 4709 21315 4743
rect 21833 4709 21867 4743
rect 29653 4709 29687 4743
rect 7481 4641 7515 4675
rect 9689 4641 9723 4675
rect 13461 4641 13495 4675
rect 15025 4641 15059 4675
rect 17325 4641 17359 4675
rect 18153 4641 18187 4675
rect 18337 4641 18371 4675
rect 18613 4641 18647 4675
rect 18705 4641 18739 4675
rect 21373 4641 21407 4675
rect 21557 4641 21591 4675
rect 23673 4641 23707 4675
rect 24317 4641 24351 4675
rect 28273 4641 28307 4675
rect 30824 4641 30858 4675
rect 6101 4573 6135 4607
rect 6377 4573 6411 4607
rect 7021 4573 7055 4607
rect 14381 4573 14415 4607
rect 15117 4573 15151 4607
rect 15209 4573 15243 4607
rect 16129 4573 16163 4607
rect 16865 4573 16899 4607
rect 17509 4573 17543 4607
rect 18981 4573 19015 4607
rect 19717 4573 19751 4607
rect 21005 4573 21039 4607
rect 24041 4573 24075 4607
rect 24225 4573 24259 4607
rect 24777 4573 24811 4607
rect 29101 4573 29135 4607
rect 29193 4573 29227 4607
rect 30665 4573 30699 4607
rect 30941 4573 30975 4607
rect 31677 4573 31711 4607
rect 31861 4573 31895 4607
rect 16957 4505 16991 4539
rect 18889 4505 18923 4539
rect 24685 4505 24719 4539
rect 31217 4505 31251 4539
rect 6469 4437 6503 4471
rect 13829 4437 13863 4471
rect 16221 4437 16255 4471
rect 18061 4437 18095 4471
rect 19625 4437 19659 4471
rect 20361 4437 20395 4471
rect 20453 4437 20487 4471
rect 25421 4437 25455 4471
rect 28641 4437 28675 4471
rect 5720 4233 5754 4267
rect 7205 4233 7239 4267
rect 12252 4233 12286 4267
rect 14092 4233 14126 4267
rect 16570 4233 16604 4267
rect 18061 4233 18095 4267
rect 19060 4233 19094 4267
rect 23397 4233 23431 4267
rect 25071 4233 25105 4267
rect 29837 4233 29871 4267
rect 31585 4233 31619 4267
rect 30389 4165 30423 4199
rect 5457 4097 5491 4131
rect 11989 4097 12023 4131
rect 13829 4097 13863 4131
rect 16313 4097 16347 4131
rect 18797 4097 18831 4131
rect 20913 4097 20947 4131
rect 22753 4097 22787 4131
rect 25329 4097 25363 4131
rect 28089 4097 28123 4131
rect 3065 4029 3099 4063
rect 3341 4029 3375 4063
rect 15945 4029 15979 4063
rect 16221 4029 16255 4063
rect 18153 4029 18187 4063
rect 18337 4029 18371 4063
rect 18429 4029 18463 4063
rect 18521 4029 18555 4063
rect 25605 4029 25639 4063
rect 30113 4029 30147 4063
rect 31401 4029 31435 4063
rect 31861 4029 31895 4063
rect 16129 3961 16163 3995
rect 21189 3961 21223 3995
rect 25513 3961 25547 3995
rect 28365 3961 28399 3995
rect 30021 3961 30055 3995
rect 3249 3893 3283 3927
rect 3525 3893 3559 3927
rect 13737 3893 13771 3927
rect 15577 3893 15611 3927
rect 15853 3893 15887 3927
rect 18705 3893 18739 3927
rect 20545 3893 20579 3927
rect 22661 3893 22695 3927
rect 23581 3893 23615 3927
rect 31677 3893 31711 3927
rect 13737 3689 13771 3723
rect 16221 3689 16255 3723
rect 16681 3689 16715 3723
rect 18429 3689 18463 3723
rect 18797 3689 18831 3723
rect 21005 3689 21039 3723
rect 21925 3689 21959 3723
rect 23121 3689 23155 3723
rect 23857 3689 23891 3723
rect 6377 3621 6411 3655
rect 14197 3621 14231 3655
rect 20269 3621 20303 3655
rect 21373 3621 21407 3655
rect 22109 3621 22143 3655
rect 30113 3621 30147 3655
rect 4261 3553 4295 3587
rect 5825 3553 5859 3587
rect 10425 3553 10459 3587
rect 13829 3553 13863 3587
rect 16773 3553 16807 3587
rect 18337 3553 18371 3587
rect 20545 3553 20579 3587
rect 21833 3553 21867 3587
rect 23213 3553 23247 3587
rect 25789 3553 25823 3587
rect 29101 3553 29135 3587
rect 30389 3553 30423 3587
rect 3249 3485 3283 3519
rect 4813 3485 4847 3519
rect 10885 3485 10919 3519
rect 13921 3485 13955 3519
rect 15669 3485 15703 3519
rect 17233 3485 17267 3519
rect 21465 3485 21499 3519
rect 21649 3485 21683 3519
rect 22753 3485 22787 3519
rect 24777 3485 24811 3519
rect 30849 3485 30883 3519
rect 20913 3417 20947 3451
rect 13829 3145 13863 3179
rect 29009 3145 29043 3179
rect 29285 3145 29319 3179
rect 31677 3145 31711 3179
rect 9689 3077 9723 3111
rect 12265 3009 12299 3043
rect 14841 3009 14875 3043
rect 16221 3009 16255 3043
rect 17693 3009 17727 3043
rect 18613 3009 18647 3043
rect 19073 3009 19107 3043
rect 19809 3009 19843 3043
rect 23949 3009 23983 3043
rect 26525 3009 26559 3043
rect 30849 3009 30883 3043
rect 4445 2941 4479 2975
rect 4537 2941 4571 2975
rect 7205 2941 7239 2975
rect 9229 2941 9263 2975
rect 9505 2941 9539 2975
rect 11621 2941 11655 2975
rect 13645 2941 13679 2975
rect 15577 2941 15611 2975
rect 17969 2941 18003 2975
rect 19349 2941 19383 2975
rect 21557 2941 21591 2975
rect 23489 2941 23523 2975
rect 26065 2941 26099 2975
rect 27721 2941 27755 2975
rect 29101 2941 29135 2975
rect 29653 2941 29687 2975
rect 31585 2941 31619 2975
rect 31861 2941 31895 2975
rect 3249 2873 3283 2907
rect 6101 2873 6135 2907
rect 8217 2873 8251 2907
rect 4721 2805 4755 2839
rect 16681 2805 16715 2839
rect 21373 2805 21407 2839
rect 27537 2805 27571 2839
rect 31401 2805 31435 2839
<< metal1 >>
rect 21450 32308 21456 32360
rect 21508 32348 21514 32360
rect 21508 32320 28672 32348
rect 21508 32308 21514 32320
rect 17770 32240 17776 32292
rect 17828 32280 17834 32292
rect 25958 32280 25964 32292
rect 17828 32252 25964 32280
rect 17828 32240 17834 32252
rect 25958 32240 25964 32252
rect 26016 32240 26022 32292
rect 28644 32224 28672 32320
rect 25774 32172 25780 32224
rect 25832 32212 25838 32224
rect 28258 32212 28264 32224
rect 25832 32184 28264 32212
rect 25832 32172 25838 32184
rect 28258 32172 28264 32184
rect 28316 32172 28322 32224
rect 28626 32172 28632 32224
rect 28684 32172 28690 32224
rect 2760 32122 32200 32144
rect 2760 32070 6946 32122
rect 6998 32070 7010 32122
rect 7062 32070 7074 32122
rect 7126 32070 7138 32122
rect 7190 32070 7202 32122
rect 7254 32070 14306 32122
rect 14358 32070 14370 32122
rect 14422 32070 14434 32122
rect 14486 32070 14498 32122
rect 14550 32070 14562 32122
rect 14614 32070 21666 32122
rect 21718 32070 21730 32122
rect 21782 32070 21794 32122
rect 21846 32070 21858 32122
rect 21910 32070 21922 32122
rect 21974 32070 29026 32122
rect 29078 32070 29090 32122
rect 29142 32070 29154 32122
rect 29206 32070 29218 32122
rect 29270 32070 29282 32122
rect 29334 32070 32200 32122
rect 2760 32048 32200 32070
rect 7101 32011 7159 32017
rect 7101 31977 7113 32011
rect 7147 32008 7159 32011
rect 7558 32008 7564 32020
rect 7147 31980 7564 32008
rect 7147 31977 7159 31980
rect 7101 31971 7159 31977
rect 7558 31968 7564 31980
rect 7616 31968 7622 32020
rect 9674 31968 9680 32020
rect 9732 31968 9738 32020
rect 10137 32011 10195 32017
rect 10137 31977 10149 32011
rect 10183 31977 10195 32011
rect 10137 31971 10195 31977
rect 1026 31900 1032 31952
rect 1084 31940 1090 31952
rect 1084 31912 3096 31940
rect 1084 31900 1090 31912
rect 3068 31881 3096 31912
rect 4154 31900 4160 31952
rect 4212 31900 4218 31952
rect 5166 31900 5172 31952
rect 5224 31940 5230 31952
rect 5629 31943 5687 31949
rect 5629 31940 5641 31943
rect 5224 31912 5641 31940
rect 5224 31900 5230 31912
rect 5629 31909 5641 31912
rect 5675 31909 5687 31943
rect 5629 31903 5687 31909
rect 6454 31900 6460 31952
rect 6512 31940 6518 31952
rect 6512 31912 6960 31940
rect 6512 31900 6518 31912
rect 3053 31875 3111 31881
rect 3053 31841 3065 31875
rect 3099 31841 3111 31875
rect 3053 31835 3111 31841
rect 3878 31832 3884 31884
rect 3936 31832 3942 31884
rect 4172 31804 4200 31900
rect 6638 31832 6644 31884
rect 6696 31832 6702 31884
rect 6932 31881 6960 31912
rect 8662 31900 8668 31952
rect 8720 31900 8726 31952
rect 9692 31940 9720 31968
rect 10152 31940 10180 31971
rect 11606 31968 11612 32020
rect 11664 32008 11670 32020
rect 11664 31980 12572 32008
rect 11664 31968 11670 31980
rect 12544 31949 12572 31980
rect 13372 31980 17356 32008
rect 12529 31943 12587 31949
rect 9692 31912 9996 31940
rect 10152 31912 12480 31940
rect 6917 31875 6975 31881
rect 6917 31841 6929 31875
rect 6963 31841 6975 31875
rect 6917 31835 6975 31841
rect 9674 31832 9680 31884
rect 9732 31832 9738 31884
rect 9968 31881 9996 31912
rect 9953 31875 10011 31881
rect 9953 31841 9965 31875
rect 9999 31841 10011 31875
rect 9953 31835 10011 31841
rect 11793 31875 11851 31881
rect 11793 31841 11805 31875
rect 11839 31872 11851 31875
rect 12342 31872 12348 31884
rect 11839 31844 12348 31872
rect 11839 31841 11851 31844
rect 11793 31835 11851 31841
rect 12342 31832 12348 31844
rect 12400 31832 12406 31884
rect 12452 31872 12480 31912
rect 12529 31909 12541 31943
rect 12575 31909 12587 31943
rect 12529 31903 12587 31909
rect 13372 31872 13400 31980
rect 14366 31900 14372 31952
rect 14424 31900 14430 31952
rect 16114 31900 16120 31952
rect 16172 31940 16178 31952
rect 16172 31912 16712 31940
rect 16172 31900 16178 31912
rect 12452 31844 13400 31872
rect 15378 31832 15384 31884
rect 15436 31832 15442 31884
rect 16393 31875 16451 31881
rect 16393 31841 16405 31875
rect 16439 31872 16451 31875
rect 16574 31872 16580 31884
rect 16439 31844 16580 31872
rect 16439 31841 16451 31844
rect 16393 31835 16451 31841
rect 16574 31832 16580 31844
rect 16632 31832 16638 31884
rect 4341 31807 4399 31813
rect 4341 31804 4353 31807
rect 4172 31776 4353 31804
rect 4341 31773 4353 31776
rect 4387 31773 4399 31807
rect 4341 31767 4399 31773
rect 14090 31764 14096 31816
rect 14148 31764 14154 31816
rect 16684 31813 16712 31912
rect 16669 31807 16727 31813
rect 16669 31773 16681 31807
rect 16715 31773 16727 31807
rect 17328 31804 17356 31980
rect 17402 31968 17408 32020
rect 17460 31968 17466 32020
rect 17862 31968 17868 32020
rect 17920 31968 17926 32020
rect 18690 31968 18696 32020
rect 18748 31968 18754 32020
rect 18782 31968 18788 32020
rect 18840 31968 18846 32020
rect 18966 31968 18972 32020
rect 19024 32008 19030 32020
rect 19024 31980 20944 32008
rect 19024 31968 19030 31980
rect 17420 31872 17448 31968
rect 17681 31875 17739 31881
rect 17681 31872 17693 31875
rect 17420 31844 17693 31872
rect 17681 31841 17693 31844
rect 17727 31841 17739 31875
rect 18708 31872 18736 31968
rect 20622 31900 20628 31952
rect 20680 31900 20686 31952
rect 18969 31875 19027 31881
rect 18969 31872 18981 31875
rect 18708 31844 18981 31872
rect 17681 31835 17739 31841
rect 18969 31841 18981 31844
rect 19015 31841 19027 31875
rect 18969 31835 19027 31841
rect 20640 31804 20668 31900
rect 20916 31881 20944 31980
rect 22002 31968 22008 32020
rect 22060 31968 22066 32020
rect 25774 31968 25780 32020
rect 25832 31968 25838 32020
rect 31018 31968 31024 32020
rect 31076 32008 31082 32020
rect 31665 32011 31723 32017
rect 31665 32008 31677 32011
rect 31076 31980 31677 32008
rect 31076 31968 31082 31980
rect 31665 31977 31677 31980
rect 31711 31977 31723 32011
rect 31665 31971 31723 31977
rect 33134 31968 33140 32020
rect 33192 31968 33198 32020
rect 20901 31875 20959 31881
rect 20901 31841 20913 31875
rect 20947 31841 20959 31875
rect 22020 31872 22048 31968
rect 23842 31900 23848 31952
rect 23900 31940 23906 31952
rect 23900 31912 24440 31940
rect 23900 31900 23906 31912
rect 22557 31875 22615 31881
rect 22557 31872 22569 31875
rect 22020 31844 22569 31872
rect 20901 31835 20959 31841
rect 22557 31841 22569 31844
rect 22603 31841 22615 31875
rect 22557 31835 22615 31841
rect 24026 31832 24032 31884
rect 24084 31832 24090 31884
rect 24412 31813 24440 31912
rect 25130 31900 25136 31952
rect 25188 31900 25194 31952
rect 21361 31807 21419 31813
rect 21361 31804 21373 31807
rect 17328 31776 18460 31804
rect 20640 31776 21373 31804
rect 16669 31767 16727 31773
rect 18432 31680 18460 31776
rect 21361 31773 21373 31776
rect 21407 31773 21419 31807
rect 21361 31767 21419 31773
rect 24397 31807 24455 31813
rect 24397 31773 24409 31807
rect 24443 31773 24455 31807
rect 25148 31804 25176 31900
rect 25498 31832 25504 31884
rect 25556 31832 25562 31884
rect 25593 31875 25651 31881
rect 25593 31841 25605 31875
rect 25639 31872 25651 31875
rect 25685 31875 25743 31881
rect 25685 31872 25697 31875
rect 25639 31844 25697 31872
rect 25639 31841 25651 31844
rect 25593 31835 25651 31841
rect 25685 31841 25697 31844
rect 25731 31872 25743 31875
rect 25792 31872 25820 31968
rect 25731 31844 25820 31872
rect 25884 31912 26280 31940
rect 25731 31841 25743 31844
rect 25685 31835 25743 31841
rect 25884 31804 25912 31912
rect 26252 31881 26280 31912
rect 26418 31900 26424 31952
rect 26476 31940 26482 31952
rect 26476 31912 27016 31940
rect 26476 31900 26482 31912
rect 26237 31875 26295 31881
rect 26237 31841 26249 31875
rect 26283 31841 26295 31875
rect 26237 31835 26295 31841
rect 26513 31875 26571 31881
rect 26513 31841 26525 31875
rect 26559 31841 26571 31875
rect 26513 31835 26571 31841
rect 25148 31776 25912 31804
rect 24397 31767 24455 31773
rect 25958 31764 25964 31816
rect 26016 31804 26022 31816
rect 26528 31804 26556 31835
rect 26988 31813 27016 31912
rect 28074 31900 28080 31952
rect 28132 31940 28138 31952
rect 28132 31912 30420 31940
rect 28132 31900 28138 31912
rect 28626 31832 28632 31884
rect 28684 31832 28690 31884
rect 28718 31832 28724 31884
rect 28776 31872 28782 31884
rect 30392 31881 30420 31912
rect 30101 31875 30159 31881
rect 30101 31872 30113 31875
rect 28776 31844 30113 31872
rect 28776 31832 28782 31844
rect 30101 31841 30113 31844
rect 30147 31841 30159 31875
rect 30101 31835 30159 31841
rect 30377 31875 30435 31881
rect 30377 31841 30389 31875
rect 30423 31841 30435 31875
rect 30377 31835 30435 31841
rect 31849 31875 31907 31881
rect 31849 31841 31861 31875
rect 31895 31872 31907 31875
rect 33152 31872 33180 31968
rect 31895 31844 33180 31872
rect 31895 31841 31907 31844
rect 31849 31835 31907 31841
rect 26016 31776 26556 31804
rect 26973 31807 27031 31813
rect 26016 31764 26022 31776
rect 26973 31773 26985 31807
rect 27019 31773 27031 31807
rect 26973 31767 27031 31773
rect 28350 31764 28356 31816
rect 28408 31804 28414 31816
rect 29089 31807 29147 31813
rect 29089 31804 29101 31807
rect 28408 31776 29101 31804
rect 28408 31764 28414 31776
rect 29089 31773 29101 31776
rect 29135 31773 29147 31807
rect 29089 31767 29147 31773
rect 19518 31696 19524 31748
rect 19576 31736 19582 31748
rect 26053 31739 26111 31745
rect 26053 31736 26065 31739
rect 19576 31708 26065 31736
rect 19576 31696 19582 31708
rect 26053 31705 26065 31708
rect 26099 31705 26111 31739
rect 26053 31699 26111 31705
rect 3237 31671 3295 31677
rect 3237 31637 3249 31671
rect 3283 31668 3295 31671
rect 11882 31668 11888 31680
rect 3283 31640 11888 31668
rect 3283 31637 3295 31640
rect 3237 31631 3295 31637
rect 11882 31628 11888 31640
rect 11940 31628 11946 31680
rect 18414 31628 18420 31680
rect 18472 31628 18478 31680
rect 22370 31628 22376 31680
rect 22428 31628 22434 31680
rect 25777 31671 25835 31677
rect 25777 31637 25789 31671
rect 25823 31668 25835 31671
rect 25958 31668 25964 31680
rect 25823 31640 25964 31668
rect 25823 31637 25835 31640
rect 25777 31631 25835 31637
rect 25958 31628 25964 31640
rect 26016 31628 26022 31680
rect 2760 31578 32200 31600
rect 2760 31526 6286 31578
rect 6338 31526 6350 31578
rect 6402 31526 6414 31578
rect 6466 31526 6478 31578
rect 6530 31526 6542 31578
rect 6594 31526 13646 31578
rect 13698 31526 13710 31578
rect 13762 31526 13774 31578
rect 13826 31526 13838 31578
rect 13890 31526 13902 31578
rect 13954 31526 21006 31578
rect 21058 31526 21070 31578
rect 21122 31526 21134 31578
rect 21186 31526 21198 31578
rect 21250 31526 21262 31578
rect 21314 31526 28366 31578
rect 28418 31526 28430 31578
rect 28482 31526 28494 31578
rect 28546 31526 28558 31578
rect 28610 31526 28622 31578
rect 28674 31526 32200 31578
rect 2760 31504 32200 31526
rect 15010 31424 15016 31476
rect 15068 31464 15074 31476
rect 15068 31436 28212 31464
rect 15068 31424 15074 31436
rect 11701 31399 11759 31405
rect 11701 31365 11713 31399
rect 11747 31396 11759 31399
rect 11747 31368 12388 31396
rect 11747 31365 11759 31368
rect 11701 31359 11759 31365
rect 2314 31288 2320 31340
rect 2372 31328 2378 31340
rect 12360 31337 12388 31368
rect 23658 31356 23664 31408
rect 23716 31396 23722 31408
rect 24578 31396 24584 31408
rect 23716 31368 24584 31396
rect 23716 31356 23722 31368
rect 24578 31356 24584 31368
rect 24636 31356 24642 31408
rect 24946 31356 24952 31408
rect 25004 31396 25010 31408
rect 25866 31396 25872 31408
rect 25004 31368 25872 31396
rect 25004 31356 25010 31368
rect 3237 31331 3295 31337
rect 3237 31328 3249 31331
rect 2372 31300 3249 31328
rect 2372 31288 2378 31300
rect 3237 31297 3249 31300
rect 3283 31297 3295 31331
rect 11057 31331 11115 31337
rect 11057 31328 11069 31331
rect 3237 31291 3295 31297
rect 10796 31300 11069 31328
rect 4154 31220 4160 31272
rect 4212 31260 4218 31272
rect 4249 31263 4307 31269
rect 4249 31260 4261 31263
rect 4212 31232 4261 31260
rect 4212 31220 4218 31232
rect 4249 31229 4261 31232
rect 4295 31229 4307 31263
rect 4249 31223 4307 31229
rect 10796 31136 10824 31300
rect 11057 31297 11069 31300
rect 11103 31297 11115 31331
rect 11057 31291 11115 31297
rect 12345 31331 12403 31337
rect 12345 31297 12357 31331
rect 12391 31297 12403 31331
rect 12345 31291 12403 31297
rect 12894 31288 12900 31340
rect 12952 31328 12958 31340
rect 13449 31331 13507 31337
rect 13449 31328 13461 31331
rect 12952 31300 13461 31328
rect 12952 31288 12958 31300
rect 13449 31297 13461 31300
rect 13495 31297 13507 31331
rect 13449 31291 13507 31297
rect 14182 31288 14188 31340
rect 14240 31328 14246 31340
rect 14550 31328 14556 31340
rect 14240 31300 14556 31328
rect 14240 31288 14246 31300
rect 14550 31288 14556 31300
rect 14608 31288 14614 31340
rect 24486 31328 24492 31340
rect 23492 31300 24492 31328
rect 11333 31263 11391 31269
rect 11333 31229 11345 31263
rect 11379 31260 11391 31263
rect 12434 31260 12440 31272
rect 11379 31232 12440 31260
rect 11379 31229 11391 31232
rect 11333 31223 11391 31229
rect 12434 31220 12440 31232
rect 12492 31260 12498 31272
rect 12989 31263 13047 31269
rect 12989 31260 13001 31263
rect 12492 31232 13001 31260
rect 12492 31220 12498 31232
rect 12989 31229 13001 31232
rect 13035 31229 13047 31263
rect 12989 31223 13047 31229
rect 15381 31263 15439 31269
rect 15381 31229 15393 31263
rect 15427 31260 15439 31263
rect 15427 31232 15976 31260
rect 15427 31229 15439 31232
rect 15381 31223 15439 31229
rect 15948 31136 15976 31232
rect 16574 31220 16580 31272
rect 16632 31220 16638 31272
rect 18046 31220 18052 31272
rect 18104 31220 18110 31272
rect 21269 31263 21327 31269
rect 21269 31229 21281 31263
rect 21315 31260 21327 31263
rect 22094 31260 22100 31272
rect 21315 31232 22100 31260
rect 21315 31229 21327 31232
rect 21269 31223 21327 31229
rect 22094 31220 22100 31232
rect 22152 31220 22158 31272
rect 23106 31220 23112 31272
rect 23164 31260 23170 31272
rect 23492 31269 23520 31300
rect 24486 31288 24492 31300
rect 24544 31288 24550 31340
rect 23477 31263 23535 31269
rect 23477 31260 23489 31263
rect 23164 31232 23489 31260
rect 23164 31220 23170 31232
rect 23477 31229 23489 31232
rect 23523 31229 23535 31263
rect 23477 31223 23535 31229
rect 23750 31220 23756 31272
rect 23808 31220 23814 31272
rect 24026 31220 24032 31272
rect 24084 31260 24090 31272
rect 24121 31263 24179 31269
rect 24121 31260 24133 31263
rect 24084 31232 24133 31260
rect 24084 31220 24090 31232
rect 24121 31229 24133 31232
rect 24167 31229 24179 31263
rect 24121 31223 24179 31229
rect 24578 31220 24584 31272
rect 24636 31220 24642 31272
rect 24670 31220 24676 31272
rect 24728 31262 24734 31272
rect 25056 31269 25084 31368
rect 25866 31356 25872 31368
rect 25924 31356 25930 31408
rect 26326 31356 26332 31408
rect 26384 31396 26390 31408
rect 27525 31399 27583 31405
rect 27525 31396 27537 31399
rect 26384 31368 27537 31396
rect 26384 31356 26390 31368
rect 27525 31365 27537 31368
rect 27571 31365 27583 31399
rect 27525 31359 27583 31365
rect 25608 31300 25820 31328
rect 24857 31263 24915 31269
rect 24857 31262 24869 31263
rect 24728 31234 24869 31262
rect 24728 31220 24734 31234
rect 24857 31229 24869 31234
rect 24903 31229 24915 31263
rect 24857 31223 24915 31229
rect 25041 31263 25099 31269
rect 25041 31229 25053 31263
rect 25087 31229 25099 31263
rect 25041 31223 25099 31229
rect 25130 31220 25136 31272
rect 25188 31260 25194 31272
rect 25225 31263 25283 31269
rect 25225 31260 25237 31263
rect 25188 31232 25237 31260
rect 25188 31220 25194 31232
rect 25225 31229 25237 31232
rect 25271 31229 25283 31263
rect 25225 31223 25283 31229
rect 25383 31263 25441 31269
rect 25383 31229 25395 31263
rect 25429 31262 25441 31263
rect 25429 31260 25544 31262
rect 25608 31260 25636 31300
rect 25429 31234 25636 31260
rect 25429 31229 25452 31234
rect 25516 31232 25636 31234
rect 25383 31223 25452 31229
rect 24302 31201 24308 31204
rect 24279 31195 24308 31201
rect 24279 31161 24291 31195
rect 24279 31155 24308 31161
rect 24302 31152 24308 31155
rect 24360 31152 24366 31204
rect 24394 31152 24400 31204
rect 24452 31152 24458 31204
rect 24486 31152 24492 31204
rect 24544 31152 24550 31204
rect 24949 31195 25007 31201
rect 24949 31161 24961 31195
rect 24995 31161 25007 31195
rect 24949 31155 25007 31161
rect 10778 31084 10784 31136
rect 10836 31084 10842 31136
rect 11241 31127 11299 31133
rect 11241 31093 11253 31127
rect 11287 31124 11299 31127
rect 11330 31124 11336 31136
rect 11287 31096 11336 31124
rect 11287 31093 11299 31096
rect 11241 31087 11299 31093
rect 11330 31084 11336 31096
rect 11388 31084 11394 31136
rect 11790 31084 11796 31136
rect 11848 31084 11854 31136
rect 15102 31084 15108 31136
rect 15160 31084 15166 31136
rect 15286 31084 15292 31136
rect 15344 31084 15350 31136
rect 15930 31084 15936 31136
rect 15988 31084 15994 31136
rect 16022 31084 16028 31136
rect 16080 31084 16086 31136
rect 17494 31084 17500 31136
rect 17552 31084 17558 31136
rect 18509 31127 18567 31133
rect 18509 31093 18521 31127
rect 18555 31124 18567 31127
rect 18598 31124 18604 31136
rect 18555 31096 18604 31124
rect 18555 31093 18567 31096
rect 18509 31087 18567 31093
rect 18598 31084 18604 31096
rect 18656 31084 18662 31136
rect 21358 31084 21364 31136
rect 21416 31084 21422 31136
rect 23569 31127 23627 31133
rect 23569 31093 23581 31127
rect 23615 31124 23627 31127
rect 23658 31124 23664 31136
rect 23615 31096 23664 31124
rect 23615 31093 23627 31096
rect 23569 31087 23627 31093
rect 23658 31084 23664 31096
rect 23716 31084 23722 31136
rect 23934 31084 23940 31136
rect 23992 31084 23998 31136
rect 24762 31084 24768 31136
rect 24820 31084 24826 31136
rect 24964 31124 24992 31155
rect 25222 31124 25228 31136
rect 24964 31096 25228 31124
rect 25222 31084 25228 31096
rect 25280 31084 25286 31136
rect 25314 31084 25320 31136
rect 25372 31124 25378 31136
rect 25424 31124 25452 31223
rect 25682 31220 25688 31272
rect 25740 31220 25746 31272
rect 25792 31260 25820 31300
rect 26050 31288 26056 31340
rect 26108 31288 26114 31340
rect 26191 31263 26249 31269
rect 25792 31256 26096 31260
rect 26191 31256 26203 31263
rect 25792 31232 26203 31256
rect 26068 31229 26203 31232
rect 26237 31260 26249 31263
rect 26237 31229 26254 31260
rect 26068 31228 26254 31229
rect 26191 31223 26249 31228
rect 26326 31220 26332 31272
rect 26384 31220 26390 31272
rect 26418 31220 26424 31272
rect 26476 31220 26482 31272
rect 26513 31263 26571 31269
rect 26513 31229 26525 31263
rect 26559 31260 26571 31263
rect 26559 31232 26648 31260
rect 26559 31229 26571 31232
rect 26513 31223 26571 31229
rect 25501 31195 25559 31201
rect 25501 31161 25513 31195
rect 25547 31161 25559 31195
rect 25501 31155 25559 31161
rect 25372 31096 25452 31124
rect 25516 31124 25544 31155
rect 25590 31152 25596 31204
rect 25648 31152 25654 31204
rect 26620 31136 26648 31232
rect 26878 31220 26884 31272
rect 26936 31220 26942 31272
rect 28184 31269 28212 31436
rect 30098 31288 30104 31340
rect 30156 31288 30162 31340
rect 34146 31288 34152 31340
rect 34204 31288 34210 31340
rect 27433 31263 27491 31269
rect 27433 31229 27445 31263
rect 27479 31260 27491 31263
rect 27709 31263 27767 31269
rect 27709 31260 27721 31263
rect 27479 31232 27721 31260
rect 27479 31229 27491 31232
rect 27433 31223 27491 31229
rect 27709 31229 27721 31232
rect 27755 31229 27767 31263
rect 27709 31223 27767 31229
rect 28169 31263 28227 31269
rect 28169 31229 28181 31263
rect 28215 31229 28227 31263
rect 28169 31223 28227 31229
rect 29638 31220 29644 31272
rect 29696 31220 29702 31272
rect 29365 31195 29423 31201
rect 29365 31161 29377 31195
rect 29411 31192 29423 31195
rect 34164 31192 34192 31288
rect 29411 31164 34192 31192
rect 29411 31161 29423 31164
rect 29365 31155 29423 31161
rect 25774 31124 25780 31136
rect 25516 31096 25780 31124
rect 25372 31084 25378 31096
rect 25774 31084 25780 31096
rect 25832 31084 25838 31136
rect 25869 31127 25927 31133
rect 25869 31093 25881 31127
rect 25915 31124 25927 31127
rect 26510 31124 26516 31136
rect 25915 31096 26516 31124
rect 25915 31093 25927 31096
rect 25869 31087 25927 31093
rect 26510 31084 26516 31096
rect 26568 31084 26574 31136
rect 26602 31084 26608 31136
rect 26660 31084 26666 31136
rect 26697 31127 26755 31133
rect 26697 31093 26709 31127
rect 26743 31124 26755 31127
rect 27154 31124 27160 31136
rect 26743 31096 27160 31124
rect 26743 31093 26755 31096
rect 26697 31087 26755 31093
rect 27154 31084 27160 31096
rect 27212 31084 27218 31136
rect 2760 31034 32200 31056
rect 2760 30982 6946 31034
rect 6998 30982 7010 31034
rect 7062 30982 7074 31034
rect 7126 30982 7138 31034
rect 7190 30982 7202 31034
rect 7254 30982 14306 31034
rect 14358 30982 14370 31034
rect 14422 30982 14434 31034
rect 14486 30982 14498 31034
rect 14550 30982 14562 31034
rect 14614 30982 21666 31034
rect 21718 30982 21730 31034
rect 21782 30982 21794 31034
rect 21846 30982 21858 31034
rect 21910 30982 21922 31034
rect 21974 30982 29026 31034
rect 29078 30982 29090 31034
rect 29142 30982 29154 31034
rect 29206 30982 29218 31034
rect 29270 30982 29282 31034
rect 29334 30982 32200 31034
rect 2760 30960 32200 30982
rect 11790 30920 11796 30932
rect 10888 30892 11796 30920
rect 10888 30861 10916 30892
rect 11790 30880 11796 30892
rect 11848 30880 11854 30932
rect 11882 30880 11888 30932
rect 11940 30920 11946 30932
rect 22370 30920 22376 30932
rect 11940 30892 18552 30920
rect 11940 30880 11946 30892
rect 10873 30855 10931 30861
rect 10873 30821 10885 30855
rect 10919 30821 10931 30855
rect 12529 30855 12587 30861
rect 12529 30852 12541 30855
rect 12098 30824 12541 30852
rect 10873 30815 10931 30821
rect 12529 30821 12541 30824
rect 12575 30821 12587 30855
rect 15286 30852 15292 30864
rect 14766 30824 15292 30852
rect 12529 30815 12587 30821
rect 15286 30812 15292 30824
rect 15344 30812 15350 30864
rect 15933 30855 15991 30861
rect 15933 30821 15945 30855
rect 15979 30852 15991 30855
rect 16022 30852 16028 30864
rect 15979 30824 16028 30852
rect 15979 30821 15991 30824
rect 15933 30815 15991 30821
rect 16022 30812 16028 30824
rect 16080 30812 16086 30864
rect 16942 30812 16948 30864
rect 17000 30812 17006 30864
rect 4430 30744 4436 30796
rect 4488 30744 4494 30796
rect 4522 30744 4528 30796
rect 4580 30744 4586 30796
rect 12434 30784 12440 30796
rect 12360 30756 12440 30784
rect 1302 30676 1308 30728
rect 1360 30716 1366 30728
rect 3237 30719 3295 30725
rect 3237 30716 3249 30719
rect 1360 30688 3249 30716
rect 1360 30676 1366 30688
rect 3237 30685 3249 30688
rect 3283 30685 3295 30719
rect 3237 30679 3295 30685
rect 4801 30719 4859 30725
rect 4801 30685 4813 30719
rect 4847 30716 4859 30719
rect 5350 30716 5356 30728
rect 4847 30688 5356 30716
rect 4847 30685 4859 30688
rect 4801 30679 4859 30685
rect 5350 30676 5356 30688
rect 5408 30676 5414 30728
rect 10597 30719 10655 30725
rect 10597 30685 10609 30719
rect 10643 30716 10655 30719
rect 10870 30716 10876 30728
rect 10643 30688 10876 30716
rect 10643 30685 10655 30688
rect 10597 30679 10655 30685
rect 10870 30676 10876 30688
rect 10928 30676 10934 30728
rect 12360 30725 12388 30756
rect 12434 30744 12440 30756
rect 12492 30744 12498 30796
rect 12618 30744 12624 30796
rect 12676 30784 12682 30796
rect 12805 30787 12863 30793
rect 12805 30784 12817 30787
rect 12676 30756 12817 30784
rect 12676 30744 12682 30756
rect 12805 30753 12817 30756
rect 12851 30753 12863 30787
rect 12805 30747 12863 30753
rect 12345 30719 12403 30725
rect 12345 30685 12357 30719
rect 12391 30685 12403 30719
rect 12345 30679 12403 30685
rect 13265 30719 13323 30725
rect 13265 30685 13277 30719
rect 13311 30685 13323 30719
rect 13265 30679 13323 30685
rect 12894 30540 12900 30592
rect 12952 30540 12958 30592
rect 13280 30580 13308 30679
rect 13538 30676 13544 30728
rect 13596 30676 13602 30728
rect 15657 30719 15715 30725
rect 15657 30716 15669 30719
rect 14936 30688 15669 30716
rect 14274 30580 14280 30592
rect 13280 30552 14280 30580
rect 14274 30540 14280 30552
rect 14332 30580 14338 30592
rect 14936 30580 14964 30688
rect 15657 30685 15669 30688
rect 15703 30716 15715 30719
rect 15703 30688 17080 30716
rect 15703 30685 15715 30688
rect 15657 30679 15715 30685
rect 15010 30608 15016 30660
rect 15068 30608 15074 30660
rect 17052 30592 17080 30688
rect 18414 30676 18420 30728
rect 18472 30676 18478 30728
rect 18524 30716 18552 30892
rect 18616 30892 22376 30920
rect 18616 30793 18644 30892
rect 22370 30880 22376 30892
rect 22428 30880 22434 30932
rect 23750 30880 23756 30932
rect 23808 30920 23814 30932
rect 24029 30923 24087 30929
rect 24029 30920 24041 30923
rect 23808 30892 24041 30920
rect 23808 30880 23814 30892
rect 24029 30889 24041 30892
rect 24075 30889 24087 30923
rect 24029 30883 24087 30889
rect 24578 30880 24584 30932
rect 24636 30920 24642 30932
rect 24946 30920 24952 30932
rect 24636 30892 24952 30920
rect 24636 30880 24642 30892
rect 24946 30880 24952 30892
rect 25004 30880 25010 30932
rect 25130 30880 25136 30932
rect 25188 30880 25194 30932
rect 25682 30880 25688 30932
rect 25740 30880 25746 30932
rect 26418 30880 26424 30932
rect 26476 30880 26482 30932
rect 27614 30920 27620 30932
rect 26528 30892 27620 30920
rect 21358 30812 21364 30864
rect 21416 30812 21422 30864
rect 24302 30812 24308 30864
rect 24360 30852 24366 30864
rect 24670 30852 24676 30864
rect 24360 30824 24676 30852
rect 24360 30812 24366 30824
rect 24670 30812 24676 30824
rect 24728 30852 24734 30864
rect 25038 30852 25044 30864
rect 24728 30824 25044 30852
rect 24728 30812 24734 30824
rect 25038 30812 25044 30824
rect 25096 30812 25102 30864
rect 25148 30852 25176 30880
rect 25148 30824 25636 30852
rect 19518 30793 19524 30796
rect 18601 30787 18659 30793
rect 18601 30753 18613 30787
rect 18647 30753 18659 30787
rect 18601 30747 18659 30753
rect 19337 30787 19395 30793
rect 19337 30753 19349 30787
rect 19383 30753 19395 30787
rect 19337 30747 19395 30753
rect 19475 30787 19524 30793
rect 19475 30753 19487 30787
rect 19521 30753 19524 30787
rect 19475 30747 19524 30753
rect 19352 30716 19380 30747
rect 19518 30744 19524 30747
rect 19576 30744 19582 30796
rect 23842 30744 23848 30796
rect 23900 30744 23906 30796
rect 24026 30744 24032 30796
rect 24084 30744 24090 30796
rect 24762 30744 24768 30796
rect 24820 30784 24826 30796
rect 25133 30787 25191 30793
rect 25133 30784 25145 30787
rect 24820 30756 25145 30784
rect 24820 30744 24826 30756
rect 25133 30753 25145 30756
rect 25179 30753 25191 30787
rect 25133 30747 25191 30753
rect 25314 30744 25320 30796
rect 25372 30744 25378 30796
rect 18524 30688 19380 30716
rect 19613 30719 19671 30725
rect 19613 30685 19625 30719
rect 19659 30716 19671 30719
rect 19659 30688 20024 30716
rect 19659 30685 19671 30688
rect 19613 30679 19671 30685
rect 17310 30608 17316 30660
rect 17368 30648 17374 30660
rect 17405 30651 17463 30657
rect 17405 30648 17417 30651
rect 17368 30620 17417 30648
rect 17368 30608 17374 30620
rect 17405 30617 17417 30620
rect 17451 30648 17463 30651
rect 17770 30648 17776 30660
rect 17451 30620 17776 30648
rect 17451 30617 17463 30620
rect 17405 30611 17463 30617
rect 17770 30608 17776 30620
rect 17828 30608 17834 30660
rect 18141 30651 18199 30657
rect 18141 30617 18153 30651
rect 18187 30648 18199 30651
rect 18782 30648 18788 30660
rect 18187 30620 18788 30648
rect 18187 30617 18199 30620
rect 18141 30611 18199 30617
rect 18782 30608 18788 30620
rect 18840 30648 18846 30660
rect 19061 30651 19119 30657
rect 19061 30648 19073 30651
rect 18840 30620 19073 30648
rect 18840 30608 18846 30620
rect 19061 30617 19073 30620
rect 19107 30617 19119 30651
rect 19061 30611 19119 30617
rect 14332 30552 14964 30580
rect 14332 30540 14338 30552
rect 15194 30540 15200 30592
rect 15252 30580 15258 30592
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 15252 30552 15485 30580
rect 15252 30540 15258 30552
rect 15473 30549 15485 30552
rect 15519 30549 15531 30583
rect 15473 30543 15531 30549
rect 17034 30540 17040 30592
rect 17092 30540 17098 30592
rect 18598 30540 18604 30592
rect 18656 30580 18662 30592
rect 19996 30580 20024 30688
rect 20346 30676 20352 30728
rect 20404 30676 20410 30728
rect 20625 30719 20683 30725
rect 20625 30685 20637 30719
rect 20671 30716 20683 30719
rect 20714 30716 20720 30728
rect 20671 30688 20720 30716
rect 20671 30685 20683 30688
rect 20625 30679 20683 30685
rect 20714 30676 20720 30688
rect 20772 30676 20778 30728
rect 22097 30719 22155 30725
rect 22097 30685 22109 30719
rect 22143 30716 22155 30719
rect 22922 30716 22928 30728
rect 22143 30688 22928 30716
rect 22143 30685 22155 30688
rect 22097 30679 22155 30685
rect 22922 30676 22928 30688
rect 22980 30676 22986 30728
rect 24044 30716 24072 30744
rect 25222 30716 25228 30728
rect 24044 30688 25228 30716
rect 25222 30676 25228 30688
rect 25280 30716 25286 30728
rect 25280 30688 25544 30716
rect 25280 30676 25286 30688
rect 25516 30657 25544 30688
rect 25501 30651 25559 30657
rect 25501 30617 25513 30651
rect 25547 30617 25559 30651
rect 25608 30648 25636 30824
rect 25700 30716 25728 30880
rect 26234 30812 26240 30864
rect 26292 30852 26298 30864
rect 26292 30824 26335 30852
rect 26292 30812 26298 30824
rect 25866 30744 25872 30796
rect 25924 30784 25930 30796
rect 26053 30787 26111 30793
rect 26053 30784 26065 30787
rect 25924 30756 26065 30784
rect 25924 30744 25930 30756
rect 26053 30753 26065 30756
rect 26099 30753 26111 30787
rect 26528 30784 26556 30892
rect 27614 30880 27620 30892
rect 27672 30880 27678 30932
rect 28166 30880 28172 30932
rect 28224 30920 28230 30932
rect 28261 30923 28319 30929
rect 28261 30920 28273 30923
rect 28224 30892 28273 30920
rect 28224 30880 28230 30892
rect 28261 30889 28273 30892
rect 28307 30920 28319 30923
rect 28718 30920 28724 30932
rect 28307 30892 28724 30920
rect 28307 30889 28319 30892
rect 28261 30883 28319 30889
rect 28718 30880 28724 30892
rect 28776 30880 28782 30932
rect 32582 30920 32588 30932
rect 30208 30892 32588 30920
rect 30208 30861 30236 30892
rect 32582 30880 32588 30892
rect 32640 30880 32646 30932
rect 30193 30855 30251 30861
rect 28014 30824 30144 30852
rect 26053 30747 26111 30753
rect 26160 30756 26556 30784
rect 26160 30716 26188 30756
rect 28258 30744 28264 30796
rect 28316 30784 28322 30796
rect 28810 30784 28816 30796
rect 28316 30756 28816 30784
rect 28316 30744 28322 30756
rect 28810 30744 28816 30756
rect 28868 30744 28874 30796
rect 28997 30787 29055 30793
rect 28997 30753 29009 30787
rect 29043 30784 29055 30787
rect 29822 30784 29828 30796
rect 29043 30756 29828 30784
rect 29043 30753 29055 30756
rect 28997 30747 29055 30753
rect 29822 30744 29828 30756
rect 29880 30744 29886 30796
rect 30116 30784 30144 30824
rect 30193 30821 30205 30855
rect 30239 30821 30251 30855
rect 30193 30815 30251 30821
rect 31570 30812 31576 30864
rect 31628 30812 31634 30864
rect 30374 30784 30380 30796
rect 30116 30756 30380 30784
rect 30374 30744 30380 30756
rect 30432 30744 30438 30796
rect 30469 30787 30527 30793
rect 30469 30753 30481 30787
rect 30515 30753 30527 30787
rect 30469 30747 30527 30753
rect 25700 30688 26188 30716
rect 26513 30719 26571 30725
rect 26513 30685 26525 30719
rect 26559 30685 26571 30719
rect 26513 30679 26571 30685
rect 26418 30648 26424 30660
rect 25608 30620 26424 30648
rect 25501 30611 25559 30617
rect 26418 30608 26424 30620
rect 26476 30608 26482 30660
rect 18656 30552 20024 30580
rect 18656 30540 18662 30552
rect 20254 30540 20260 30592
rect 20312 30540 20318 30592
rect 22278 30540 22284 30592
rect 22336 30540 22342 30592
rect 24578 30540 24584 30592
rect 24636 30540 24642 30592
rect 26234 30540 26240 30592
rect 26292 30580 26298 30592
rect 26528 30580 26556 30679
rect 26786 30676 26792 30728
rect 26844 30676 26850 30728
rect 29730 30676 29736 30728
rect 29788 30716 29794 30728
rect 30484 30716 30512 30747
rect 29788 30688 30512 30716
rect 29788 30676 29794 30688
rect 26292 30552 26556 30580
rect 26292 30540 26298 30552
rect 28718 30540 28724 30592
rect 28776 30540 28782 30592
rect 2760 30490 32200 30512
rect 2760 30438 6286 30490
rect 6338 30438 6350 30490
rect 6402 30438 6414 30490
rect 6466 30438 6478 30490
rect 6530 30438 6542 30490
rect 6594 30438 13646 30490
rect 13698 30438 13710 30490
rect 13762 30438 13774 30490
rect 13826 30438 13838 30490
rect 13890 30438 13902 30490
rect 13954 30438 21006 30490
rect 21058 30438 21070 30490
rect 21122 30438 21134 30490
rect 21186 30438 21198 30490
rect 21250 30438 21262 30490
rect 21314 30438 28366 30490
rect 28418 30438 28430 30490
rect 28482 30438 28494 30490
rect 28546 30438 28558 30490
rect 28610 30438 28622 30490
rect 28674 30438 32200 30490
rect 2760 30416 32200 30438
rect 14645 30379 14703 30385
rect 14645 30345 14657 30379
rect 14691 30345 14703 30379
rect 16574 30376 16580 30388
rect 14645 30339 14703 30345
rect 12342 30268 12348 30320
rect 12400 30268 12406 30320
rect 2774 30200 2780 30252
rect 2832 30240 2838 30252
rect 3237 30243 3295 30249
rect 3237 30240 3249 30243
rect 2832 30212 3249 30240
rect 2832 30200 2838 30212
rect 3237 30209 3249 30212
rect 3283 30209 3295 30243
rect 3237 30203 3295 30209
rect 9674 30200 9680 30252
rect 9732 30200 9738 30252
rect 10597 30243 10655 30249
rect 10597 30209 10609 30243
rect 10643 30240 10655 30243
rect 10870 30240 10876 30252
rect 10643 30212 10876 30240
rect 10643 30209 10655 30212
rect 10597 30203 10655 30209
rect 10870 30200 10876 30212
rect 10928 30200 10934 30252
rect 12805 30243 12863 30249
rect 12805 30209 12817 30243
rect 12851 30240 12863 30243
rect 14182 30240 14188 30252
rect 12851 30212 14188 30240
rect 12851 30209 12863 30212
rect 12805 30203 12863 30209
rect 14182 30200 14188 30212
rect 14240 30200 14246 30252
rect 14274 30200 14280 30252
rect 14332 30240 14338 30252
rect 14553 30243 14611 30249
rect 14553 30240 14565 30243
rect 14332 30212 14565 30240
rect 14332 30200 14338 30212
rect 14553 30209 14565 30212
rect 14599 30209 14611 30243
rect 14553 30203 14611 30209
rect 4433 30175 4491 30181
rect 4433 30141 4445 30175
rect 4479 30172 4491 30175
rect 4522 30172 4528 30184
rect 4479 30144 4528 30172
rect 4479 30141 4491 30144
rect 4433 30135 4491 30141
rect 4522 30132 4528 30144
rect 4580 30132 4586 30184
rect 8205 30175 8263 30181
rect 8205 30172 8217 30175
rect 7668 30144 8217 30172
rect 7668 30048 7696 30144
rect 8205 30141 8217 30144
rect 8251 30141 8263 30175
rect 8205 30135 8263 30141
rect 11974 30132 11980 30184
rect 12032 30132 12038 30184
rect 10318 30064 10324 30116
rect 10376 30104 10382 30116
rect 10873 30107 10931 30113
rect 10873 30104 10885 30107
rect 10376 30076 10885 30104
rect 10376 30064 10382 30076
rect 10873 30073 10885 30076
rect 10919 30073 10931 30107
rect 10873 30067 10931 30073
rect 12894 30064 12900 30116
rect 12952 30104 12958 30116
rect 14277 30107 14335 30113
rect 12952 30076 13110 30104
rect 12952 30064 12958 30076
rect 14277 30073 14289 30107
rect 14323 30104 14335 30107
rect 14660 30104 14688 30339
rect 16546 30336 16580 30376
rect 16632 30336 16638 30388
rect 16942 30336 16948 30388
rect 17000 30336 17006 30388
rect 17310 30336 17316 30388
rect 17368 30336 17374 30388
rect 20714 30336 20720 30388
rect 20772 30376 20778 30388
rect 22094 30376 22100 30388
rect 20772 30348 20944 30376
rect 20772 30336 20778 30348
rect 16025 30311 16083 30317
rect 16025 30277 16037 30311
rect 16071 30308 16083 30311
rect 16546 30308 16574 30336
rect 16071 30280 16574 30308
rect 16071 30277 16083 30280
rect 16025 30271 16083 30277
rect 14734 30200 14740 30252
rect 14792 30240 14798 30252
rect 15194 30240 15200 30252
rect 14792 30212 15200 30240
rect 14792 30200 14798 30212
rect 15194 30200 15200 30212
rect 15252 30240 15258 30252
rect 16577 30243 16635 30249
rect 16577 30240 16589 30243
rect 15252 30212 16589 30240
rect 15252 30200 15258 30212
rect 16577 30209 16589 30212
rect 16623 30209 16635 30243
rect 17328 30240 17356 30336
rect 18966 30268 18972 30320
rect 19024 30268 19030 30320
rect 20916 30317 20944 30348
rect 21008 30348 22100 30376
rect 20901 30311 20959 30317
rect 20901 30277 20913 30311
rect 20947 30277 20959 30311
rect 20901 30271 20959 30277
rect 16577 30203 16635 30209
rect 16776 30212 17356 30240
rect 15013 30175 15071 30181
rect 15013 30141 15025 30175
rect 15059 30172 15071 30175
rect 15102 30172 15108 30184
rect 15059 30144 15108 30172
rect 15059 30141 15071 30144
rect 15013 30135 15071 30141
rect 15102 30132 15108 30144
rect 15160 30132 15166 30184
rect 16393 30175 16451 30181
rect 16393 30141 16405 30175
rect 16439 30172 16451 30175
rect 16776 30172 16804 30212
rect 17494 30200 17500 30252
rect 17552 30200 17558 30252
rect 19334 30240 19340 30252
rect 19260 30212 19340 30240
rect 16439 30144 16804 30172
rect 16853 30175 16911 30181
rect 16439 30141 16451 30144
rect 16393 30135 16451 30141
rect 16853 30141 16865 30175
rect 16899 30141 16911 30175
rect 16853 30135 16911 30141
rect 14323 30076 14688 30104
rect 14323 30073 14335 30076
rect 14277 30067 14335 30073
rect 16298 30064 16304 30116
rect 16356 30104 16362 30116
rect 16485 30107 16543 30113
rect 16485 30104 16497 30107
rect 16356 30076 16497 30104
rect 16356 30064 16362 30076
rect 16485 30073 16497 30076
rect 16531 30073 16543 30107
rect 16485 30067 16543 30073
rect 7650 29996 7656 30048
rect 7708 29996 7714 30048
rect 8294 29996 8300 30048
rect 8352 29996 8358 30048
rect 8754 29996 8760 30048
rect 8812 30036 8818 30048
rect 9125 30039 9183 30045
rect 9125 30036 9137 30039
rect 8812 30008 9137 30036
rect 8812 29996 8818 30008
rect 9125 30005 9137 30008
rect 9171 30005 9183 30039
rect 9125 29999 9183 30005
rect 11882 29996 11888 30048
rect 11940 30036 11946 30048
rect 15105 30039 15163 30045
rect 15105 30036 15117 30039
rect 11940 30008 15117 30036
rect 11940 29996 11946 30008
rect 15105 30005 15117 30008
rect 15151 30005 15163 30039
rect 15105 29999 15163 30005
rect 15930 29996 15936 30048
rect 15988 30036 15994 30048
rect 16868 30036 16896 30135
rect 17034 30132 17040 30184
rect 17092 30172 17098 30184
rect 19260 30181 19288 30212
rect 19334 30200 19340 30212
rect 19392 30240 19398 30252
rect 21008 30240 21036 30348
rect 22094 30336 22100 30348
rect 22152 30376 22158 30388
rect 22554 30376 22560 30388
rect 22152 30348 22560 30376
rect 22152 30336 22158 30348
rect 22554 30336 22560 30348
rect 22612 30336 22618 30388
rect 23477 30379 23535 30385
rect 23477 30345 23489 30379
rect 23523 30376 23535 30379
rect 23842 30376 23848 30388
rect 23523 30348 23848 30376
rect 23523 30345 23535 30348
rect 23477 30339 23535 30345
rect 23842 30336 23848 30348
rect 23900 30336 23906 30388
rect 23934 30336 23940 30388
rect 23992 30376 23998 30388
rect 24394 30376 24400 30388
rect 23992 30348 24400 30376
rect 23992 30336 23998 30348
rect 24394 30336 24400 30348
rect 24452 30336 24458 30388
rect 24946 30336 24952 30388
rect 25004 30336 25010 30388
rect 25314 30336 25320 30388
rect 25372 30336 25378 30388
rect 26878 30376 26884 30388
rect 26252 30348 26884 30376
rect 24964 30308 24992 30336
rect 25409 30311 25467 30317
rect 25409 30308 25421 30311
rect 24964 30280 25421 30308
rect 25409 30277 25421 30280
rect 25455 30277 25467 30311
rect 25409 30271 25467 30277
rect 26053 30311 26111 30317
rect 26053 30277 26065 30311
rect 26099 30308 26111 30311
rect 26252 30308 26280 30348
rect 26878 30336 26884 30348
rect 26936 30336 26942 30388
rect 27522 30336 27528 30388
rect 27580 30376 27586 30388
rect 27580 30348 27752 30376
rect 27580 30336 27586 30348
rect 26099 30280 26280 30308
rect 27724 30308 27752 30348
rect 28810 30336 28816 30388
rect 28868 30376 28874 30388
rect 28868 30348 30144 30376
rect 28868 30336 28874 30348
rect 28537 30311 28595 30317
rect 28537 30308 28549 30311
rect 27724 30280 28549 30308
rect 26099 30277 26111 30280
rect 26053 30271 26111 30277
rect 28537 30277 28549 30280
rect 28583 30308 28595 30311
rect 28721 30311 28779 30317
rect 28721 30308 28733 30311
rect 28583 30280 28733 30308
rect 28583 30277 28595 30280
rect 28537 30271 28595 30277
rect 28721 30277 28733 30280
rect 28767 30277 28779 30311
rect 28721 30271 28779 30277
rect 19392 30212 21036 30240
rect 21453 30243 21511 30249
rect 19392 30200 19398 30212
rect 17221 30175 17279 30181
rect 17221 30172 17233 30175
rect 17092 30144 17233 30172
rect 17092 30132 17098 30144
rect 17221 30141 17233 30144
rect 17267 30141 17279 30175
rect 17221 30135 17279 30141
rect 19245 30175 19303 30181
rect 19245 30141 19257 30175
rect 19291 30141 19303 30175
rect 19245 30135 19303 30141
rect 20254 30132 20260 30184
rect 20312 30132 20318 30184
rect 20456 30181 20484 30212
rect 21453 30209 21465 30243
rect 21499 30209 21511 30243
rect 21453 30203 21511 30209
rect 21729 30243 21787 30249
rect 21729 30209 21741 30243
rect 21775 30240 21787 30243
rect 22094 30240 22100 30252
rect 21775 30212 22100 30240
rect 21775 30209 21787 30212
rect 21729 30203 21787 30209
rect 20441 30175 20499 30181
rect 20441 30141 20453 30175
rect 20487 30141 20499 30175
rect 21468 30172 21496 30203
rect 22094 30200 22100 30212
rect 22152 30240 22158 30252
rect 23474 30240 23480 30252
rect 22152 30212 23480 30240
rect 22152 30200 22158 30212
rect 23474 30200 23480 30212
rect 23532 30240 23538 30252
rect 23569 30243 23627 30249
rect 23569 30240 23581 30243
rect 23532 30212 23581 30240
rect 23532 30200 23538 30212
rect 23569 30209 23581 30212
rect 23615 30209 23627 30243
rect 23569 30203 23627 30209
rect 23845 30243 23903 30249
rect 23845 30209 23857 30243
rect 23891 30240 23903 30243
rect 24578 30240 24584 30252
rect 23891 30212 24584 30240
rect 23891 30209 23903 30212
rect 23845 30203 23903 30209
rect 24578 30200 24584 30212
rect 24636 30200 24642 30252
rect 25222 30200 25228 30252
rect 25280 30240 25286 30252
rect 26068 30240 26096 30271
rect 27062 30240 27068 30252
rect 25280 30212 25636 30240
rect 25280 30200 25286 30212
rect 21542 30172 21548 30184
rect 21468 30144 21548 30172
rect 20441 30135 20499 30141
rect 21542 30132 21548 30144
rect 21600 30132 21606 30184
rect 25498 30172 25504 30184
rect 24978 30144 25504 30172
rect 25498 30132 25504 30144
rect 25556 30132 25562 30184
rect 25608 30181 25636 30212
rect 25792 30212 26096 30240
rect 26160 30212 27068 30240
rect 25792 30181 25820 30212
rect 25593 30175 25651 30181
rect 25593 30141 25605 30175
rect 25639 30141 25651 30175
rect 25593 30135 25651 30141
rect 25777 30175 25835 30181
rect 25777 30141 25789 30175
rect 25823 30141 25835 30175
rect 25777 30135 25835 30141
rect 25866 30132 25872 30184
rect 25924 30172 25930 30184
rect 26160 30172 26188 30212
rect 27062 30200 27068 30212
rect 27120 30200 27126 30252
rect 27154 30200 27160 30252
rect 27212 30240 27218 30252
rect 27525 30243 27583 30249
rect 27525 30240 27537 30243
rect 27212 30212 27537 30240
rect 27212 30200 27218 30212
rect 27525 30209 27537 30212
rect 27571 30209 27583 30243
rect 27525 30203 27583 30209
rect 27801 30243 27859 30249
rect 27801 30209 27813 30243
rect 27847 30240 27859 30243
rect 30116 30240 30144 30348
rect 30374 30336 30380 30388
rect 30432 30336 30438 30388
rect 30392 30308 30420 30336
rect 30929 30311 30987 30317
rect 30929 30308 30941 30311
rect 30392 30280 30941 30308
rect 30929 30277 30941 30280
rect 30975 30277 30987 30311
rect 30929 30271 30987 30277
rect 33042 30240 33048 30252
rect 27847 30212 28948 30240
rect 27847 30209 27859 30212
rect 27801 30203 27859 30209
rect 28920 30184 28948 30212
rect 29196 30212 30052 30240
rect 30116 30212 31064 30240
rect 25924 30144 26188 30172
rect 25924 30132 25930 30144
rect 27890 30132 27896 30184
rect 27948 30132 27954 30184
rect 28258 30132 28264 30184
rect 28316 30172 28322 30184
rect 28629 30175 28687 30181
rect 28629 30172 28641 30175
rect 28316 30144 28641 30172
rect 28316 30132 28322 30144
rect 28629 30141 28641 30144
rect 28675 30141 28687 30175
rect 28629 30135 28687 30141
rect 28902 30132 28908 30184
rect 28960 30132 28966 30184
rect 29196 30181 29224 30212
rect 30024 30184 30052 30212
rect 29148 30175 29224 30181
rect 29148 30141 29160 30175
rect 29194 30144 29224 30175
rect 29194 30141 29206 30144
rect 29148 30135 29206 30141
rect 29914 30132 29920 30184
rect 29972 30132 29978 30184
rect 30006 30132 30012 30184
rect 30064 30132 30070 30184
rect 30650 30132 30656 30184
rect 30708 30132 30714 30184
rect 30926 30132 30932 30184
rect 30984 30172 30990 30184
rect 31036 30181 31064 30212
rect 31864 30212 33048 30240
rect 31864 30181 31892 30212
rect 33042 30200 33048 30212
rect 33100 30200 33106 30252
rect 31021 30175 31079 30181
rect 31021 30172 31033 30175
rect 30984 30144 31033 30172
rect 30984 30132 30990 30144
rect 31021 30141 31033 30144
rect 31067 30172 31079 30175
rect 31389 30175 31447 30181
rect 31389 30172 31401 30175
rect 31067 30144 31401 30172
rect 31067 30141 31079 30144
rect 31021 30135 31079 30141
rect 31389 30141 31401 30144
rect 31435 30141 31447 30175
rect 31389 30135 31447 30141
rect 31849 30175 31907 30181
rect 31849 30141 31861 30175
rect 31895 30141 31907 30175
rect 31849 30135 31907 30141
rect 19153 30107 19211 30113
rect 19153 30104 19165 30107
rect 18722 30076 19165 30104
rect 19153 30073 19165 30076
rect 19199 30073 19211 30107
rect 19153 30067 19211 30073
rect 19613 30107 19671 30113
rect 19613 30073 19625 30107
rect 19659 30104 19671 30107
rect 21269 30107 21327 30113
rect 19659 30076 20944 30104
rect 19659 30073 19671 30076
rect 19613 30067 19671 30073
rect 19904 30048 19932 30076
rect 15988 30008 16896 30036
rect 15988 29996 15994 30008
rect 19702 29996 19708 30048
rect 19760 29996 19766 30048
rect 19886 29996 19892 30048
rect 19944 29996 19950 30048
rect 20438 29996 20444 30048
rect 20496 30036 20502 30048
rect 20533 30039 20591 30045
rect 20533 30036 20545 30039
rect 20496 30008 20545 30036
rect 20496 29996 20502 30008
rect 20533 30005 20545 30008
rect 20579 30005 20591 30039
rect 20916 30036 20944 30076
rect 21269 30073 21281 30107
rect 21315 30104 21327 30107
rect 21315 30076 21772 30104
rect 21315 30073 21327 30076
rect 21269 30067 21327 30073
rect 21361 30039 21419 30045
rect 21361 30036 21373 30039
rect 20916 30008 21373 30036
rect 20533 29999 20591 30005
rect 21361 30005 21373 30008
rect 21407 30005 21419 30039
rect 21744 30036 21772 30076
rect 22002 30064 22008 30116
rect 22060 30064 22066 30116
rect 22738 30064 22744 30116
rect 22796 30064 22802 30116
rect 25958 30064 25964 30116
rect 26016 30104 26022 30116
rect 26016 30076 26358 30104
rect 26016 30064 26022 30076
rect 28350 30064 28356 30116
rect 28408 30104 28414 30116
rect 28408 30076 29316 30104
rect 28408 30064 28414 30076
rect 22278 30036 22284 30048
rect 21744 30008 22284 30036
rect 21361 29999 21419 30005
rect 22278 29996 22284 30008
rect 22336 29996 22342 30048
rect 22922 29996 22928 30048
rect 22980 30036 22986 30048
rect 27154 30036 27160 30048
rect 22980 30008 27160 30036
rect 22980 29996 22986 30008
rect 27154 29996 27160 30008
rect 27212 29996 27218 30048
rect 27246 29996 27252 30048
rect 27304 30036 27310 30048
rect 29288 30045 29316 30076
rect 29089 30039 29147 30045
rect 29089 30036 29101 30039
rect 27304 30008 29101 30036
rect 27304 29996 27310 30008
rect 29089 30005 29101 30008
rect 29135 30005 29147 30039
rect 29089 29999 29147 30005
rect 29273 30039 29331 30045
rect 29273 30005 29285 30039
rect 29319 30005 29331 30039
rect 29273 29999 29331 30005
rect 29362 29996 29368 30048
rect 29420 29996 29426 30048
rect 29546 29996 29552 30048
rect 29604 30036 29610 30048
rect 30101 30039 30159 30045
rect 30101 30036 30113 30039
rect 29604 30008 30113 30036
rect 29604 29996 29610 30008
rect 30101 30005 30113 30008
rect 30147 30005 30159 30039
rect 30101 29999 30159 30005
rect 31294 29996 31300 30048
rect 31352 29996 31358 30048
rect 31478 29996 31484 30048
rect 31536 30036 31542 30048
rect 31665 30039 31723 30045
rect 31665 30036 31677 30039
rect 31536 30008 31677 30036
rect 31536 29996 31542 30008
rect 31665 30005 31677 30008
rect 31711 30005 31723 30039
rect 31665 29999 31723 30005
rect 2760 29946 32200 29968
rect 2760 29894 6946 29946
rect 6998 29894 7010 29946
rect 7062 29894 7074 29946
rect 7126 29894 7138 29946
rect 7190 29894 7202 29946
rect 7254 29894 14306 29946
rect 14358 29894 14370 29946
rect 14422 29894 14434 29946
rect 14486 29894 14498 29946
rect 14550 29894 14562 29946
rect 14614 29894 21666 29946
rect 21718 29894 21730 29946
rect 21782 29894 21794 29946
rect 21846 29894 21858 29946
rect 21910 29894 21922 29946
rect 21974 29894 29026 29946
rect 29078 29894 29090 29946
rect 29142 29894 29154 29946
rect 29206 29894 29218 29946
rect 29270 29894 29282 29946
rect 29334 29894 32200 29946
rect 2760 29872 32200 29894
rect 4430 29792 4436 29844
rect 4488 29832 4494 29844
rect 4525 29835 4583 29841
rect 4525 29832 4537 29835
rect 4488 29804 4537 29832
rect 4488 29792 4494 29804
rect 4525 29801 4537 29804
rect 4571 29801 4583 29835
rect 4525 29795 4583 29801
rect 9674 29792 9680 29844
rect 9732 29832 9738 29844
rect 9769 29835 9827 29841
rect 9769 29832 9781 29835
rect 9732 29804 9781 29832
rect 9732 29792 9738 29804
rect 9769 29801 9781 29804
rect 9815 29801 9827 29835
rect 9769 29795 9827 29801
rect 10318 29792 10324 29844
rect 10376 29792 10382 29844
rect 11974 29792 11980 29844
rect 12032 29792 12038 29844
rect 12342 29792 12348 29844
rect 12400 29792 12406 29844
rect 12989 29835 13047 29841
rect 12989 29801 13001 29835
rect 13035 29832 13047 29835
rect 13538 29832 13544 29844
rect 13035 29804 13544 29832
rect 13035 29801 13047 29804
rect 12989 29795 13047 29801
rect 13538 29792 13544 29804
rect 13596 29792 13602 29844
rect 13909 29835 13967 29841
rect 13909 29801 13921 29835
rect 13955 29832 13967 29835
rect 15010 29832 15016 29844
rect 13955 29804 15016 29832
rect 13955 29801 13967 29804
rect 13909 29795 13967 29801
rect 15010 29792 15016 29804
rect 15068 29792 15074 29844
rect 15194 29792 15200 29844
rect 15252 29832 15258 29844
rect 15565 29835 15623 29841
rect 15565 29832 15577 29835
rect 15252 29804 15577 29832
rect 15252 29792 15258 29804
rect 15565 29801 15577 29804
rect 15611 29801 15623 29835
rect 15565 29795 15623 29801
rect 17221 29835 17279 29841
rect 17221 29801 17233 29835
rect 17267 29832 17279 29835
rect 18046 29832 18052 29844
rect 17267 29804 18052 29832
rect 17267 29801 17279 29804
rect 17221 29795 17279 29801
rect 8294 29724 8300 29776
rect 8352 29764 8358 29776
rect 11425 29767 11483 29773
rect 8352 29736 8786 29764
rect 8352 29724 8358 29736
rect 11425 29733 11437 29767
rect 11471 29764 11483 29767
rect 12360 29764 12388 29792
rect 15102 29764 15108 29776
rect 11471 29736 12388 29764
rect 14108 29736 15108 29764
rect 11471 29733 11483 29736
rect 11425 29727 11483 29733
rect 3142 29656 3148 29708
rect 3200 29656 3206 29708
rect 4709 29699 4767 29705
rect 4709 29665 4721 29699
rect 4755 29696 4767 29699
rect 12069 29699 12127 29705
rect 4755 29668 5120 29696
rect 4755 29665 4767 29668
rect 4709 29659 4767 29665
rect 3510 29588 3516 29640
rect 3568 29588 3574 29640
rect 5092 29501 5120 29668
rect 12069 29665 12081 29699
rect 12115 29665 12127 29699
rect 14108 29696 14136 29736
rect 15102 29724 15108 29736
rect 15160 29724 15166 29776
rect 15580 29764 15608 29795
rect 18046 29792 18052 29804
rect 18104 29792 18110 29844
rect 18966 29792 18972 29844
rect 19024 29792 19030 29844
rect 20346 29832 20352 29844
rect 19444 29804 20352 29832
rect 16853 29767 16911 29773
rect 15580 29736 16528 29764
rect 12069 29659 12127 29665
rect 12176 29668 14136 29696
rect 14645 29699 14703 29705
rect 7374 29588 7380 29640
rect 7432 29628 7438 29640
rect 8021 29631 8079 29637
rect 8021 29628 8033 29631
rect 7432 29600 8033 29628
rect 7432 29588 7438 29600
rect 8021 29597 8033 29600
rect 8067 29597 8079 29631
rect 8021 29591 8079 29597
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 10965 29631 11023 29637
rect 10965 29597 10977 29631
rect 11011 29628 11023 29631
rect 11011 29600 11100 29628
rect 11011 29597 11023 29600
rect 10965 29591 11023 29597
rect 11072 29569 11100 29600
rect 11238 29588 11244 29640
rect 11296 29628 11302 29640
rect 11517 29631 11575 29637
rect 11517 29628 11529 29631
rect 11296 29600 11529 29628
rect 11296 29588 11302 29600
rect 11517 29597 11529 29600
rect 11563 29597 11575 29631
rect 11517 29591 11575 29597
rect 11606 29588 11612 29640
rect 11664 29588 11670 29640
rect 12084 29572 12112 29659
rect 11057 29563 11115 29569
rect 11057 29529 11069 29563
rect 11103 29529 11115 29563
rect 11057 29523 11115 29529
rect 12066 29520 12072 29572
rect 12124 29520 12130 29572
rect 5077 29495 5135 29501
rect 5077 29461 5089 29495
rect 5123 29492 5135 29495
rect 12176 29492 12204 29668
rect 14645 29665 14657 29699
rect 14691 29696 14703 29699
rect 14826 29696 14832 29708
rect 14691 29668 14832 29696
rect 14691 29665 14703 29668
rect 14645 29659 14703 29665
rect 14826 29656 14832 29668
rect 14884 29656 14890 29708
rect 14921 29699 14979 29705
rect 14921 29665 14933 29699
rect 14967 29696 14979 29699
rect 16298 29696 16304 29708
rect 14967 29668 16304 29696
rect 14967 29665 14979 29668
rect 14921 29659 14979 29665
rect 16298 29656 16304 29668
rect 16356 29696 16362 29708
rect 16393 29699 16451 29705
rect 16393 29696 16405 29699
rect 16356 29668 16405 29696
rect 16356 29656 16362 29668
rect 16393 29665 16405 29668
rect 16439 29665 16451 29699
rect 16393 29659 16451 29665
rect 12437 29631 12495 29637
rect 12437 29597 12449 29631
rect 12483 29628 12495 29631
rect 12483 29600 13584 29628
rect 12483 29597 12495 29600
rect 12437 29591 12495 29597
rect 13556 29569 13584 29600
rect 13630 29588 13636 29640
rect 13688 29628 13694 29640
rect 14001 29631 14059 29637
rect 14001 29628 14013 29631
rect 13688 29600 14013 29628
rect 13688 29588 13694 29600
rect 14001 29597 14013 29600
rect 14047 29597 14059 29631
rect 14001 29591 14059 29597
rect 14090 29588 14096 29640
rect 14148 29588 14154 29640
rect 14553 29631 14611 29637
rect 14553 29597 14565 29631
rect 14599 29628 14611 29631
rect 14734 29628 14740 29640
rect 14599 29600 14740 29628
rect 14599 29597 14611 29600
rect 14553 29591 14611 29597
rect 14734 29588 14740 29600
rect 14792 29588 14798 29640
rect 15013 29631 15071 29637
rect 15013 29597 15025 29631
rect 15059 29597 15071 29631
rect 15013 29591 15071 29597
rect 13541 29563 13599 29569
rect 13541 29529 13553 29563
rect 13587 29529 13599 29563
rect 15028 29560 15056 29591
rect 15746 29588 15752 29640
rect 15804 29588 15810 29640
rect 13541 29523 13599 29529
rect 13648 29532 15056 29560
rect 16500 29560 16528 29736
rect 16853 29733 16865 29767
rect 16899 29764 16911 29767
rect 18984 29764 19012 29792
rect 16899 29736 19012 29764
rect 16899 29733 16911 29736
rect 16853 29727 16911 29733
rect 19334 29724 19340 29776
rect 19392 29724 19398 29776
rect 17681 29699 17739 29705
rect 16684 29668 17448 29696
rect 16574 29588 16580 29640
rect 16632 29588 16638 29640
rect 16684 29560 16712 29668
rect 17420 29637 17448 29668
rect 17681 29665 17693 29699
rect 17727 29696 17739 29699
rect 18506 29696 18512 29708
rect 17727 29668 18512 29696
rect 17727 29665 17739 29668
rect 17681 29659 17739 29665
rect 18506 29656 18512 29668
rect 18564 29656 18570 29708
rect 19245 29699 19303 29705
rect 19245 29665 19257 29699
rect 19291 29696 19303 29699
rect 19352 29696 19380 29724
rect 19444 29705 19472 29804
rect 20346 29792 20352 29804
rect 20404 29792 20410 29844
rect 20714 29792 20720 29844
rect 20772 29832 20778 29844
rect 21177 29835 21235 29841
rect 21177 29832 21189 29835
rect 20772 29804 21189 29832
rect 20772 29792 20778 29804
rect 21177 29801 21189 29804
rect 21223 29832 21235 29835
rect 21450 29832 21456 29844
rect 21223 29804 21456 29832
rect 21223 29801 21235 29804
rect 21177 29795 21235 29801
rect 21450 29792 21456 29804
rect 21508 29792 21514 29844
rect 22002 29792 22008 29844
rect 22060 29792 22066 29844
rect 22738 29792 22744 29844
rect 22796 29792 22802 29844
rect 23750 29792 23756 29844
rect 23808 29792 23814 29844
rect 24486 29792 24492 29844
rect 24544 29832 24550 29844
rect 24762 29832 24768 29844
rect 24544 29804 24768 29832
rect 24544 29792 24550 29804
rect 24762 29792 24768 29804
rect 24820 29832 24826 29844
rect 25133 29835 25191 29841
rect 25133 29832 25145 29835
rect 24820 29804 25145 29832
rect 24820 29792 24826 29804
rect 25133 29801 25145 29804
rect 25179 29801 25191 29835
rect 25133 29795 25191 29801
rect 25682 29792 25688 29844
rect 25740 29792 25746 29844
rect 25777 29835 25835 29841
rect 25777 29801 25789 29835
rect 25823 29832 25835 29835
rect 26326 29832 26332 29844
rect 25823 29804 26332 29832
rect 25823 29801 25835 29804
rect 25777 29795 25835 29801
rect 26326 29792 26332 29804
rect 26384 29792 26390 29844
rect 27617 29835 27675 29841
rect 27617 29801 27629 29835
rect 27663 29832 27675 29835
rect 27890 29832 27896 29844
rect 27663 29804 27896 29832
rect 27663 29801 27675 29804
rect 27617 29795 27675 29801
rect 27890 29792 27896 29804
rect 27948 29792 27954 29844
rect 28813 29835 28871 29841
rect 28813 29801 28825 29835
rect 28859 29801 28871 29835
rect 28813 29795 28871 29801
rect 19702 29724 19708 29776
rect 19760 29724 19766 29776
rect 20438 29724 20444 29776
rect 20496 29724 20502 29776
rect 22020 29764 22048 29792
rect 23477 29767 23535 29773
rect 23477 29764 23489 29767
rect 22020 29736 23489 29764
rect 23477 29733 23489 29736
rect 23523 29733 23535 29767
rect 23477 29727 23535 29733
rect 19291 29668 19380 29696
rect 19429 29699 19487 29705
rect 19291 29665 19303 29668
rect 19245 29659 19303 29665
rect 19429 29665 19441 29699
rect 19475 29665 19487 29699
rect 19429 29659 19487 29665
rect 22554 29656 22560 29708
rect 22612 29696 22618 29708
rect 22649 29699 22707 29705
rect 22649 29696 22661 29699
rect 22612 29668 22661 29696
rect 22612 29656 22618 29668
rect 22649 29665 22661 29668
rect 22695 29665 22707 29699
rect 22649 29659 22707 29665
rect 23017 29699 23075 29705
rect 23017 29665 23029 29699
rect 23063 29696 23075 29699
rect 23106 29696 23112 29708
rect 23063 29668 23112 29696
rect 23063 29665 23075 29668
rect 23017 29659 23075 29665
rect 23106 29656 23112 29668
rect 23164 29656 23170 29708
rect 23201 29699 23259 29705
rect 23201 29665 23213 29699
rect 23247 29665 23259 29699
rect 23201 29659 23259 29665
rect 23293 29699 23351 29705
rect 23293 29665 23305 29699
rect 23339 29696 23351 29699
rect 23768 29696 23796 29792
rect 23339 29668 23796 29696
rect 23860 29736 25268 29764
rect 23339 29665 23351 29668
rect 23293 29659 23351 29665
rect 16761 29631 16819 29637
rect 16761 29597 16773 29631
rect 16807 29628 16819 29631
rect 17405 29631 17463 29637
rect 16807 29600 16896 29628
rect 16807 29597 16819 29600
rect 16761 29591 16819 29597
rect 16500 29532 16712 29560
rect 5123 29464 12204 29492
rect 5123 29461 5135 29464
rect 5077 29455 5135 29461
rect 13446 29452 13452 29504
rect 13504 29492 13510 29504
rect 13648 29492 13676 29532
rect 16868 29504 16896 29600
rect 17405 29597 17417 29631
rect 17451 29597 17463 29631
rect 17405 29591 17463 29597
rect 17589 29631 17647 29637
rect 17589 29597 17601 29631
rect 17635 29628 17647 29631
rect 17770 29628 17776 29640
rect 17635 29600 17776 29628
rect 17635 29597 17647 29600
rect 17589 29591 17647 29597
rect 17420 29560 17448 29591
rect 17770 29588 17776 29600
rect 17828 29588 17834 29640
rect 18690 29628 18696 29640
rect 17972 29600 18696 29628
rect 17972 29560 18000 29600
rect 18690 29588 18696 29600
rect 18748 29588 18754 29640
rect 18877 29631 18935 29637
rect 18877 29597 18889 29631
rect 18923 29597 18935 29631
rect 23216 29628 23244 29659
rect 23658 29628 23664 29640
rect 23216 29600 23664 29628
rect 18877 29591 18935 29597
rect 17420 29532 18000 29560
rect 18049 29563 18107 29569
rect 18049 29529 18061 29563
rect 18095 29560 18107 29563
rect 18892 29560 18920 29591
rect 23658 29588 23664 29600
rect 23716 29628 23722 29640
rect 23860 29628 23888 29736
rect 25240 29708 25268 29736
rect 24394 29656 24400 29708
rect 24452 29656 24458 29708
rect 24489 29699 24547 29705
rect 24489 29665 24501 29699
rect 24535 29665 24547 29699
rect 24489 29659 24547 29665
rect 24581 29699 24639 29705
rect 24581 29665 24593 29699
rect 24627 29665 24639 29699
rect 24581 29659 24639 29665
rect 23716 29600 23888 29628
rect 24121 29631 24179 29637
rect 23716 29588 23722 29600
rect 24121 29597 24133 29631
rect 24167 29628 24179 29631
rect 24213 29631 24271 29637
rect 24213 29628 24225 29631
rect 24167 29600 24225 29628
rect 24167 29597 24179 29600
rect 24121 29591 24179 29597
rect 24213 29597 24225 29600
rect 24259 29597 24271 29631
rect 24213 29591 24271 29597
rect 18095 29532 18920 29560
rect 23293 29563 23351 29569
rect 18095 29529 18107 29532
rect 18049 29523 18107 29529
rect 23293 29529 23305 29563
rect 23339 29560 23351 29563
rect 24504 29560 24532 29659
rect 24596 29628 24624 29659
rect 24670 29656 24676 29708
rect 24728 29705 24734 29708
rect 24728 29699 24757 29705
rect 24745 29665 24757 29699
rect 24728 29659 24757 29665
rect 24728 29656 24734 29659
rect 25222 29656 25228 29708
rect 25280 29656 25286 29708
rect 25317 29699 25375 29705
rect 25317 29665 25329 29699
rect 25363 29696 25375 29699
rect 25593 29699 25651 29705
rect 25593 29696 25605 29699
rect 25363 29668 25605 29696
rect 25363 29665 25375 29668
rect 25317 29659 25375 29665
rect 25593 29665 25605 29668
rect 25639 29696 25651 29699
rect 25700 29696 25728 29792
rect 26050 29764 26056 29776
rect 25792 29736 26056 29764
rect 25792 29705 25820 29736
rect 26050 29724 26056 29736
rect 26108 29724 26114 29776
rect 28718 29764 28724 29776
rect 27370 29736 28724 29764
rect 28718 29724 28724 29736
rect 28776 29724 28782 29776
rect 28828 29764 28856 29795
rect 28994 29792 29000 29844
rect 29052 29792 29058 29844
rect 29270 29792 29276 29844
rect 29328 29832 29334 29844
rect 29730 29832 29736 29844
rect 29328 29804 29736 29832
rect 29328 29792 29334 29804
rect 29730 29792 29736 29804
rect 29788 29792 29794 29844
rect 29914 29792 29920 29844
rect 29972 29792 29978 29844
rect 30190 29792 30196 29844
rect 30248 29792 30254 29844
rect 29932 29764 29960 29792
rect 28828 29736 29960 29764
rect 31662 29724 31668 29776
rect 31720 29724 31726 29776
rect 25639 29668 25728 29696
rect 25777 29699 25835 29705
rect 25639 29665 25651 29668
rect 25593 29659 25651 29665
rect 25777 29665 25789 29699
rect 25823 29665 25835 29699
rect 28938 29699 28996 29705
rect 28938 29696 28950 29699
rect 25777 29659 25835 29665
rect 28000 29668 28950 29696
rect 28000 29640 28028 29668
rect 28938 29665 28950 29668
rect 28984 29665 28996 29699
rect 28938 29659 28996 29665
rect 29178 29656 29184 29708
rect 29236 29696 29242 29708
rect 29457 29699 29515 29705
rect 29457 29696 29469 29699
rect 29236 29668 29469 29696
rect 29236 29656 29242 29668
rect 29457 29665 29469 29668
rect 29503 29665 29515 29699
rect 29457 29659 29515 29665
rect 30285 29699 30343 29705
rect 30285 29665 30297 29699
rect 30331 29696 30343 29699
rect 30374 29696 30380 29708
rect 30331 29668 30380 29696
rect 30331 29665 30343 29668
rect 30285 29659 30343 29665
rect 30374 29656 30380 29668
rect 30432 29656 30438 29708
rect 30469 29699 30527 29705
rect 30469 29665 30481 29699
rect 30515 29665 30527 29699
rect 30469 29659 30527 29665
rect 24857 29631 24915 29637
rect 24596 29600 24808 29628
rect 24780 29572 24808 29600
rect 24857 29597 24869 29631
rect 24903 29628 24915 29631
rect 24949 29631 25007 29637
rect 24949 29628 24961 29631
rect 24903 29600 24961 29628
rect 24903 29597 24915 29600
rect 24857 29591 24915 29597
rect 24949 29597 24961 29600
rect 24995 29597 25007 29631
rect 24949 29591 25007 29597
rect 25869 29631 25927 29637
rect 25869 29597 25881 29631
rect 25915 29597 25927 29631
rect 25869 29591 25927 29597
rect 26145 29631 26203 29637
rect 26145 29597 26157 29631
rect 26191 29628 26203 29631
rect 27709 29631 27767 29637
rect 27709 29628 27721 29631
rect 26191 29600 27721 29628
rect 26191 29597 26203 29600
rect 26145 29591 26203 29597
rect 27709 29597 27721 29600
rect 27755 29597 27767 29631
rect 27709 29591 27767 29597
rect 23339 29532 24532 29560
rect 23339 29529 23351 29532
rect 23293 29523 23351 29529
rect 24762 29520 24768 29572
rect 24820 29520 24826 29572
rect 13504 29464 13676 29492
rect 13504 29452 13510 29464
rect 14366 29452 14372 29504
rect 14424 29452 14430 29504
rect 16850 29452 16856 29504
rect 16908 29452 16914 29504
rect 18322 29452 18328 29504
rect 18380 29452 18386 29504
rect 19150 29452 19156 29504
rect 19208 29452 19214 29504
rect 21542 29452 21548 29504
rect 21600 29452 21606 29504
rect 23750 29452 23756 29504
rect 23808 29492 23814 29504
rect 24872 29492 24900 29591
rect 23808 29464 24900 29492
rect 23808 29452 23814 29464
rect 24946 29452 24952 29504
rect 25004 29492 25010 29504
rect 25501 29495 25559 29501
rect 25501 29492 25513 29495
rect 25004 29464 25513 29492
rect 25004 29452 25010 29464
rect 25501 29461 25513 29464
rect 25547 29461 25559 29495
rect 25884 29492 25912 29591
rect 27982 29588 27988 29640
rect 28040 29588 28046 29640
rect 28350 29588 28356 29640
rect 28408 29588 28414 29640
rect 30484 29628 30512 29659
rect 28966 29600 30512 29628
rect 27154 29520 27160 29572
rect 27212 29560 27218 29572
rect 28966 29560 28994 29600
rect 27212 29532 28994 29560
rect 27212 29520 27218 29532
rect 26142 29492 26148 29504
rect 25884 29464 26148 29492
rect 25501 29455 25559 29461
rect 26142 29452 26148 29464
rect 26200 29452 26206 29504
rect 26234 29452 26240 29504
rect 26292 29492 26298 29504
rect 29270 29492 29276 29504
rect 26292 29464 29276 29492
rect 26292 29452 26298 29464
rect 29270 29452 29276 29464
rect 29328 29452 29334 29504
rect 29365 29495 29423 29501
rect 29365 29461 29377 29495
rect 29411 29492 29423 29495
rect 29546 29492 29552 29504
rect 29411 29464 29552 29492
rect 29411 29461 29423 29464
rect 29365 29455 29423 29461
rect 29546 29452 29552 29464
rect 29604 29452 29610 29504
rect 30009 29495 30067 29501
rect 30009 29461 30021 29495
rect 30055 29492 30067 29495
rect 31386 29492 31392 29504
rect 30055 29464 31392 29492
rect 30055 29461 30067 29464
rect 30009 29455 30067 29461
rect 31386 29452 31392 29464
rect 31444 29452 31450 29504
rect 2760 29402 32200 29424
rect 2760 29350 6286 29402
rect 6338 29350 6350 29402
rect 6402 29350 6414 29402
rect 6466 29350 6478 29402
rect 6530 29350 6542 29402
rect 6594 29350 13646 29402
rect 13698 29350 13710 29402
rect 13762 29350 13774 29402
rect 13826 29350 13838 29402
rect 13890 29350 13902 29402
rect 13954 29350 21006 29402
rect 21058 29350 21070 29402
rect 21122 29350 21134 29402
rect 21186 29350 21198 29402
rect 21250 29350 21262 29402
rect 21314 29350 28366 29402
rect 28418 29350 28430 29402
rect 28482 29350 28494 29402
rect 28546 29350 28558 29402
rect 28610 29350 28622 29402
rect 28674 29350 32200 29402
rect 2760 29328 32200 29350
rect 3513 29291 3571 29297
rect 3513 29257 3525 29291
rect 3559 29288 3571 29291
rect 3878 29288 3884 29300
rect 3559 29260 3884 29288
rect 3559 29257 3571 29260
rect 3513 29251 3571 29257
rect 3878 29248 3884 29260
rect 3936 29248 3942 29300
rect 8021 29291 8079 29297
rect 8021 29257 8033 29291
rect 8067 29288 8079 29291
rect 8294 29288 8300 29300
rect 8067 29260 8300 29288
rect 8067 29257 8079 29260
rect 8021 29251 8079 29257
rect 8294 29248 8300 29260
rect 8352 29248 8358 29300
rect 14366 29248 14372 29300
rect 14424 29248 14430 29300
rect 18322 29248 18328 29300
rect 18380 29248 18386 29300
rect 19705 29291 19763 29297
rect 19705 29257 19717 29291
rect 19751 29288 19763 29291
rect 20254 29288 20260 29300
rect 19751 29260 20260 29288
rect 19751 29257 19763 29260
rect 19705 29251 19763 29257
rect 20254 29248 20260 29260
rect 20312 29248 20318 29300
rect 21992 29291 22050 29297
rect 21992 29257 22004 29291
rect 22038 29288 22050 29291
rect 23569 29291 23627 29297
rect 23569 29288 23581 29291
rect 22038 29260 23581 29288
rect 22038 29257 22050 29260
rect 21992 29251 22050 29257
rect 23569 29257 23581 29260
rect 23615 29257 23627 29291
rect 26234 29288 26240 29300
rect 23569 29251 23627 29257
rect 23860 29260 26240 29288
rect 7745 29223 7803 29229
rect 7745 29189 7757 29223
rect 7791 29220 7803 29223
rect 8386 29220 8392 29232
rect 7791 29192 8392 29220
rect 7791 29189 7803 29192
rect 7745 29183 7803 29189
rect 8386 29180 8392 29192
rect 8444 29180 8450 29232
rect 11606 29220 11612 29232
rect 10888 29192 11612 29220
rect 5537 29155 5595 29161
rect 5537 29152 5549 29155
rect 3896 29124 5549 29152
rect 3896 29070 3924 29124
rect 5537 29121 5549 29124
rect 5583 29121 5595 29155
rect 8573 29155 8631 29161
rect 8573 29152 8585 29155
rect 5537 29115 5595 29121
rect 8312 29124 8585 29152
rect 5261 29087 5319 29093
rect 5261 29053 5273 29087
rect 5307 29053 5319 29087
rect 5261 29047 5319 29053
rect 5629 29087 5687 29093
rect 5629 29053 5641 29087
rect 5675 29053 5687 29087
rect 5629 29047 5687 29053
rect 4982 28976 4988 29028
rect 5040 28976 5046 29028
rect 4246 28908 4252 28960
rect 4304 28948 4310 28960
rect 5276 28948 5304 29047
rect 5644 29016 5672 29047
rect 7650 29044 7656 29096
rect 7708 29044 7714 29096
rect 6178 29016 6184 29028
rect 5644 28988 6184 29016
rect 6178 28976 6184 28988
rect 6236 29016 6242 29028
rect 7668 29016 7696 29044
rect 6236 28988 7696 29016
rect 6236 28976 6242 28988
rect 4304 28920 5304 28948
rect 4304 28908 4310 28920
rect 6822 28908 6828 28960
rect 6880 28948 6886 28960
rect 8312 28948 8340 29124
rect 8573 29121 8585 29124
rect 8619 29152 8631 29155
rect 9769 29155 9827 29161
rect 9769 29152 9781 29155
rect 8619 29124 9781 29152
rect 8619 29121 8631 29124
rect 8573 29115 8631 29121
rect 9769 29121 9781 29124
rect 9815 29152 9827 29155
rect 10778 29152 10784 29164
rect 9815 29124 10784 29152
rect 9815 29121 9827 29124
rect 9769 29115 9827 29121
rect 10778 29112 10784 29124
rect 10836 29152 10842 29164
rect 10888 29161 10916 29192
rect 11606 29180 11612 29192
rect 11664 29220 11670 29232
rect 11664 29192 12434 29220
rect 11664 29180 11670 29192
rect 10873 29155 10931 29161
rect 10873 29152 10885 29155
rect 10836 29124 10885 29152
rect 10836 29112 10842 29124
rect 10873 29121 10885 29124
rect 10919 29121 10931 29155
rect 10873 29115 10931 29121
rect 11146 29112 11152 29164
rect 11204 29152 11210 29164
rect 11882 29152 11888 29164
rect 11204 29124 11888 29152
rect 11204 29112 11210 29124
rect 11882 29112 11888 29124
rect 11940 29112 11946 29164
rect 12406 29152 12434 29192
rect 13173 29155 13231 29161
rect 13173 29152 13185 29155
rect 12406 29124 13185 29152
rect 13173 29121 13185 29124
rect 13219 29152 13231 29155
rect 14090 29152 14096 29164
rect 13219 29124 14096 29152
rect 13219 29121 13231 29124
rect 13173 29115 13231 29121
rect 14090 29112 14096 29124
rect 14148 29112 14154 29164
rect 14384 29152 14412 29248
rect 15381 29155 15439 29161
rect 15381 29152 15393 29155
rect 14384 29124 15393 29152
rect 15381 29121 15393 29124
rect 15427 29121 15439 29155
rect 15381 29115 15439 29121
rect 17313 29155 17371 29161
rect 17313 29121 17325 29155
rect 17359 29152 17371 29155
rect 18340 29152 18368 29248
rect 18690 29180 18696 29232
rect 18748 29220 18754 29232
rect 19521 29223 19579 29229
rect 19521 29220 19533 29223
rect 18748 29192 19533 29220
rect 18748 29180 18754 29192
rect 19521 29189 19533 29192
rect 19567 29220 19579 29223
rect 21542 29220 21548 29232
rect 19567 29192 21548 29220
rect 19567 29189 19579 29192
rect 19521 29183 19579 29189
rect 17359 29124 18368 29152
rect 17359 29121 17371 29124
rect 17313 29115 17371 29121
rect 18506 29112 18512 29164
rect 18564 29152 18570 29164
rect 20272 29161 20300 29192
rect 21542 29180 21548 29192
rect 21600 29180 21606 29232
rect 18785 29155 18843 29161
rect 18785 29152 18797 29155
rect 18564 29124 18797 29152
rect 18564 29112 18570 29124
rect 18785 29121 18797 29124
rect 18831 29152 18843 29155
rect 20257 29155 20315 29161
rect 18831 29124 20208 29152
rect 18831 29121 18843 29124
rect 18785 29115 18843 29121
rect 8389 29087 8447 29093
rect 8389 29053 8401 29087
rect 8435 29084 8447 29087
rect 8754 29084 8760 29096
rect 8435 29056 8760 29084
rect 8435 29053 8447 29056
rect 8389 29047 8447 29053
rect 8754 29044 8760 29056
rect 8812 29044 8818 29096
rect 8846 29044 8852 29096
rect 8904 29044 8910 29096
rect 11790 29044 11796 29096
rect 11848 29044 11854 29096
rect 12526 29044 12532 29096
rect 12584 29044 12590 29096
rect 13354 29044 13360 29096
rect 13412 29044 13418 29096
rect 14182 29044 14188 29096
rect 14240 29084 14246 29096
rect 14645 29087 14703 29093
rect 14645 29084 14657 29087
rect 14240 29056 14657 29084
rect 14240 29044 14246 29056
rect 14645 29053 14657 29056
rect 14691 29053 14703 29087
rect 14645 29047 14703 29053
rect 15933 29087 15991 29093
rect 15933 29053 15945 29087
rect 15979 29053 15991 29087
rect 15933 29047 15991 29053
rect 9493 29019 9551 29025
rect 9493 29016 9505 29019
rect 9232 28988 9505 29016
rect 6880 28920 8340 28948
rect 8481 28951 8539 28957
rect 6880 28908 6886 28920
rect 8481 28917 8493 28951
rect 8527 28948 8539 28951
rect 9232 28948 9260 28988
rect 9493 28985 9505 28988
rect 9539 29016 9551 29019
rect 9950 29016 9956 29028
rect 9539 28988 9956 29016
rect 9539 28985 9551 28988
rect 9493 28979 9551 28985
rect 9950 28976 9956 28988
rect 10008 28976 10014 29028
rect 11149 29019 11207 29025
rect 11149 28985 11161 29019
rect 11195 29016 11207 29019
rect 11238 29016 11244 29028
rect 11195 28988 11244 29016
rect 11195 28985 11207 28988
rect 11149 28979 11207 28985
rect 11238 28976 11244 28988
rect 11296 28976 11302 29028
rect 12434 28976 12440 29028
rect 12492 29016 12498 29028
rect 13538 29016 13544 29028
rect 12492 28988 13544 29016
rect 12492 28976 12498 28988
rect 13538 28976 13544 28988
rect 13596 29016 13602 29028
rect 14001 29019 14059 29025
rect 14001 29016 14013 29019
rect 13596 28988 14013 29016
rect 13596 28976 13602 28988
rect 14001 28985 14013 28988
rect 14047 28985 14059 29019
rect 14001 28979 14059 28985
rect 15948 28960 15976 29047
rect 16114 29044 16120 29096
rect 16172 29084 16178 29096
rect 16209 29087 16267 29093
rect 16209 29084 16221 29087
rect 16172 29056 16221 29084
rect 16172 29044 16178 29056
rect 16209 29053 16221 29056
rect 16255 29053 16267 29087
rect 16209 29047 16267 29053
rect 17034 29044 17040 29096
rect 17092 29044 17098 29096
rect 19150 29084 19156 29096
rect 18446 29056 19156 29084
rect 19150 29044 19156 29056
rect 19208 29044 19214 29096
rect 20180 29084 20208 29124
rect 20257 29121 20269 29155
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 21729 29155 21787 29161
rect 21729 29121 21741 29155
rect 21775 29152 21787 29155
rect 22094 29152 22100 29164
rect 21775 29124 22100 29152
rect 21775 29121 21787 29124
rect 21729 29115 21787 29121
rect 22094 29112 22100 29124
rect 22152 29112 22158 29164
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29152 23535 29155
rect 23750 29152 23756 29164
rect 23523 29124 23756 29152
rect 23523 29121 23535 29124
rect 23477 29115 23535 29121
rect 23750 29112 23756 29124
rect 23808 29112 23814 29164
rect 23860 29084 23888 29260
rect 26234 29248 26240 29260
rect 26292 29248 26298 29300
rect 26329 29291 26387 29297
rect 26329 29257 26341 29291
rect 26375 29257 26387 29291
rect 26329 29251 26387 29257
rect 24946 29180 24952 29232
rect 25004 29180 25010 29232
rect 26344 29220 26372 29251
rect 26786 29248 26792 29300
rect 26844 29288 26850 29300
rect 26881 29291 26939 29297
rect 26881 29288 26893 29291
rect 26844 29260 26893 29288
rect 26844 29248 26850 29260
rect 26881 29257 26893 29260
rect 26927 29257 26939 29291
rect 26881 29251 26939 29257
rect 27522 29248 27528 29300
rect 27580 29248 27586 29300
rect 27614 29248 27620 29300
rect 27672 29248 27678 29300
rect 28258 29248 28264 29300
rect 28316 29248 28322 29300
rect 28994 29248 29000 29300
rect 29052 29248 29058 29300
rect 29168 29291 29226 29297
rect 29168 29257 29180 29291
rect 29214 29288 29226 29291
rect 29362 29288 29368 29300
rect 29214 29260 29368 29288
rect 29214 29257 29226 29260
rect 29168 29251 29226 29257
rect 29362 29248 29368 29260
rect 29420 29248 29426 29300
rect 30650 29248 30656 29300
rect 30708 29248 30714 29300
rect 31294 29248 31300 29300
rect 31352 29248 31358 29300
rect 27540 29220 27568 29248
rect 25148 29192 26280 29220
rect 26344 29192 27568 29220
rect 27632 29220 27660 29248
rect 28353 29223 28411 29229
rect 28353 29220 28365 29223
rect 27632 29192 28365 29220
rect 24213 29155 24271 29161
rect 24213 29121 24225 29155
rect 24259 29152 24271 29155
rect 24964 29152 24992 29180
rect 25148 29164 25176 29192
rect 24259 29124 24992 29152
rect 24259 29121 24271 29124
rect 24213 29115 24271 29121
rect 25130 29112 25136 29164
rect 25188 29112 25194 29164
rect 25222 29112 25228 29164
rect 25280 29112 25286 29164
rect 26050 29112 26056 29164
rect 26108 29112 26114 29164
rect 20180 29056 20944 29084
rect 16850 28976 16856 29028
rect 16908 28976 16914 29028
rect 20073 29019 20131 29025
rect 20073 28985 20085 29019
rect 20119 29016 20131 29019
rect 20714 29016 20720 29028
rect 20119 28988 20720 29016
rect 20119 28985 20131 28988
rect 20073 28979 20131 28985
rect 20714 28976 20720 28988
rect 20772 28976 20778 29028
rect 20916 29016 20944 29056
rect 23492 29056 23888 29084
rect 24949 29087 25007 29093
rect 20916 28988 22416 29016
rect 8527 28920 9260 28948
rect 8527 28917 8539 28920
rect 8481 28911 8539 28917
rect 14090 28908 14096 28960
rect 14148 28908 14154 28960
rect 14642 28908 14648 28960
rect 14700 28948 14706 28960
rect 14829 28951 14887 28957
rect 14829 28948 14841 28951
rect 14700 28920 14841 28948
rect 14700 28908 14706 28920
rect 14829 28917 14841 28920
rect 14875 28917 14887 28951
rect 14829 28911 14887 28917
rect 15838 28908 15844 28960
rect 15896 28908 15902 28960
rect 15930 28908 15936 28960
rect 15988 28908 15994 28960
rect 20165 28951 20223 28957
rect 20165 28917 20177 28951
rect 20211 28948 20223 28951
rect 20438 28948 20444 28960
rect 20211 28920 20444 28948
rect 20211 28917 20223 28920
rect 20165 28911 20223 28917
rect 20438 28908 20444 28920
rect 20496 28908 20502 28960
rect 22388 28948 22416 28988
rect 22646 28976 22652 29028
rect 22704 28976 22710 29028
rect 23492 29016 23520 29056
rect 24949 29053 24961 29087
rect 24995 29053 25007 29087
rect 24949 29047 25007 29053
rect 25041 29087 25099 29093
rect 25041 29053 25053 29087
rect 25087 29084 25099 29087
rect 26068 29084 26096 29112
rect 26252 29093 26280 29192
rect 28353 29189 28365 29192
rect 28399 29189 28411 29223
rect 28353 29183 28411 29189
rect 26510 29112 26516 29164
rect 26568 29152 26574 29164
rect 27433 29155 27491 29161
rect 27433 29152 27445 29155
rect 26568 29124 27445 29152
rect 26568 29112 26574 29124
rect 27433 29121 27445 29124
rect 27479 29121 27491 29155
rect 27433 29115 27491 29121
rect 27893 29155 27951 29161
rect 27893 29121 27905 29155
rect 27939 29152 27951 29155
rect 28166 29152 28172 29164
rect 27939 29124 28172 29152
rect 27939 29121 27951 29124
rect 27893 29115 27951 29121
rect 28166 29112 28172 29124
rect 28224 29112 28230 29164
rect 29012 29152 29040 29248
rect 31312 29152 31340 29248
rect 28736 29124 29040 29152
rect 30300 29124 31340 29152
rect 25087 29056 26096 29084
rect 25087 29053 25099 29056
rect 25041 29047 25099 29053
rect 24029 29019 24087 29025
rect 24029 29016 24041 29019
rect 23308 28988 23520 29016
rect 23584 28988 24041 29016
rect 23308 28948 23336 28988
rect 23584 28960 23612 28988
rect 24029 28985 24041 28988
rect 24075 28985 24087 29019
rect 24964 29016 24992 29047
rect 25130 29016 25136 29028
rect 24964 28988 25136 29016
rect 24029 28979 24087 28985
rect 25130 28976 25136 28988
rect 25188 28976 25194 29028
rect 26068 29016 26096 29056
rect 26237 29087 26295 29093
rect 26237 29053 26249 29087
rect 26283 29053 26295 29087
rect 26237 29047 26295 29053
rect 26605 29087 26663 29093
rect 26605 29053 26617 29087
rect 26651 29053 26663 29087
rect 26605 29047 26663 29053
rect 26697 29087 26755 29093
rect 26697 29053 26709 29087
rect 26743 29053 26755 29087
rect 26697 29047 26755 29053
rect 26620 29016 26648 29047
rect 26068 28988 26648 29016
rect 26712 29016 26740 29047
rect 27614 29044 27620 29096
rect 27672 29084 27678 29096
rect 27801 29087 27859 29093
rect 27801 29084 27813 29087
rect 27672 29056 27813 29084
rect 27672 29044 27678 29056
rect 27801 29053 27813 29056
rect 27847 29053 27859 29087
rect 27801 29047 27859 29053
rect 27982 29044 27988 29096
rect 28040 29044 28046 29096
rect 28077 29087 28135 29093
rect 28077 29053 28089 29087
rect 28123 29084 28135 29087
rect 28626 29084 28632 29096
rect 28123 29056 28632 29084
rect 28123 29053 28135 29056
rect 28077 29047 28135 29053
rect 28626 29044 28632 29056
rect 28684 29084 28690 29096
rect 28736 29093 28764 29124
rect 28721 29087 28779 29093
rect 28721 29084 28733 29087
rect 28684 29056 28733 29084
rect 28684 29044 28690 29056
rect 28721 29053 28733 29056
rect 28767 29053 28779 29087
rect 28721 29047 28779 29053
rect 28902 29044 28908 29096
rect 28960 29044 28966 29096
rect 30300 29070 30328 29124
rect 31386 29112 31392 29164
rect 31444 29152 31450 29164
rect 31444 29124 31708 29152
rect 31444 29112 31450 29124
rect 30926 29044 30932 29096
rect 30984 29044 30990 29096
rect 31680 29093 31708 29124
rect 31665 29087 31723 29093
rect 31665 29053 31677 29087
rect 31711 29053 31723 29087
rect 31665 29047 31723 29053
rect 27890 29016 27896 29028
rect 26712 28988 27896 29016
rect 22388 28920 23336 28948
rect 23566 28908 23572 28960
rect 23624 28908 23630 28960
rect 23934 28908 23940 28960
rect 23992 28908 23998 28960
rect 26050 28908 26056 28960
rect 26108 28908 26114 28960
rect 26418 28908 26424 28960
rect 26476 28948 26482 28960
rect 26712 28948 26740 28988
rect 27890 28976 27896 28988
rect 27948 29016 27954 29028
rect 28537 29019 28595 29025
rect 28537 29016 28549 29019
rect 27948 28988 28549 29016
rect 27948 28976 27954 28988
rect 28537 28985 28549 28988
rect 28583 28985 28595 29019
rect 28537 28979 28595 28985
rect 30760 28988 30972 29016
rect 26476 28920 26740 28948
rect 26476 28908 26482 28920
rect 26878 28908 26884 28960
rect 26936 28948 26942 28960
rect 30006 28948 30012 28960
rect 26936 28920 30012 28948
rect 26936 28908 26942 28920
rect 30006 28908 30012 28920
rect 30064 28948 30070 28960
rect 30760 28948 30788 28988
rect 30064 28920 30788 28948
rect 30064 28908 30070 28920
rect 30834 28908 30840 28960
rect 30892 28908 30898 28960
rect 30944 28948 30972 28988
rect 31294 28976 31300 29028
rect 31352 29016 31358 29028
rect 31389 29019 31447 29025
rect 31389 29016 31401 29019
rect 31352 28988 31401 29016
rect 31352 28976 31358 28988
rect 31389 28985 31401 28988
rect 31435 28985 31447 29019
rect 31389 28979 31447 28985
rect 31662 28948 31668 28960
rect 30944 28920 31668 28948
rect 31662 28908 31668 28920
rect 31720 28908 31726 28960
rect 2760 28858 32200 28880
rect 2760 28806 6946 28858
rect 6998 28806 7010 28858
rect 7062 28806 7074 28858
rect 7126 28806 7138 28858
rect 7190 28806 7202 28858
rect 7254 28806 14306 28858
rect 14358 28806 14370 28858
rect 14422 28806 14434 28858
rect 14486 28806 14498 28858
rect 14550 28806 14562 28858
rect 14614 28806 21666 28858
rect 21718 28806 21730 28858
rect 21782 28806 21794 28858
rect 21846 28806 21858 28858
rect 21910 28806 21922 28858
rect 21974 28806 29026 28858
rect 29078 28806 29090 28858
rect 29142 28806 29154 28858
rect 29206 28806 29218 28858
rect 29270 28806 29282 28858
rect 29334 28806 32200 28858
rect 2760 28784 32200 28806
rect 8021 28747 8079 28753
rect 8021 28713 8033 28747
rect 8067 28744 8079 28747
rect 8846 28744 8852 28756
rect 8067 28716 8852 28744
rect 8067 28713 8079 28716
rect 8021 28707 8079 28713
rect 8846 28704 8852 28716
rect 8904 28704 8910 28756
rect 12526 28704 12532 28756
rect 12584 28744 12590 28756
rect 12621 28747 12679 28753
rect 12621 28744 12633 28747
rect 12584 28716 12633 28744
rect 12584 28704 12590 28716
rect 12621 28713 12633 28716
rect 12667 28713 12679 28747
rect 12621 28707 12679 28713
rect 14642 28704 14648 28756
rect 14700 28704 14706 28756
rect 15746 28704 15752 28756
rect 15804 28704 15810 28756
rect 22646 28704 22652 28756
rect 22704 28704 22710 28756
rect 23566 28704 23572 28756
rect 23624 28704 23630 28756
rect 23934 28704 23940 28756
rect 23992 28744 23998 28756
rect 24581 28747 24639 28753
rect 24581 28744 24593 28747
rect 23992 28716 24593 28744
rect 23992 28704 23998 28716
rect 24581 28713 24593 28716
rect 24627 28713 24639 28747
rect 24581 28707 24639 28713
rect 26973 28747 27031 28753
rect 26973 28713 26985 28747
rect 27019 28744 27031 28747
rect 27062 28744 27068 28756
rect 27019 28716 27068 28744
rect 27019 28713 27031 28716
rect 26973 28707 27031 28713
rect 27062 28704 27068 28716
rect 27120 28704 27126 28756
rect 27522 28744 27528 28756
rect 27356 28716 27528 28744
rect 5258 28636 5264 28688
rect 5316 28636 5322 28688
rect 12805 28679 12863 28685
rect 12805 28676 12817 28679
rect 12374 28648 12817 28676
rect 12805 28645 12817 28648
rect 12851 28645 12863 28679
rect 12805 28639 12863 28645
rect 14277 28679 14335 28685
rect 14277 28645 14289 28679
rect 14323 28676 14335 28679
rect 14660 28676 14688 28704
rect 15838 28676 15844 28688
rect 14323 28648 14688 28676
rect 15502 28648 15844 28676
rect 14323 28645 14335 28648
rect 14277 28639 14335 28645
rect 15838 28636 15844 28648
rect 15896 28636 15902 28688
rect 20346 28636 20352 28688
rect 20404 28676 20410 28688
rect 21358 28676 21364 28688
rect 20404 28648 21364 28676
rect 20404 28636 20410 28648
rect 21358 28636 21364 28648
rect 21416 28676 21422 28688
rect 23474 28676 23480 28688
rect 21416 28648 23480 28676
rect 21416 28636 21422 28648
rect 23474 28636 23480 28648
rect 23532 28636 23538 28688
rect 6457 28611 6515 28617
rect 6457 28608 6469 28611
rect 5736 28580 6469 28608
rect 3973 28543 4031 28549
rect 3973 28509 3985 28543
rect 4019 28509 4031 28543
rect 3973 28503 4031 28509
rect 4249 28543 4307 28549
rect 4249 28509 4261 28543
rect 4295 28540 4307 28543
rect 5442 28540 5448 28552
rect 4295 28512 5448 28540
rect 4295 28509 4307 28512
rect 4249 28503 4307 28509
rect 3988 28404 4016 28503
rect 5442 28500 5448 28512
rect 5500 28500 5506 28552
rect 5736 28549 5764 28580
rect 6457 28577 6469 28580
rect 6503 28608 6515 28611
rect 6638 28608 6644 28620
rect 6503 28580 6644 28608
rect 6503 28577 6515 28580
rect 6457 28571 6515 28577
rect 6638 28568 6644 28580
rect 6696 28568 6702 28620
rect 8386 28568 8392 28620
rect 8444 28568 8450 28620
rect 10870 28608 10876 28620
rect 9784 28580 10876 28608
rect 5721 28543 5779 28549
rect 5721 28509 5733 28543
rect 5767 28509 5779 28543
rect 5721 28503 5779 28509
rect 7193 28543 7251 28549
rect 7193 28509 7205 28543
rect 7239 28509 7251 28543
rect 7193 28503 7251 28509
rect 6638 28432 6644 28484
rect 6696 28472 6702 28484
rect 7208 28472 7236 28503
rect 9490 28500 9496 28552
rect 9548 28500 9554 28552
rect 9784 28549 9812 28580
rect 10870 28568 10876 28580
rect 10928 28568 10934 28620
rect 12894 28568 12900 28620
rect 12952 28568 12958 28620
rect 15930 28568 15936 28620
rect 15988 28608 15994 28620
rect 16025 28611 16083 28617
rect 16025 28608 16037 28611
rect 15988 28580 16037 28608
rect 15988 28568 15994 28580
rect 16025 28577 16037 28580
rect 16071 28608 16083 28611
rect 16301 28611 16359 28617
rect 16301 28608 16313 28611
rect 16071 28580 16313 28608
rect 16071 28577 16083 28580
rect 16025 28571 16083 28577
rect 16301 28577 16313 28580
rect 16347 28577 16359 28611
rect 16301 28571 16359 28577
rect 22094 28568 22100 28620
rect 22152 28608 22158 28620
rect 22554 28608 22560 28620
rect 22152 28580 22560 28608
rect 22152 28568 22158 28580
rect 22554 28568 22560 28580
rect 22612 28568 22618 28620
rect 9769 28543 9827 28549
rect 9769 28540 9781 28543
rect 9692 28512 9781 28540
rect 6696 28444 7236 28472
rect 6696 28432 6702 28444
rect 9692 28416 9720 28512
rect 9769 28509 9781 28512
rect 9815 28509 9827 28543
rect 9769 28503 9827 28509
rect 10226 28500 10232 28552
rect 10284 28500 10290 28552
rect 10781 28543 10839 28549
rect 10781 28509 10793 28543
rect 10827 28540 10839 28543
rect 11149 28543 11207 28549
rect 11149 28540 11161 28543
rect 10827 28512 11161 28540
rect 10827 28509 10839 28512
rect 10781 28503 10839 28509
rect 11149 28509 11161 28512
rect 11195 28509 11207 28543
rect 11149 28503 11207 28509
rect 13998 28500 14004 28552
rect 14056 28500 14062 28552
rect 17126 28500 17132 28552
rect 17184 28500 17190 28552
rect 19794 28500 19800 28552
rect 19852 28500 19858 28552
rect 23584 28540 23612 28704
rect 24026 28676 24032 28688
rect 23676 28648 24032 28676
rect 23676 28617 23704 28648
rect 24026 28636 24032 28648
rect 24084 28676 24090 28688
rect 27356 28685 27384 28716
rect 27522 28704 27528 28716
rect 27580 28704 27586 28756
rect 28626 28704 28632 28756
rect 28684 28704 28690 28756
rect 28997 28747 29055 28753
rect 28997 28713 29009 28747
rect 29043 28744 29055 28747
rect 31021 28747 31079 28753
rect 31021 28744 31033 28747
rect 29043 28716 31033 28744
rect 29043 28713 29055 28716
rect 28997 28707 29055 28713
rect 31021 28713 31033 28716
rect 31067 28744 31079 28747
rect 31110 28744 31116 28756
rect 31067 28716 31116 28744
rect 31067 28713 31079 28716
rect 31021 28707 31079 28713
rect 31110 28704 31116 28716
rect 31168 28704 31174 28756
rect 24397 28679 24455 28685
rect 24397 28676 24409 28679
rect 24084 28648 24409 28676
rect 24084 28636 24090 28648
rect 24397 28645 24409 28648
rect 24443 28645 24455 28679
rect 24397 28639 24455 28645
rect 27157 28679 27215 28685
rect 27157 28645 27169 28679
rect 27203 28645 27215 28679
rect 27157 28639 27215 28645
rect 27341 28679 27399 28685
rect 27341 28645 27353 28679
rect 27387 28645 27399 28679
rect 27341 28639 27399 28645
rect 27448 28648 28120 28676
rect 23661 28611 23719 28617
rect 23661 28577 23673 28611
rect 23707 28577 23719 28611
rect 23661 28571 23719 28577
rect 23750 28568 23756 28620
rect 23808 28568 23814 28620
rect 24489 28611 24547 28617
rect 24489 28577 24501 28611
rect 24535 28577 24547 28611
rect 24489 28571 24547 28577
rect 24673 28611 24731 28617
rect 24673 28577 24685 28611
rect 24719 28608 24731 28611
rect 25130 28608 25136 28620
rect 24719 28580 25136 28608
rect 24719 28577 24731 28580
rect 24673 28571 24731 28577
rect 24504 28540 24532 28571
rect 25130 28568 25136 28580
rect 25188 28608 25194 28620
rect 27172 28608 27200 28639
rect 27448 28608 27476 28648
rect 25188 28580 27108 28608
rect 27172 28580 27476 28608
rect 25188 28568 25194 28580
rect 23584 28512 24532 28540
rect 26970 28500 26976 28552
rect 27028 28500 27034 28552
rect 27080 28540 27108 28580
rect 27522 28568 27528 28620
rect 27580 28568 27586 28620
rect 27617 28611 27675 28617
rect 27617 28577 27629 28611
rect 27663 28608 27675 28611
rect 27706 28608 27712 28620
rect 27663 28580 27712 28608
rect 27663 28577 27675 28580
rect 27617 28571 27675 28577
rect 27706 28568 27712 28580
rect 27764 28568 27770 28620
rect 27801 28611 27859 28617
rect 27801 28577 27813 28611
rect 27847 28577 27859 28611
rect 27801 28571 27859 28577
rect 27540 28540 27568 28568
rect 27080 28512 27568 28540
rect 26988 28472 27016 28500
rect 26988 28444 27292 28472
rect 4246 28404 4252 28416
rect 3988 28376 4252 28404
rect 4246 28364 4252 28376
rect 4304 28364 4310 28416
rect 5810 28364 5816 28416
rect 5868 28364 5874 28416
rect 7834 28364 7840 28416
rect 7892 28364 7898 28416
rect 9674 28364 9680 28416
rect 9732 28364 9738 28416
rect 13909 28407 13967 28413
rect 13909 28373 13921 28407
rect 13955 28404 13967 28407
rect 14642 28404 14648 28416
rect 13955 28376 14648 28404
rect 13955 28373 13967 28376
rect 13909 28367 13967 28373
rect 14642 28364 14648 28376
rect 14700 28364 14706 28416
rect 15933 28407 15991 28413
rect 15933 28373 15945 28407
rect 15979 28404 15991 28407
rect 16022 28404 16028 28416
rect 15979 28376 16028 28404
rect 15979 28373 15991 28376
rect 15933 28367 15991 28373
rect 16022 28364 16028 28376
rect 16080 28364 16086 28416
rect 16206 28364 16212 28416
rect 16264 28364 16270 28416
rect 16574 28364 16580 28416
rect 16632 28364 16638 28416
rect 17770 28364 17776 28416
rect 17828 28364 17834 28416
rect 20438 28364 20444 28416
rect 20496 28364 20502 28416
rect 26418 28364 26424 28416
rect 26476 28404 26482 28416
rect 27157 28407 27215 28413
rect 27157 28404 27169 28407
rect 26476 28376 27169 28404
rect 26476 28364 26482 28376
rect 27157 28373 27169 28376
rect 27203 28373 27215 28407
rect 27264 28404 27292 28444
rect 27430 28432 27436 28484
rect 27488 28472 27494 28484
rect 27525 28475 27583 28481
rect 27525 28472 27537 28475
rect 27488 28444 27537 28472
rect 27488 28432 27494 28444
rect 27525 28441 27537 28444
rect 27571 28441 27583 28475
rect 27816 28472 27844 28571
rect 27890 28568 27896 28620
rect 27948 28568 27954 28620
rect 28092 28617 28120 28648
rect 28077 28611 28135 28617
rect 28077 28577 28089 28611
rect 28123 28608 28135 28611
rect 28644 28608 28672 28704
rect 28905 28679 28963 28685
rect 28905 28676 28917 28679
rect 28123 28580 28672 28608
rect 28736 28648 28917 28676
rect 28123 28577 28135 28580
rect 28077 28571 28135 28577
rect 28166 28500 28172 28552
rect 28224 28540 28230 28552
rect 28736 28540 28764 28648
rect 28905 28645 28917 28648
rect 28951 28645 28963 28679
rect 28905 28639 28963 28645
rect 29181 28679 29239 28685
rect 29181 28645 29193 28679
rect 29227 28676 29239 28679
rect 29546 28676 29552 28688
rect 29227 28648 29552 28676
rect 29227 28645 29239 28648
rect 29181 28639 29239 28645
rect 29546 28636 29552 28648
rect 29604 28636 29610 28688
rect 30834 28676 30840 28688
rect 30774 28648 30840 28676
rect 30834 28636 30840 28648
rect 30892 28636 30898 28688
rect 31662 28636 31668 28688
rect 31720 28636 31726 28688
rect 28810 28568 28816 28620
rect 28868 28568 28874 28620
rect 31389 28611 31447 28617
rect 31389 28577 31401 28611
rect 31435 28577 31447 28611
rect 31389 28571 31447 28577
rect 28224 28512 28764 28540
rect 28224 28500 28230 28512
rect 28902 28500 28908 28552
rect 28960 28540 28966 28552
rect 29273 28543 29331 28549
rect 29273 28540 29285 28543
rect 28960 28512 29285 28540
rect 28960 28500 28966 28512
rect 29273 28509 29285 28512
rect 29319 28509 29331 28543
rect 29273 28503 29331 28509
rect 29549 28543 29607 28549
rect 29549 28509 29561 28543
rect 29595 28540 29607 28543
rect 29595 28512 31156 28540
rect 29595 28509 29607 28512
rect 29549 28503 29607 28509
rect 29178 28472 29184 28484
rect 27816 28444 29184 28472
rect 27525 28435 27583 28441
rect 29178 28432 29184 28444
rect 29236 28432 29242 28484
rect 31128 28481 31156 28512
rect 31202 28500 31208 28552
rect 31260 28540 31266 28552
rect 31297 28543 31355 28549
rect 31297 28540 31309 28543
rect 31260 28512 31309 28540
rect 31260 28500 31266 28512
rect 31297 28509 31309 28512
rect 31343 28509 31355 28543
rect 31297 28503 31355 28509
rect 31113 28475 31171 28481
rect 31113 28441 31125 28475
rect 31159 28441 31171 28475
rect 31113 28435 31171 28441
rect 27985 28407 28043 28413
rect 27985 28404 27997 28407
rect 27264 28376 27997 28404
rect 27157 28367 27215 28373
rect 27985 28373 27997 28376
rect 28031 28373 28043 28407
rect 27985 28367 28043 28373
rect 30190 28364 30196 28416
rect 30248 28404 30254 28416
rect 31404 28404 31432 28571
rect 31757 28543 31815 28549
rect 31757 28509 31769 28543
rect 31803 28540 31815 28543
rect 31803 28512 32260 28540
rect 31803 28509 31815 28512
rect 31757 28503 31815 28509
rect 30248 28376 31432 28404
rect 30248 28364 30254 28376
rect 2760 28314 32200 28336
rect 2760 28262 6286 28314
rect 6338 28262 6350 28314
rect 6402 28262 6414 28314
rect 6466 28262 6478 28314
rect 6530 28262 6542 28314
rect 6594 28262 13646 28314
rect 13698 28262 13710 28314
rect 13762 28262 13774 28314
rect 13826 28262 13838 28314
rect 13890 28262 13902 28314
rect 13954 28262 21006 28314
rect 21058 28262 21070 28314
rect 21122 28262 21134 28314
rect 21186 28262 21198 28314
rect 21250 28262 21262 28314
rect 21314 28262 28366 28314
rect 28418 28262 28430 28314
rect 28482 28262 28494 28314
rect 28546 28262 28558 28314
rect 28610 28262 28622 28314
rect 28674 28262 32200 28314
rect 2760 28240 32200 28262
rect 4982 28160 4988 28212
rect 5040 28200 5046 28212
rect 5261 28203 5319 28209
rect 5261 28200 5273 28203
rect 5040 28172 5273 28200
rect 5040 28160 5046 28172
rect 5261 28169 5273 28172
rect 5307 28169 5319 28203
rect 5261 28163 5319 28169
rect 5442 28160 5448 28212
rect 5500 28160 5506 28212
rect 5810 28160 5816 28212
rect 5868 28160 5874 28212
rect 9309 28203 9367 28209
rect 9309 28169 9321 28203
rect 9355 28200 9367 28203
rect 9490 28200 9496 28212
rect 9355 28172 9496 28200
rect 9355 28169 9367 28172
rect 9309 28163 9367 28169
rect 9490 28160 9496 28172
rect 9548 28160 9554 28212
rect 10226 28160 10232 28212
rect 10284 28200 10290 28212
rect 10689 28203 10747 28209
rect 10689 28200 10701 28203
rect 10284 28172 10701 28200
rect 10284 28160 10290 28172
rect 10689 28169 10701 28172
rect 10735 28169 10747 28203
rect 12066 28200 12072 28212
rect 10689 28163 10747 28169
rect 10796 28172 12072 28200
rect 3878 28024 3884 28076
rect 3936 28024 3942 28076
rect 4709 28067 4767 28073
rect 4709 28033 4721 28067
rect 4755 28064 4767 28067
rect 4755 28036 5580 28064
rect 4755 28033 4767 28036
rect 4709 28027 4767 28033
rect 5552 27940 5580 28036
rect 5828 28005 5856 28160
rect 10796 28132 10824 28172
rect 12066 28160 12072 28172
rect 12124 28200 12130 28212
rect 12894 28200 12900 28212
rect 12124 28172 12900 28200
rect 12124 28160 12130 28172
rect 12894 28160 12900 28172
rect 12952 28200 12958 28212
rect 13081 28203 13139 28209
rect 12952 28172 13032 28200
rect 12952 28160 12958 28172
rect 5920 28104 7420 28132
rect 5920 28005 5948 28104
rect 5997 28067 6055 28073
rect 5997 28033 6009 28067
rect 6043 28033 6055 28067
rect 7392 28064 7420 28104
rect 10428 28104 10824 28132
rect 7392 28036 10364 28064
rect 5997 28027 6055 28033
rect 5813 27999 5871 28005
rect 5813 27965 5825 27999
rect 5859 27965 5871 27999
rect 5813 27959 5871 27965
rect 5905 27999 5963 28005
rect 5905 27965 5917 27999
rect 5951 27965 5963 27999
rect 5905 27959 5963 27965
rect 4433 27931 4491 27937
rect 4433 27897 4445 27931
rect 4479 27928 4491 27931
rect 4893 27931 4951 27937
rect 4893 27928 4905 27931
rect 4479 27900 4905 27928
rect 4479 27897 4491 27900
rect 4433 27891 4491 27897
rect 4893 27897 4905 27900
rect 4939 27897 4951 27931
rect 4893 27891 4951 27897
rect 5534 27888 5540 27940
rect 5592 27928 5598 27940
rect 6012 27928 6040 28027
rect 7285 27999 7343 28005
rect 7285 27965 7297 27999
rect 7331 27965 7343 27999
rect 7285 27959 7343 27965
rect 6457 27931 6515 27937
rect 6457 27928 6469 27931
rect 5592 27900 6469 27928
rect 5592 27888 5598 27900
rect 6457 27897 6469 27900
rect 6503 27928 6515 27931
rect 6822 27928 6828 27940
rect 6503 27900 6828 27928
rect 6503 27897 6515 27900
rect 6457 27891 6515 27897
rect 6822 27888 6828 27900
rect 6880 27888 6886 27940
rect 7300 27928 7328 27959
rect 9858 27956 9864 28008
rect 9916 27956 9922 28008
rect 7561 27931 7619 27937
rect 7300 27900 7420 27928
rect 7392 27872 7420 27900
rect 7561 27897 7573 27931
rect 7607 27928 7619 27931
rect 7834 27928 7840 27940
rect 7607 27900 7840 27928
rect 7607 27897 7619 27900
rect 7561 27891 7619 27897
rect 7834 27888 7840 27900
rect 7892 27888 7898 27940
rect 9766 27928 9772 27940
rect 8786 27900 9772 27928
rect 9766 27888 9772 27900
rect 9824 27888 9830 27940
rect 10336 27928 10364 28036
rect 10428 28005 10456 28104
rect 10870 28092 10876 28144
rect 10928 28092 10934 28144
rect 10888 28064 10916 28092
rect 11333 28067 11391 28073
rect 11333 28064 11345 28067
rect 10888 28036 11345 28064
rect 11333 28033 11345 28036
rect 11379 28033 11391 28067
rect 11333 28027 11391 28033
rect 10413 27999 10471 28005
rect 10413 27965 10425 27999
rect 10459 27965 10471 27999
rect 10413 27959 10471 27965
rect 10594 27956 10600 28008
rect 10652 27996 10658 28008
rect 10873 27999 10931 28005
rect 10873 27996 10885 27999
rect 10652 27968 10885 27996
rect 10652 27956 10658 27968
rect 10873 27965 10885 27968
rect 10919 27965 10931 27999
rect 10873 27959 10931 27965
rect 10965 27999 11023 28005
rect 10965 27965 10977 27999
rect 11011 27996 11023 27999
rect 11146 27996 11152 28008
rect 11011 27968 11152 27996
rect 11011 27965 11023 27968
rect 10965 27959 11023 27965
rect 11146 27956 11152 27968
rect 11204 27956 11210 28008
rect 11241 27999 11299 28005
rect 11241 27965 11253 27999
rect 11287 27996 11299 27999
rect 13004 27996 13032 28172
rect 13081 28169 13093 28203
rect 13127 28200 13139 28203
rect 13354 28200 13360 28212
rect 13127 28172 13360 28200
rect 13127 28169 13139 28172
rect 13081 28163 13139 28169
rect 13354 28160 13360 28172
rect 13412 28160 13418 28212
rect 15565 28203 15623 28209
rect 13556 28172 15148 28200
rect 13556 28008 13584 28172
rect 14090 28024 14096 28076
rect 14148 28024 14154 28076
rect 15120 28064 15148 28172
rect 15565 28169 15577 28203
rect 15611 28200 15623 28203
rect 16114 28200 16120 28212
rect 15611 28172 16120 28200
rect 15611 28169 15623 28172
rect 15565 28163 15623 28169
rect 16114 28160 16120 28172
rect 16172 28160 16178 28212
rect 19429 28203 19487 28209
rect 19429 28169 19441 28203
rect 19475 28200 19487 28203
rect 19794 28200 19800 28212
rect 19475 28172 19800 28200
rect 19475 28169 19487 28172
rect 19429 28163 19487 28169
rect 19794 28160 19800 28172
rect 19852 28160 19858 28212
rect 23842 28160 23848 28212
rect 23900 28200 23906 28212
rect 23937 28203 23995 28209
rect 23937 28200 23949 28203
rect 23900 28172 23949 28200
rect 23900 28160 23906 28172
rect 23937 28169 23949 28172
rect 23983 28169 23995 28203
rect 23937 28163 23995 28169
rect 24026 28160 24032 28212
rect 24084 28160 24090 28212
rect 26513 28203 26571 28209
rect 26513 28169 26525 28203
rect 26559 28200 26571 28203
rect 26602 28200 26608 28212
rect 26559 28172 26608 28200
rect 26559 28169 26571 28172
rect 26513 28163 26571 28169
rect 26602 28160 26608 28172
rect 26660 28160 26666 28212
rect 28534 28160 28540 28212
rect 28592 28200 28598 28212
rect 28718 28200 28724 28212
rect 28592 28172 28724 28200
rect 28592 28160 28598 28172
rect 28718 28160 28724 28172
rect 28776 28160 28782 28212
rect 28810 28160 28816 28212
rect 28868 28160 28874 28212
rect 29454 28160 29460 28212
rect 29512 28200 29518 28212
rect 29825 28203 29883 28209
rect 29825 28200 29837 28203
rect 29512 28172 29837 28200
rect 29512 28160 29518 28172
rect 29825 28169 29837 28172
rect 29871 28200 29883 28203
rect 30190 28200 30196 28212
rect 29871 28172 30196 28200
rect 29871 28169 29883 28172
rect 29825 28163 29883 28169
rect 30190 28160 30196 28172
rect 30248 28160 30254 28212
rect 30374 28160 30380 28212
rect 30432 28200 30438 28212
rect 30837 28203 30895 28209
rect 30837 28200 30849 28203
rect 30432 28172 30849 28200
rect 30432 28160 30438 28172
rect 30837 28169 30849 28172
rect 30883 28169 30895 28203
rect 30837 28163 30895 28169
rect 31021 28203 31079 28209
rect 31021 28169 31033 28203
rect 31067 28200 31079 28203
rect 32232 28200 32260 28512
rect 31067 28172 32260 28200
rect 31067 28169 31079 28172
rect 31021 28163 31079 28169
rect 15841 28067 15899 28073
rect 15841 28064 15853 28067
rect 15120 28036 15853 28064
rect 15841 28033 15853 28036
rect 15887 28064 15899 28067
rect 15930 28064 15936 28076
rect 15887 28036 15936 28064
rect 15887 28033 15899 28036
rect 15841 28027 15899 28033
rect 15930 28024 15936 28036
rect 15988 28024 15994 28076
rect 17034 28024 17040 28076
rect 17092 28064 17098 28076
rect 17681 28067 17739 28073
rect 17681 28064 17693 28067
rect 17092 28036 17693 28064
rect 17092 28024 17098 28036
rect 17681 28033 17693 28036
rect 17727 28033 17739 28067
rect 17681 28027 17739 28033
rect 13357 27999 13415 28005
rect 13357 27996 13369 27999
rect 11287 27968 11376 27996
rect 13004 27968 13369 27996
rect 11287 27965 11299 27968
rect 11241 27959 11299 27965
rect 10502 27928 10508 27940
rect 10336 27900 10508 27928
rect 10502 27888 10508 27900
rect 10560 27888 10566 27940
rect 11054 27888 11060 27940
rect 11112 27888 11118 27940
rect 4801 27863 4859 27869
rect 4801 27829 4813 27863
rect 4847 27860 4859 27863
rect 6546 27860 6552 27872
rect 4847 27832 6552 27860
rect 4847 27829 4859 27832
rect 4801 27823 4859 27829
rect 6546 27820 6552 27832
rect 6604 27820 6610 27872
rect 7193 27863 7251 27869
rect 7193 27829 7205 27863
rect 7239 27860 7251 27863
rect 7282 27860 7288 27872
rect 7239 27832 7288 27860
rect 7239 27829 7251 27832
rect 7193 27823 7251 27829
rect 7282 27820 7288 27832
rect 7340 27820 7346 27872
rect 7374 27820 7380 27872
rect 7432 27820 7438 27872
rect 9030 27820 9036 27872
rect 9088 27820 9094 27872
rect 10318 27820 10324 27872
rect 10376 27820 10382 27872
rect 11348 27860 11376 27968
rect 13357 27965 13369 27968
rect 13403 27996 13415 27999
rect 13538 27996 13544 28008
rect 13403 27968 13544 27996
rect 13403 27965 13415 27968
rect 13357 27959 13415 27965
rect 13538 27956 13544 27968
rect 13596 27956 13602 28008
rect 13817 27999 13875 28005
rect 13817 27965 13829 27999
rect 13863 27965 13875 27999
rect 16206 27996 16212 28008
rect 15226 27968 16212 27996
rect 13817 27959 13875 27965
rect 11606 27888 11612 27940
rect 11664 27888 11670 27940
rect 13265 27931 13323 27937
rect 13265 27928 13277 27931
rect 12834 27900 13277 27928
rect 13265 27897 13277 27900
rect 13311 27897 13323 27931
rect 13832 27928 13860 27959
rect 16206 27956 16212 27968
rect 16264 27956 16270 28008
rect 19702 27956 19708 28008
rect 19760 27996 19766 28008
rect 22094 27996 22100 28008
rect 19760 27968 22100 27996
rect 19760 27956 19766 27968
rect 22094 27956 22100 27968
rect 22152 27956 22158 28008
rect 23106 27956 23112 28008
rect 23164 27996 23170 28008
rect 23566 28005 23572 28008
rect 23293 27999 23351 28005
rect 23293 27996 23305 27999
rect 23164 27968 23305 27996
rect 23164 27956 23170 27968
rect 23293 27965 23305 27968
rect 23339 27965 23351 27999
rect 23293 27959 23351 27965
rect 23551 27999 23572 28005
rect 23551 27965 23563 27999
rect 23551 27959 23572 27965
rect 23566 27956 23572 27959
rect 23624 27956 23630 28008
rect 23658 27956 23664 28008
rect 23716 27956 23722 28008
rect 24044 28005 24072 28160
rect 24486 28092 24492 28144
rect 24544 28132 24550 28144
rect 24544 28104 24716 28132
rect 24544 28092 24550 28104
rect 24688 28073 24716 28104
rect 27614 28092 27620 28144
rect 27672 28092 27678 28144
rect 28258 28092 28264 28144
rect 28316 28092 28322 28144
rect 24673 28067 24731 28073
rect 24673 28033 24685 28067
rect 24719 28033 24731 28067
rect 24673 28027 24731 28033
rect 24765 28067 24823 28073
rect 24765 28033 24777 28067
rect 24811 28064 24823 28067
rect 24811 28036 25176 28064
rect 24811 28033 24823 28036
rect 24765 28027 24823 28033
rect 25148 28008 25176 28036
rect 26050 28024 26056 28076
rect 26108 28024 26114 28076
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28064 26295 28067
rect 27525 28067 27583 28073
rect 27525 28064 27537 28067
rect 26283 28036 27537 28064
rect 26283 28033 26295 28036
rect 26237 28027 26295 28033
rect 27525 28033 27537 28036
rect 27571 28033 27583 28067
rect 27632 28064 27660 28092
rect 27890 28064 27896 28076
rect 27632 28036 27896 28064
rect 27525 28027 27583 28033
rect 27890 28024 27896 28036
rect 27948 28064 27954 28076
rect 28718 28064 28724 28076
rect 27948 28036 28724 28064
rect 27948 28024 27954 28036
rect 28718 28024 28724 28036
rect 28776 28024 28782 28076
rect 28828 28064 28856 28160
rect 29178 28092 29184 28144
rect 29236 28132 29242 28144
rect 29638 28132 29644 28144
rect 29236 28104 29644 28132
rect 29236 28092 29242 28104
rect 29638 28092 29644 28104
rect 29696 28132 29702 28144
rect 29914 28132 29920 28144
rect 29696 28104 29920 28132
rect 29696 28092 29702 28104
rect 29914 28092 29920 28104
rect 29972 28092 29978 28144
rect 31110 28092 31116 28144
rect 31168 28092 31174 28144
rect 29362 28064 29368 28076
rect 28828 28036 29368 28064
rect 29362 28024 29368 28036
rect 29420 28024 29426 28076
rect 30190 28024 30196 28076
rect 30248 28064 30254 28076
rect 30377 28067 30435 28073
rect 30377 28064 30389 28067
rect 30248 28036 30389 28064
rect 30248 28024 30254 28036
rect 30377 28033 30389 28036
rect 30423 28033 30435 28067
rect 30377 28027 30435 28033
rect 24029 27999 24087 28005
rect 24029 27965 24041 27999
rect 24075 27965 24087 27999
rect 24029 27959 24087 27965
rect 24394 27956 24400 28008
rect 24452 27996 24458 28008
rect 24489 27999 24547 28005
rect 24489 27996 24501 27999
rect 24452 27968 24501 27996
rect 24452 27956 24458 27968
rect 24489 27965 24501 27968
rect 24535 27965 24547 27999
rect 24489 27959 24547 27965
rect 24578 27956 24584 28008
rect 24636 27956 24642 28008
rect 25041 27999 25099 28005
rect 25041 27965 25053 27999
rect 25087 27965 25099 27999
rect 25041 27959 25099 27965
rect 13998 27928 14004 27940
rect 13832 27900 14004 27928
rect 13265 27891 13323 27897
rect 13998 27888 14004 27900
rect 14056 27888 14062 27940
rect 16669 27931 16727 27937
rect 16669 27897 16681 27931
rect 16715 27928 16727 27931
rect 16715 27900 17080 27928
rect 16715 27897 16727 27900
rect 16669 27891 16727 27897
rect 11422 27860 11428 27872
rect 11348 27832 11428 27860
rect 11422 27820 11428 27832
rect 11480 27860 11486 27872
rect 13725 27863 13783 27869
rect 13725 27860 13737 27863
rect 11480 27832 13737 27860
rect 11480 27820 11486 27832
rect 13725 27829 13737 27832
rect 13771 27860 13783 27863
rect 16298 27860 16304 27872
rect 13771 27832 16304 27860
rect 13771 27829 13783 27832
rect 13725 27823 13783 27829
rect 16298 27820 16304 27832
rect 16356 27820 16362 27872
rect 17052 27869 17080 27900
rect 17954 27888 17960 27940
rect 18012 27888 18018 27940
rect 19613 27931 19671 27937
rect 19613 27928 19625 27931
rect 19182 27900 19625 27928
rect 19613 27897 19625 27900
rect 19659 27897 19671 27931
rect 25056 27928 25084 27959
rect 25130 27956 25136 28008
rect 25188 27956 25194 28008
rect 25593 27999 25651 28005
rect 25593 27965 25605 27999
rect 25639 27996 25651 27999
rect 26145 27999 26203 28005
rect 26145 27996 26157 27999
rect 25639 27968 26157 27996
rect 25639 27965 25651 27968
rect 25593 27959 25651 27965
rect 26145 27965 26157 27968
rect 26191 27965 26203 27999
rect 26145 27959 26203 27965
rect 26694 27956 26700 28008
rect 26752 27956 26758 28008
rect 26878 27956 26884 28008
rect 26936 27956 26942 28008
rect 27614 27956 27620 28008
rect 27672 27996 27678 28008
rect 28077 27999 28135 28005
rect 28077 27996 28089 27999
rect 27672 27968 28089 27996
rect 27672 27956 27678 27968
rect 28077 27965 28089 27968
rect 28123 27965 28135 27999
rect 28077 27959 28135 27965
rect 28445 27999 28503 28005
rect 28445 27965 28457 27999
rect 28491 27965 28503 27999
rect 28445 27959 28503 27965
rect 28537 27999 28595 28005
rect 28537 27965 28549 27999
rect 28583 27965 28595 27999
rect 28537 27959 28595 27965
rect 19613 27891 19671 27897
rect 24228 27900 25636 27928
rect 17037 27863 17095 27869
rect 17037 27829 17049 27863
rect 17083 27860 17095 27863
rect 17586 27860 17592 27872
rect 17083 27832 17592 27860
rect 17083 27829 17095 27832
rect 17037 27823 17095 27829
rect 17586 27820 17592 27832
rect 17644 27820 17650 27872
rect 22738 27820 22744 27872
rect 22796 27820 22802 27872
rect 24228 27869 24256 27900
rect 25608 27872 25636 27900
rect 26418 27888 26424 27940
rect 26476 27888 26482 27940
rect 27157 27931 27215 27937
rect 27157 27897 27169 27931
rect 27203 27928 27215 27931
rect 27246 27928 27252 27940
rect 27203 27900 27252 27928
rect 27203 27897 27215 27900
rect 27157 27891 27215 27897
rect 27246 27888 27252 27900
rect 27304 27888 27310 27940
rect 27341 27931 27399 27937
rect 27341 27897 27353 27931
rect 27387 27928 27399 27931
rect 27522 27928 27528 27940
rect 27387 27900 27528 27928
rect 27387 27897 27399 27900
rect 27341 27891 27399 27897
rect 27522 27888 27528 27900
rect 27580 27928 27586 27940
rect 28166 27928 28172 27940
rect 27580 27900 28172 27928
rect 27580 27888 27586 27900
rect 28166 27888 28172 27900
rect 28224 27928 28230 27940
rect 28460 27928 28488 27959
rect 28224 27900 28488 27928
rect 28552 27928 28580 27959
rect 28626 27956 28632 28008
rect 28684 27956 28690 28008
rect 29549 27999 29607 28005
rect 29549 27965 29561 27999
rect 29595 27998 29607 27999
rect 29595 27996 29684 27998
rect 30098 27996 30104 28008
rect 29595 27970 30104 27996
rect 29595 27965 29607 27970
rect 29656 27968 30104 27970
rect 28736 27934 28994 27962
rect 29549 27959 29607 27965
rect 30098 27956 30104 27968
rect 30156 27956 30162 28008
rect 31128 27996 31156 28092
rect 31205 27999 31263 28005
rect 31205 27996 31217 27999
rect 31128 27968 31217 27996
rect 31205 27965 31217 27968
rect 31251 27965 31263 27999
rect 31205 27959 31263 27965
rect 28736 27928 28764 27934
rect 28552 27900 28764 27928
rect 28966 27928 28994 27934
rect 29454 27928 29460 27940
rect 28966 27900 29460 27928
rect 28224 27888 28230 27900
rect 24213 27863 24271 27869
rect 24213 27829 24225 27863
rect 24259 27829 24271 27863
rect 24213 27823 24271 27829
rect 24302 27820 24308 27872
rect 24360 27820 24366 27872
rect 25590 27820 25596 27872
rect 25648 27820 25654 27872
rect 25866 27820 25872 27872
rect 25924 27860 25930 27872
rect 26329 27863 26387 27869
rect 26329 27860 26341 27863
rect 25924 27832 26341 27860
rect 25924 27820 25930 27832
rect 26329 27829 26341 27832
rect 26375 27829 26387 27863
rect 26329 27823 26387 27829
rect 26970 27820 26976 27872
rect 27028 27820 27034 27872
rect 27798 27820 27804 27872
rect 27856 27860 27862 27872
rect 28552 27860 28580 27900
rect 29454 27888 29460 27900
rect 29512 27888 29518 27940
rect 30653 27931 30711 27937
rect 30653 27928 30665 27931
rect 29748 27900 30665 27928
rect 27856 27832 28580 27860
rect 27856 27820 27862 27832
rect 28810 27820 28816 27872
rect 28868 27860 28874 27872
rect 28997 27863 29055 27869
rect 28997 27860 29009 27863
rect 28868 27832 29009 27860
rect 28868 27820 28874 27832
rect 28997 27829 29009 27832
rect 29043 27829 29055 27863
rect 28997 27823 29055 27829
rect 29641 27863 29699 27869
rect 29641 27829 29653 27863
rect 29687 27860 29699 27863
rect 29748 27860 29776 27900
rect 30653 27897 30665 27900
rect 30699 27928 30711 27931
rect 30699 27900 31248 27928
rect 30699 27897 30711 27900
rect 30653 27891 30711 27897
rect 31220 27872 31248 27900
rect 29687 27832 29776 27860
rect 29687 27829 29699 27832
rect 29641 27823 29699 27829
rect 29914 27820 29920 27872
rect 29972 27860 29978 27872
rect 30193 27863 30251 27869
rect 30193 27860 30205 27863
rect 29972 27832 30205 27860
rect 29972 27820 29978 27832
rect 30193 27829 30205 27832
rect 30239 27829 30251 27863
rect 30193 27823 30251 27829
rect 30285 27863 30343 27869
rect 30285 27829 30297 27863
rect 30331 27860 30343 27863
rect 30742 27860 30748 27872
rect 30331 27832 30748 27860
rect 30331 27829 30343 27832
rect 30285 27823 30343 27829
rect 30742 27820 30748 27832
rect 30800 27820 30806 27872
rect 30834 27820 30840 27872
rect 30892 27869 30898 27872
rect 30892 27863 30911 27869
rect 30899 27829 30911 27863
rect 30892 27823 30911 27829
rect 30892 27820 30898 27823
rect 31202 27820 31208 27872
rect 31260 27820 31266 27872
rect 31846 27820 31852 27872
rect 31904 27820 31910 27872
rect 2760 27770 32200 27792
rect 2760 27718 6946 27770
rect 6998 27718 7010 27770
rect 7062 27718 7074 27770
rect 7126 27718 7138 27770
rect 7190 27718 7202 27770
rect 7254 27718 14306 27770
rect 14358 27718 14370 27770
rect 14422 27718 14434 27770
rect 14486 27718 14498 27770
rect 14550 27718 14562 27770
rect 14614 27718 21666 27770
rect 21718 27718 21730 27770
rect 21782 27718 21794 27770
rect 21846 27718 21858 27770
rect 21910 27718 21922 27770
rect 21974 27718 29026 27770
rect 29078 27718 29090 27770
rect 29142 27718 29154 27770
rect 29206 27718 29218 27770
rect 29270 27718 29282 27770
rect 29334 27718 32200 27770
rect 2760 27696 32200 27718
rect 5258 27616 5264 27668
rect 5316 27616 5322 27668
rect 6457 27659 6515 27665
rect 6457 27625 6469 27659
rect 6503 27656 6515 27659
rect 6638 27656 6644 27668
rect 6503 27628 6644 27656
rect 6503 27625 6515 27628
rect 6457 27619 6515 27625
rect 6638 27616 6644 27628
rect 6696 27616 6702 27668
rect 7282 27656 7288 27668
rect 7116 27628 7288 27656
rect 5077 27591 5135 27597
rect 5077 27557 5089 27591
rect 5123 27588 5135 27591
rect 5276 27588 5304 27616
rect 5123 27560 5304 27588
rect 5123 27557 5135 27560
rect 5077 27551 5135 27557
rect 6546 27548 6552 27600
rect 6604 27588 6610 27600
rect 6733 27591 6791 27597
rect 6733 27588 6745 27591
rect 6604 27560 6745 27588
rect 6604 27548 6610 27560
rect 6733 27557 6745 27560
rect 6779 27588 6791 27591
rect 6914 27588 6920 27600
rect 6779 27560 6920 27588
rect 6779 27557 6791 27560
rect 6733 27551 6791 27557
rect 6914 27548 6920 27560
rect 6972 27548 6978 27600
rect 4433 27523 4491 27529
rect 4433 27489 4445 27523
rect 4479 27489 4491 27523
rect 4433 27483 4491 27489
rect 5169 27523 5227 27529
rect 5169 27489 5181 27523
rect 5215 27520 5227 27523
rect 6178 27520 6184 27532
rect 5215 27492 6184 27520
rect 5215 27489 5227 27492
rect 5169 27483 5227 27489
rect 1302 27412 1308 27464
rect 1360 27452 1366 27464
rect 3237 27455 3295 27461
rect 3237 27452 3249 27455
rect 1360 27424 3249 27452
rect 1360 27412 1366 27424
rect 3237 27421 3249 27424
rect 3283 27421 3295 27455
rect 4448 27452 4476 27483
rect 6178 27480 6184 27492
rect 6236 27480 6242 27532
rect 6641 27523 6699 27529
rect 6641 27520 6653 27523
rect 6564 27492 6653 27520
rect 4448 27424 5672 27452
rect 3237 27415 3295 27421
rect 5534 27276 5540 27328
rect 5592 27276 5598 27328
rect 5644 27316 5672 27424
rect 6564 27384 6592 27492
rect 6641 27489 6653 27492
rect 6687 27489 6699 27523
rect 6641 27483 6699 27489
rect 6822 27480 6828 27532
rect 6880 27480 6886 27532
rect 7009 27523 7067 27529
rect 7009 27489 7021 27523
rect 7055 27520 7067 27523
rect 7116 27520 7144 27628
rect 7282 27616 7288 27628
rect 7340 27656 7346 27668
rect 8938 27656 8944 27668
rect 7340 27628 8944 27656
rect 7340 27616 7346 27628
rect 8938 27616 8944 27628
rect 8996 27616 9002 27668
rect 10318 27616 10324 27668
rect 10376 27656 10382 27668
rect 10376 27628 10732 27656
rect 10376 27616 10382 27628
rect 7190 27548 7196 27600
rect 7248 27588 7254 27600
rect 8849 27591 8907 27597
rect 8849 27588 8861 27591
rect 7248 27560 8861 27588
rect 7248 27548 7254 27560
rect 8849 27557 8861 27560
rect 8895 27557 8907 27591
rect 8849 27551 8907 27557
rect 9674 27548 9680 27600
rect 9732 27588 9738 27600
rect 10704 27588 10732 27628
rect 11606 27616 11612 27668
rect 11664 27656 11670 27668
rect 11885 27659 11943 27665
rect 11885 27656 11897 27659
rect 11664 27628 11897 27656
rect 11664 27616 11670 27628
rect 11885 27625 11897 27628
rect 11931 27625 11943 27659
rect 11885 27619 11943 27625
rect 13998 27616 14004 27668
rect 14056 27656 14062 27668
rect 14734 27656 14740 27668
rect 14056 27628 14740 27656
rect 14056 27616 14062 27628
rect 14734 27616 14740 27628
rect 14792 27616 14798 27668
rect 17865 27659 17923 27665
rect 17865 27625 17877 27659
rect 17911 27656 17923 27659
rect 17954 27656 17960 27668
rect 17911 27628 17960 27656
rect 17911 27625 17923 27628
rect 17865 27619 17923 27625
rect 17954 27616 17960 27628
rect 18012 27616 18018 27668
rect 23934 27656 23940 27668
rect 22940 27628 23940 27656
rect 9732 27560 10088 27588
rect 10704 27560 10810 27588
rect 9732 27548 9738 27560
rect 7055 27492 7144 27520
rect 7055 27489 7067 27492
rect 7009 27483 7067 27489
rect 9030 27480 9036 27532
rect 9088 27520 9094 27532
rect 10060 27529 10088 27560
rect 12434 27548 12440 27600
rect 12492 27548 12498 27600
rect 13446 27548 13452 27600
rect 13504 27588 13510 27600
rect 13909 27591 13967 27597
rect 13909 27588 13921 27591
rect 13504 27560 13921 27588
rect 13504 27548 13510 27560
rect 13909 27557 13921 27560
rect 13955 27588 13967 27591
rect 14645 27591 14703 27597
rect 14645 27588 14657 27591
rect 13955 27560 14657 27588
rect 13955 27557 13967 27560
rect 13909 27551 13967 27557
rect 14645 27557 14657 27560
rect 14691 27588 14703 27591
rect 14918 27588 14924 27600
rect 14691 27560 14924 27588
rect 14691 27557 14703 27560
rect 14645 27551 14703 27557
rect 14918 27548 14924 27560
rect 14976 27548 14982 27600
rect 16022 27548 16028 27600
rect 16080 27548 16086 27600
rect 17589 27591 17647 27597
rect 17589 27557 17601 27591
rect 17635 27588 17647 27591
rect 20438 27588 20444 27600
rect 17635 27560 20444 27588
rect 17635 27557 17647 27560
rect 17589 27551 17647 27557
rect 20438 27548 20444 27560
rect 20496 27548 20502 27600
rect 22940 27588 22968 27628
rect 23934 27616 23940 27628
rect 23992 27656 23998 27668
rect 23992 27628 24348 27656
rect 23992 27616 23998 27628
rect 24320 27600 24348 27628
rect 24394 27616 24400 27668
rect 24452 27656 24458 27668
rect 24762 27656 24768 27668
rect 24452 27628 24768 27656
rect 24452 27616 24458 27628
rect 24762 27616 24768 27628
rect 24820 27656 24826 27668
rect 25317 27659 25375 27665
rect 25317 27656 25329 27659
rect 24820 27628 25329 27656
rect 24820 27616 24826 27628
rect 25317 27625 25329 27628
rect 25363 27656 25375 27659
rect 25682 27656 25688 27668
rect 25363 27628 25688 27656
rect 25363 27625 25375 27628
rect 25317 27619 25375 27625
rect 25682 27616 25688 27628
rect 25740 27656 25746 27668
rect 26878 27656 26884 27668
rect 25740 27628 26884 27656
rect 25740 27616 25746 27628
rect 26878 27616 26884 27628
rect 26936 27616 26942 27668
rect 28166 27616 28172 27668
rect 28224 27656 28230 27668
rect 30374 27656 30380 27668
rect 28224 27628 30380 27656
rect 28224 27616 28230 27628
rect 30374 27616 30380 27628
rect 30432 27616 30438 27668
rect 30742 27616 30748 27668
rect 30800 27616 30806 27668
rect 30908 27659 30966 27665
rect 30908 27656 30920 27659
rect 30852 27628 30920 27656
rect 21744 27560 22968 27588
rect 23017 27591 23075 27597
rect 9401 27523 9459 27529
rect 9401 27520 9413 27523
rect 9088 27492 9413 27520
rect 9088 27480 9094 27492
rect 9401 27489 9413 27492
rect 9447 27489 9459 27523
rect 9401 27483 9459 27489
rect 9769 27523 9827 27529
rect 9769 27489 9781 27523
rect 9815 27489 9827 27523
rect 9769 27483 9827 27489
rect 10045 27523 10103 27529
rect 10045 27489 10057 27523
rect 10091 27489 10103 27523
rect 10045 27483 10103 27489
rect 7101 27455 7159 27461
rect 7101 27421 7113 27455
rect 7147 27421 7159 27455
rect 7101 27415 7159 27421
rect 6564 27356 6776 27384
rect 6638 27316 6644 27328
rect 5644 27288 6644 27316
rect 6638 27276 6644 27288
rect 6696 27276 6702 27328
rect 6748 27316 6776 27356
rect 6822 27344 6828 27396
rect 6880 27384 6886 27396
rect 7116 27384 7144 27415
rect 8110 27412 8116 27464
rect 8168 27412 8174 27464
rect 9784 27452 9812 27483
rect 12158 27480 12164 27532
rect 12216 27480 12222 27532
rect 14277 27523 14335 27529
rect 14277 27489 14289 27523
rect 14323 27520 14335 27523
rect 14458 27520 14464 27532
rect 14323 27492 14464 27520
rect 14323 27489 14335 27492
rect 14277 27483 14335 27489
rect 14458 27480 14464 27492
rect 14516 27480 14522 27532
rect 16298 27480 16304 27532
rect 16356 27520 16362 27532
rect 16758 27520 16764 27532
rect 16356 27492 16764 27520
rect 16356 27480 16362 27492
rect 16758 27480 16764 27492
rect 16816 27520 16822 27532
rect 17313 27523 17371 27529
rect 17313 27520 17325 27523
rect 16816 27492 17325 27520
rect 16816 27480 16822 27492
rect 17313 27489 17325 27492
rect 17359 27489 17371 27523
rect 17313 27483 17371 27489
rect 9784 27424 10088 27452
rect 6880 27356 7144 27384
rect 9677 27387 9735 27393
rect 6880 27344 6886 27356
rect 9677 27353 9689 27387
rect 9723 27384 9735 27387
rect 9766 27384 9772 27396
rect 9723 27356 9772 27384
rect 9723 27353 9735 27356
rect 9677 27347 9735 27353
rect 9766 27344 9772 27356
rect 9824 27344 9830 27396
rect 10060 27328 10088 27424
rect 10318 27412 10324 27464
rect 10376 27412 10382 27464
rect 12069 27455 12127 27461
rect 12069 27421 12081 27455
rect 12115 27421 12127 27455
rect 12069 27415 12127 27421
rect 11790 27344 11796 27396
rect 11848 27344 11854 27396
rect 12084 27384 12112 27415
rect 12526 27412 12532 27464
rect 12584 27412 12590 27464
rect 12897 27455 12955 27461
rect 12897 27421 12909 27455
rect 12943 27452 12955 27455
rect 13541 27455 13599 27461
rect 13541 27452 13553 27455
rect 12943 27424 13553 27452
rect 12943 27421 12955 27424
rect 12897 27415 12955 27421
rect 13541 27421 13553 27424
rect 13587 27452 13599 27455
rect 14185 27455 14243 27461
rect 14185 27452 14197 27455
rect 13587 27424 14197 27452
rect 13587 27421 13599 27424
rect 13541 27415 13599 27421
rect 14185 27421 14197 27424
rect 14231 27452 14243 27455
rect 14366 27452 14372 27464
rect 14231 27424 14372 27452
rect 14231 27421 14243 27424
rect 14185 27415 14243 27421
rect 12342 27384 12348 27396
rect 12084 27356 12348 27384
rect 12342 27344 12348 27356
rect 12400 27384 12406 27396
rect 12912 27384 12940 27415
rect 14366 27412 14372 27424
rect 14424 27412 14430 27464
rect 14553 27455 14611 27461
rect 14553 27421 14565 27455
rect 14599 27421 14611 27455
rect 14553 27415 14611 27421
rect 12400 27356 12940 27384
rect 12400 27344 12406 27356
rect 7650 27316 7656 27328
rect 6748 27288 7656 27316
rect 7650 27276 7656 27288
rect 7708 27276 7714 27328
rect 7745 27319 7803 27325
rect 7745 27285 7757 27319
rect 7791 27316 7803 27319
rect 8386 27316 8392 27328
rect 7791 27288 8392 27316
rect 7791 27285 7803 27288
rect 7745 27279 7803 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8754 27276 8760 27328
rect 8812 27276 8818 27328
rect 10042 27276 10048 27328
rect 10100 27276 10106 27328
rect 14001 27319 14059 27325
rect 14001 27285 14013 27319
rect 14047 27316 14059 27319
rect 14182 27316 14188 27328
rect 14047 27288 14188 27316
rect 14047 27285 14059 27288
rect 14001 27279 14059 27285
rect 14182 27276 14188 27288
rect 14240 27276 14246 27328
rect 14568 27316 14596 27415
rect 14734 27412 14740 27464
rect 14792 27412 14798 27464
rect 15010 27412 15016 27464
rect 15068 27412 15074 27464
rect 16485 27455 16543 27461
rect 16485 27421 16497 27455
rect 16531 27452 16543 27455
rect 17126 27452 17132 27464
rect 16531 27424 17132 27452
rect 16531 27421 16543 27424
rect 16485 27415 16543 27421
rect 17126 27412 17132 27424
rect 17184 27412 17190 27464
rect 17328 27452 17356 27483
rect 17494 27480 17500 27532
rect 17552 27480 17558 27532
rect 17678 27480 17684 27532
rect 17736 27480 17742 27532
rect 18966 27480 18972 27532
rect 19024 27520 19030 27532
rect 19153 27523 19211 27529
rect 19153 27520 19165 27523
rect 19024 27492 19165 27520
rect 19024 27480 19030 27492
rect 19153 27489 19165 27492
rect 19199 27520 19211 27523
rect 19702 27520 19708 27532
rect 19199 27492 19708 27520
rect 19199 27489 19211 27492
rect 19153 27483 19211 27489
rect 19702 27480 19708 27492
rect 19760 27480 19766 27532
rect 21744 27529 21772 27560
rect 23017 27557 23029 27591
rect 23063 27588 23075 27591
rect 23566 27588 23572 27600
rect 23063 27560 23572 27588
rect 23063 27557 23075 27560
rect 23017 27551 23075 27557
rect 23566 27548 23572 27560
rect 23624 27588 23630 27600
rect 24026 27588 24032 27600
rect 23624 27560 24032 27588
rect 23624 27548 23630 27560
rect 24026 27548 24032 27560
rect 24084 27548 24090 27600
rect 24302 27548 24308 27600
rect 24360 27548 24366 27600
rect 25593 27591 25651 27597
rect 25593 27557 25605 27591
rect 25639 27588 25651 27591
rect 26418 27588 26424 27600
rect 25639 27560 26424 27588
rect 25639 27557 25651 27560
rect 25593 27551 25651 27557
rect 26418 27548 26424 27560
rect 26476 27548 26482 27600
rect 27338 27548 27344 27600
rect 27396 27588 27402 27600
rect 30558 27588 30564 27600
rect 27396 27560 27752 27588
rect 27396 27548 27402 27560
rect 21729 27523 21787 27529
rect 21729 27489 21741 27523
rect 21775 27489 21787 27523
rect 21729 27483 21787 27489
rect 21913 27523 21971 27529
rect 21913 27489 21925 27523
rect 21959 27489 21971 27523
rect 21913 27483 21971 27489
rect 18509 27455 18567 27461
rect 18509 27452 18521 27455
rect 17328 27424 18521 27452
rect 18509 27421 18521 27424
rect 18555 27421 18567 27455
rect 18509 27415 18567 27421
rect 19242 27412 19248 27464
rect 19300 27412 19306 27464
rect 19794 27412 19800 27464
rect 19852 27452 19858 27464
rect 20533 27455 20591 27461
rect 20533 27452 20545 27455
rect 19852 27424 20545 27452
rect 19852 27412 19858 27424
rect 20533 27421 20545 27424
rect 20579 27421 20591 27455
rect 21928 27452 21956 27483
rect 22002 27480 22008 27532
rect 22060 27480 22066 27532
rect 23201 27523 23259 27529
rect 23201 27489 23213 27523
rect 23247 27489 23259 27523
rect 23201 27483 23259 27489
rect 23293 27523 23351 27529
rect 23293 27489 23305 27523
rect 23339 27489 23351 27523
rect 23293 27483 23351 27489
rect 22738 27452 22744 27464
rect 21928 27424 22744 27452
rect 20533 27415 20591 27421
rect 22738 27412 22744 27424
rect 22796 27412 22802 27464
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27421 22891 27455
rect 22833 27415 22891 27421
rect 21913 27387 21971 27393
rect 21913 27353 21925 27387
rect 21959 27384 21971 27387
rect 22848 27384 22876 27415
rect 23106 27412 23112 27464
rect 23164 27412 23170 27464
rect 21959 27356 22876 27384
rect 23017 27387 23075 27393
rect 21959 27353 21971 27356
rect 21913 27347 21971 27353
rect 23017 27353 23029 27387
rect 23063 27384 23075 27387
rect 23124 27384 23152 27412
rect 23063 27356 23152 27384
rect 23063 27353 23075 27356
rect 23017 27347 23075 27353
rect 16850 27316 16856 27328
rect 14568 27288 16856 27316
rect 16850 27276 16856 27288
rect 16908 27276 16914 27328
rect 17126 27276 17132 27328
rect 17184 27316 17190 27328
rect 17678 27316 17684 27328
rect 17184 27288 17684 27316
rect 17184 27276 17190 27288
rect 17678 27276 17684 27288
rect 17736 27276 17742 27328
rect 19058 27276 19064 27328
rect 19116 27276 19122 27328
rect 19150 27276 19156 27328
rect 19208 27316 19214 27328
rect 19889 27319 19947 27325
rect 19889 27316 19901 27319
rect 19208 27288 19901 27316
rect 19208 27276 19214 27288
rect 19889 27285 19901 27288
rect 19935 27285 19947 27319
rect 19889 27279 19947 27285
rect 19978 27276 19984 27328
rect 20036 27276 20042 27328
rect 22094 27276 22100 27328
rect 22152 27276 22158 27328
rect 22186 27276 22192 27328
rect 22244 27316 22250 27328
rect 22281 27319 22339 27325
rect 22281 27316 22293 27319
rect 22244 27288 22293 27316
rect 22244 27276 22250 27288
rect 22281 27285 22293 27288
rect 22327 27285 22339 27319
rect 22281 27279 22339 27285
rect 23106 27276 23112 27328
rect 23164 27316 23170 27328
rect 23216 27316 23244 27483
rect 23308 27452 23336 27483
rect 23382 27480 23388 27532
rect 23440 27520 23446 27532
rect 23477 27523 23535 27529
rect 23477 27520 23489 27523
rect 23440 27492 23489 27520
rect 23440 27480 23446 27492
rect 23477 27489 23489 27492
rect 23523 27520 23535 27523
rect 25133 27523 25191 27529
rect 25133 27520 25145 27523
rect 23523 27492 25145 27520
rect 23523 27489 23535 27492
rect 23477 27483 23535 27489
rect 25133 27489 25145 27492
rect 25179 27489 25191 27523
rect 25133 27483 25191 27489
rect 25225 27523 25283 27529
rect 25225 27489 25237 27523
rect 25271 27489 25283 27523
rect 25225 27483 25283 27489
rect 25869 27523 25927 27529
rect 25869 27489 25881 27523
rect 25915 27520 25927 27523
rect 26050 27520 26056 27532
rect 25915 27492 26056 27520
rect 25915 27489 25927 27492
rect 25869 27483 25927 27489
rect 23308 27424 23612 27452
rect 23584 27328 23612 27424
rect 23658 27412 23664 27464
rect 23716 27452 23722 27464
rect 24578 27452 24584 27464
rect 23716 27424 24584 27452
rect 23716 27412 23722 27424
rect 24578 27412 24584 27424
rect 24636 27452 24642 27464
rect 24857 27455 24915 27461
rect 24857 27452 24869 27455
rect 24636 27424 24869 27452
rect 24636 27412 24642 27424
rect 24857 27421 24869 27424
rect 24903 27452 24915 27455
rect 25240 27452 25268 27483
rect 26050 27480 26056 27492
rect 26108 27480 26114 27532
rect 27614 27520 27620 27532
rect 26804 27492 27620 27520
rect 24903 27424 25268 27452
rect 25777 27455 25835 27461
rect 24903 27421 24915 27424
rect 24857 27415 24915 27421
rect 25777 27421 25789 27455
rect 25823 27452 25835 27455
rect 26804 27452 26832 27492
rect 27614 27480 27620 27492
rect 27672 27480 27678 27532
rect 27724 27529 27752 27560
rect 28092 27560 30564 27588
rect 28092 27529 28120 27560
rect 30558 27548 30564 27560
rect 30616 27548 30622 27600
rect 30852 27532 30880 27628
rect 30908 27625 30920 27628
rect 30954 27625 30966 27659
rect 30908 27619 30966 27625
rect 31110 27548 31116 27600
rect 31168 27588 31174 27600
rect 31846 27588 31852 27600
rect 31168 27560 31852 27588
rect 31168 27548 31174 27560
rect 31846 27548 31852 27560
rect 31904 27548 31910 27600
rect 27709 27523 27767 27529
rect 27709 27489 27721 27523
rect 27755 27520 27767 27523
rect 28077 27523 28135 27529
rect 28077 27520 28089 27523
rect 27755 27492 28089 27520
rect 27755 27489 27767 27492
rect 27709 27483 27767 27489
rect 28077 27489 28089 27492
rect 28123 27489 28135 27523
rect 28077 27483 28135 27489
rect 28166 27480 28172 27532
rect 28224 27520 28230 27532
rect 28261 27523 28319 27529
rect 28261 27520 28273 27523
rect 28224 27492 28273 27520
rect 28224 27480 28230 27492
rect 28261 27489 28273 27492
rect 28307 27489 28319 27523
rect 28261 27483 28319 27489
rect 28534 27480 28540 27532
rect 28592 27520 28598 27532
rect 28813 27523 28871 27529
rect 28813 27520 28825 27523
rect 28592 27492 28825 27520
rect 28592 27480 28598 27492
rect 28813 27489 28825 27492
rect 28859 27520 28871 27523
rect 28994 27520 29000 27532
rect 28859 27492 29000 27520
rect 28859 27489 28871 27492
rect 28813 27483 28871 27489
rect 28994 27480 29000 27492
rect 29052 27480 29058 27532
rect 29273 27523 29331 27529
rect 29273 27489 29285 27523
rect 29319 27520 29331 27523
rect 29546 27520 29552 27532
rect 29319 27492 29552 27520
rect 29319 27489 29331 27492
rect 29273 27483 29331 27489
rect 29546 27480 29552 27492
rect 29604 27480 29610 27532
rect 29730 27480 29736 27532
rect 29788 27480 29794 27532
rect 30834 27480 30840 27532
rect 30892 27480 30898 27532
rect 31205 27523 31263 27529
rect 31205 27489 31217 27523
rect 31251 27520 31263 27523
rect 31294 27520 31300 27532
rect 31251 27492 31300 27520
rect 31251 27489 31263 27492
rect 31205 27483 31263 27489
rect 31294 27480 31300 27492
rect 31352 27480 31358 27532
rect 25823 27424 26832 27452
rect 25823 27421 25835 27424
rect 25777 27415 25835 27421
rect 26878 27412 26884 27464
rect 26936 27412 26942 27464
rect 24026 27344 24032 27396
rect 24084 27384 24090 27396
rect 24121 27387 24179 27393
rect 24121 27384 24133 27387
rect 24084 27356 24133 27384
rect 24084 27344 24090 27356
rect 24121 27353 24133 27356
rect 24167 27384 24179 27387
rect 24167 27356 24532 27384
rect 24167 27353 24179 27356
rect 24121 27347 24179 27353
rect 24504 27328 24532 27356
rect 24946 27344 24952 27396
rect 25004 27344 25010 27396
rect 26786 27384 26792 27396
rect 25424 27356 26792 27384
rect 23164 27288 23244 27316
rect 23164 27276 23170 27288
rect 23566 27276 23572 27328
rect 23624 27276 23630 27328
rect 24210 27276 24216 27328
rect 24268 27276 24274 27328
rect 24486 27276 24492 27328
rect 24544 27276 24550 27328
rect 24578 27276 24584 27328
rect 24636 27316 24642 27328
rect 25424 27316 25452 27356
rect 26786 27344 26792 27356
rect 26844 27384 26850 27396
rect 27430 27384 27436 27396
rect 26844 27356 27436 27384
rect 26844 27344 26850 27356
rect 27430 27344 27436 27356
rect 27488 27344 27494 27396
rect 27632 27384 27660 27480
rect 27982 27412 27988 27464
rect 28040 27452 28046 27464
rect 28626 27452 28632 27464
rect 28040 27424 28632 27452
rect 28040 27412 28046 27424
rect 28626 27412 28632 27424
rect 28684 27412 28690 27464
rect 29457 27455 29515 27461
rect 29457 27421 29469 27455
rect 29503 27452 29515 27455
rect 29503 27424 30052 27452
rect 29503 27421 29515 27424
rect 29457 27415 29515 27421
rect 29089 27387 29147 27393
rect 29089 27384 29101 27387
rect 27632 27356 29101 27384
rect 29089 27353 29101 27356
rect 29135 27353 29147 27387
rect 29089 27347 29147 27353
rect 29546 27344 29552 27396
rect 29604 27344 29610 27396
rect 24636 27288 25452 27316
rect 24636 27276 24642 27288
rect 25498 27276 25504 27328
rect 25556 27276 25562 27328
rect 25590 27276 25596 27328
rect 25648 27276 25654 27328
rect 26050 27276 26056 27328
rect 26108 27276 26114 27328
rect 26326 27276 26332 27328
rect 26384 27276 26390 27328
rect 26602 27276 26608 27328
rect 26660 27316 26666 27328
rect 28169 27319 28227 27325
rect 28169 27316 28181 27319
rect 26660 27288 28181 27316
rect 26660 27276 26666 27288
rect 28169 27285 28181 27288
rect 28215 27285 28227 27319
rect 28169 27279 28227 27285
rect 28721 27319 28779 27325
rect 28721 27285 28733 27319
rect 28767 27316 28779 27319
rect 28902 27316 28908 27328
rect 28767 27288 28908 27316
rect 28767 27285 28779 27288
rect 28721 27279 28779 27285
rect 28902 27276 28908 27288
rect 28960 27276 28966 27328
rect 29564 27316 29592 27344
rect 30024 27325 30052 27424
rect 30374 27412 30380 27464
rect 30432 27412 30438 27464
rect 30650 27412 30656 27464
rect 30708 27412 30714 27464
rect 30926 27412 30932 27464
rect 30984 27452 30990 27464
rect 31389 27455 31447 27461
rect 31389 27452 31401 27455
rect 30984 27424 31401 27452
rect 30984 27412 30990 27424
rect 31389 27421 31401 27424
rect 31435 27421 31447 27455
rect 31389 27415 31447 27421
rect 30392 27384 30420 27412
rect 30392 27356 30972 27384
rect 29641 27319 29699 27325
rect 29641 27316 29653 27319
rect 29564 27288 29653 27316
rect 29641 27285 29653 27288
rect 29687 27285 29699 27319
rect 29641 27279 29699 27285
rect 30009 27319 30067 27325
rect 30009 27285 30021 27319
rect 30055 27316 30067 27319
rect 30466 27316 30472 27328
rect 30055 27288 30472 27316
rect 30055 27285 30067 27288
rect 30009 27279 30067 27285
rect 30466 27276 30472 27288
rect 30524 27276 30530 27328
rect 30944 27325 30972 27356
rect 30929 27319 30987 27325
rect 30929 27285 30941 27319
rect 30975 27285 30987 27319
rect 30929 27279 30987 27285
rect 2760 27226 32200 27248
rect 2760 27174 6286 27226
rect 6338 27174 6350 27226
rect 6402 27174 6414 27226
rect 6466 27174 6478 27226
rect 6530 27174 6542 27226
rect 6594 27174 13646 27226
rect 13698 27174 13710 27226
rect 13762 27174 13774 27226
rect 13826 27174 13838 27226
rect 13890 27174 13902 27226
rect 13954 27174 21006 27226
rect 21058 27174 21070 27226
rect 21122 27174 21134 27226
rect 21186 27174 21198 27226
rect 21250 27174 21262 27226
rect 21314 27174 28366 27226
rect 28418 27174 28430 27226
rect 28482 27174 28494 27226
rect 28546 27174 28558 27226
rect 28610 27174 28622 27226
rect 28674 27174 32200 27226
rect 2760 27152 32200 27174
rect 7009 27115 7067 27121
rect 7009 27081 7021 27115
rect 7055 27112 7067 27115
rect 8110 27112 8116 27124
rect 7055 27084 8116 27112
rect 7055 27081 7067 27084
rect 7009 27075 7067 27081
rect 8110 27072 8116 27084
rect 8168 27072 8174 27124
rect 9585 27115 9643 27121
rect 9585 27081 9597 27115
rect 9631 27112 9643 27115
rect 9858 27112 9864 27124
rect 9631 27084 9864 27112
rect 9631 27081 9643 27084
rect 9585 27075 9643 27081
rect 9858 27072 9864 27084
rect 9916 27072 9922 27124
rect 10318 27072 10324 27124
rect 10376 27112 10382 27124
rect 10689 27115 10747 27121
rect 10689 27112 10701 27115
rect 10376 27084 10701 27112
rect 10376 27072 10382 27084
rect 10689 27081 10701 27084
rect 10735 27081 10747 27115
rect 10689 27075 10747 27081
rect 11146 27072 11152 27124
rect 11204 27112 11210 27124
rect 11422 27112 11428 27124
rect 11204 27084 11428 27112
rect 11204 27072 11210 27084
rect 11422 27072 11428 27084
rect 11480 27072 11486 27124
rect 14921 27115 14979 27121
rect 14921 27081 14933 27115
rect 14967 27112 14979 27115
rect 15010 27112 15016 27124
rect 14967 27084 15016 27112
rect 14967 27081 14979 27084
rect 14921 27075 14979 27081
rect 15010 27072 15016 27084
rect 15068 27072 15074 27124
rect 17494 27112 17500 27124
rect 16546 27084 17500 27112
rect 8849 27047 8907 27053
rect 8849 27044 8861 27047
rect 8680 27016 8861 27044
rect 8481 26979 8539 26985
rect 8481 26945 8493 26979
rect 8527 26976 8539 26979
rect 8680 26976 8708 27016
rect 8849 27013 8861 27016
rect 8895 27013 8907 27047
rect 8849 27007 8907 27013
rect 8938 27004 8944 27056
rect 8996 27044 9002 27056
rect 8996 27016 10180 27044
rect 8996 27004 9002 27016
rect 8527 26948 8708 26976
rect 8527 26945 8539 26948
rect 8481 26939 8539 26945
rect 9950 26936 9956 26988
rect 10008 26936 10014 26988
rect 6178 26868 6184 26920
rect 6236 26908 6242 26920
rect 6825 26911 6883 26917
rect 6825 26908 6837 26911
rect 6236 26880 6837 26908
rect 6236 26868 6242 26880
rect 6825 26877 6837 26880
rect 6871 26877 6883 26911
rect 6825 26871 6883 26877
rect 8757 26911 8815 26917
rect 8757 26877 8769 26911
rect 8803 26877 8815 26911
rect 8757 26871 8815 26877
rect 6638 26732 6644 26784
rect 6696 26772 6702 26784
rect 6733 26775 6791 26781
rect 6733 26772 6745 26775
rect 6696 26744 6745 26772
rect 6696 26732 6702 26744
rect 6733 26741 6745 26744
rect 6779 26741 6791 26775
rect 6840 26772 6868 26871
rect 7742 26800 7748 26852
rect 7800 26800 7806 26852
rect 8478 26800 8484 26852
rect 8536 26840 8542 26852
rect 8772 26840 8800 26871
rect 9398 26868 9404 26920
rect 9456 26868 9462 26920
rect 9674 26868 9680 26920
rect 9732 26908 9738 26920
rect 9769 26911 9827 26917
rect 9769 26908 9781 26911
rect 9732 26880 9781 26908
rect 9732 26868 9738 26880
rect 9769 26877 9781 26880
rect 9815 26877 9827 26911
rect 9769 26871 9827 26877
rect 9861 26911 9919 26917
rect 9861 26877 9873 26911
rect 9907 26908 9919 26911
rect 9968 26908 9996 26936
rect 10152 26917 10180 27016
rect 10594 27004 10600 27056
rect 10652 27044 10658 27056
rect 14645 27047 14703 27053
rect 10652 27016 11376 27044
rect 10652 27004 10658 27016
rect 10873 26979 10931 26985
rect 10873 26945 10885 26979
rect 10919 26976 10931 26979
rect 10919 26948 11192 26976
rect 10919 26945 10931 26948
rect 10873 26939 10931 26945
rect 9907 26880 9996 26908
rect 10137 26911 10195 26917
rect 9907 26877 9919 26880
rect 9861 26871 9919 26877
rect 10137 26877 10149 26911
rect 10183 26877 10195 26911
rect 10137 26871 10195 26877
rect 9582 26840 9588 26852
rect 8536 26812 9588 26840
rect 8536 26800 8542 26812
rect 9582 26800 9588 26812
rect 9640 26800 9646 26852
rect 9953 26843 10011 26849
rect 9953 26840 9965 26843
rect 9876 26812 9965 26840
rect 9876 26784 9904 26812
rect 9953 26809 9965 26812
rect 9999 26809 10011 26843
rect 10152 26840 10180 26871
rect 10962 26868 10968 26920
rect 11020 26868 11026 26920
rect 11164 26908 11192 26948
rect 11238 26936 11244 26988
rect 11296 26936 11302 26988
rect 11348 26985 11376 27016
rect 14645 27013 14657 27047
rect 14691 27044 14703 27047
rect 16546 27044 16574 27084
rect 17494 27072 17500 27084
rect 17552 27072 17558 27124
rect 19978 27072 19984 27124
rect 20036 27072 20042 27124
rect 23106 27072 23112 27124
rect 23164 27112 23170 27124
rect 23658 27112 23664 27124
rect 23164 27084 23664 27112
rect 23164 27072 23170 27084
rect 23658 27072 23664 27084
rect 23716 27072 23722 27124
rect 24210 27072 24216 27124
rect 24268 27072 24274 27124
rect 26326 27121 26332 27124
rect 26316 27115 26332 27121
rect 26316 27081 26328 27115
rect 26316 27075 26332 27081
rect 26326 27072 26332 27075
rect 26384 27072 26390 27124
rect 27801 27115 27859 27121
rect 27801 27081 27813 27115
rect 27847 27112 27859 27115
rect 27982 27112 27988 27124
rect 27847 27084 27988 27112
rect 27847 27081 27859 27084
rect 27801 27075 27859 27081
rect 27982 27072 27988 27084
rect 28040 27072 28046 27124
rect 29822 27112 29828 27124
rect 28092 27084 29828 27112
rect 14691 27016 16574 27044
rect 14691 27013 14703 27016
rect 14645 27007 14703 27013
rect 11333 26979 11391 26985
rect 11333 26945 11345 26979
rect 11379 26976 11391 26979
rect 11701 26979 11759 26985
rect 11701 26976 11713 26979
rect 11379 26948 11713 26976
rect 11379 26945 11391 26948
rect 11333 26939 11391 26945
rect 11701 26945 11713 26948
rect 11747 26976 11759 26979
rect 11747 26948 12480 26976
rect 11747 26945 11759 26948
rect 11701 26939 11759 26945
rect 11164 26880 12112 26908
rect 11146 26840 11152 26852
rect 10152 26812 11152 26840
rect 9953 26803 10011 26809
rect 11146 26800 11152 26812
rect 11204 26800 11210 26852
rect 12084 26849 12112 26880
rect 12452 26852 12480 26948
rect 14366 26936 14372 26988
rect 14424 26976 14430 26988
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 14424 26948 15117 26976
rect 14424 26936 14430 26948
rect 15105 26945 15117 26948
rect 15151 26976 15163 26979
rect 15473 26979 15531 26985
rect 15151 26948 15332 26976
rect 15151 26945 15163 26948
rect 15105 26939 15163 26945
rect 14090 26868 14096 26920
rect 14148 26868 14154 26920
rect 14918 26868 14924 26920
rect 14976 26868 14982 26920
rect 15194 26868 15200 26920
rect 15252 26868 15258 26920
rect 15304 26908 15332 26948
rect 15473 26945 15485 26979
rect 15519 26976 15531 26979
rect 17770 26976 17776 26988
rect 15519 26948 17776 26976
rect 15519 26945 15531 26948
rect 15473 26939 15531 26945
rect 17770 26936 17776 26948
rect 17828 26936 17834 26988
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26976 19855 26979
rect 19996 26976 20024 27072
rect 23201 27047 23259 27053
rect 23201 27013 23213 27047
rect 23247 27013 23259 27047
rect 23201 27007 23259 27013
rect 19843 26948 20024 26976
rect 20073 26979 20131 26985
rect 19843 26945 19855 26948
rect 19797 26939 19855 26945
rect 20073 26945 20085 26979
rect 20119 26976 20131 26979
rect 20530 26976 20536 26988
rect 20119 26948 20536 26976
rect 20119 26945 20131 26948
rect 20073 26939 20131 26945
rect 20530 26936 20536 26948
rect 20588 26976 20594 26988
rect 21358 26976 21364 26988
rect 20588 26948 21364 26976
rect 20588 26936 20594 26948
rect 21358 26936 21364 26948
rect 21416 26936 21422 26988
rect 21637 26979 21695 26985
rect 21637 26945 21649 26979
rect 21683 26976 21695 26979
rect 23216 26976 23244 27007
rect 21683 26948 23244 26976
rect 23845 26979 23903 26985
rect 21683 26945 21695 26948
rect 21637 26939 21695 26945
rect 23845 26945 23857 26979
rect 23891 26976 23903 26979
rect 24228 26976 24256 27072
rect 25774 27044 25780 27056
rect 23891 26948 24256 26976
rect 23891 26945 23903 26948
rect 23845 26939 23903 26945
rect 16301 26911 16359 26917
rect 16301 26908 16313 26911
rect 15304 26880 16313 26908
rect 16301 26877 16313 26880
rect 16347 26877 16359 26911
rect 16301 26871 16359 26877
rect 17310 26868 17316 26920
rect 17368 26868 17374 26920
rect 24118 26908 24124 26920
rect 22940 26880 24124 26908
rect 12069 26843 12127 26849
rect 11440 26812 11744 26840
rect 7834 26772 7840 26784
rect 6840 26744 7840 26772
rect 6733 26735 6791 26741
rect 7834 26732 7840 26744
rect 7892 26732 7898 26784
rect 9858 26732 9864 26784
rect 9916 26732 9922 26784
rect 10042 26732 10048 26784
rect 10100 26772 10106 26784
rect 11440 26772 11468 26812
rect 10100 26744 11468 26772
rect 11716 26772 11744 26812
rect 12069 26809 12081 26843
rect 12115 26840 12127 26843
rect 12342 26840 12348 26852
rect 12115 26812 12348 26840
rect 12115 26809 12127 26812
rect 12069 26803 12127 26809
rect 12342 26800 12348 26812
rect 12400 26800 12406 26852
rect 12434 26800 12440 26852
rect 12492 26840 12498 26852
rect 14936 26840 14964 26868
rect 15565 26843 15623 26849
rect 15565 26840 15577 26843
rect 12492 26812 15577 26840
rect 12492 26800 12498 26812
rect 15565 26809 15577 26812
rect 15611 26840 15623 26843
rect 16025 26843 16083 26849
rect 16025 26840 16037 26843
rect 15611 26812 16037 26840
rect 15611 26809 15623 26812
rect 15565 26803 15623 26809
rect 16025 26809 16037 26812
rect 16071 26840 16083 26843
rect 17126 26840 17132 26852
rect 16071 26812 17132 26840
rect 16071 26809 16083 26812
rect 16025 26803 16083 26809
rect 17126 26800 17132 26812
rect 17184 26840 17190 26852
rect 17184 26812 17540 26840
rect 17184 26800 17190 26812
rect 17512 26784 17540 26812
rect 19058 26800 19064 26852
rect 19116 26800 19122 26852
rect 19518 26800 19524 26852
rect 19576 26840 19582 26852
rect 19576 26812 20208 26840
rect 19576 26800 19582 26812
rect 12618 26772 12624 26784
rect 11716 26744 12624 26772
rect 10100 26732 10106 26744
rect 12618 26732 12624 26744
rect 12676 26732 12682 26784
rect 13909 26775 13967 26781
rect 13909 26741 13921 26775
rect 13955 26772 13967 26775
rect 14918 26772 14924 26784
rect 13955 26744 14924 26772
rect 13955 26741 13967 26744
rect 13909 26735 13967 26741
rect 14918 26732 14924 26744
rect 14976 26732 14982 26784
rect 16666 26732 16672 26784
rect 16724 26732 16730 26784
rect 17494 26732 17500 26784
rect 17552 26732 17558 26784
rect 18325 26775 18383 26781
rect 18325 26741 18337 26775
rect 18371 26772 18383 26775
rect 20070 26772 20076 26784
rect 18371 26744 20076 26772
rect 18371 26741 18383 26744
rect 18325 26735 18383 26741
rect 20070 26732 20076 26744
rect 20128 26732 20134 26784
rect 20180 26772 20208 26812
rect 22094 26800 22100 26852
rect 22152 26800 22158 26852
rect 22940 26772 22968 26880
rect 24118 26868 24124 26880
rect 24176 26868 24182 26920
rect 24228 26908 24256 26948
rect 24688 27016 25780 27044
rect 24397 26911 24455 26917
rect 24397 26908 24409 26911
rect 24228 26880 24409 26908
rect 24397 26877 24409 26880
rect 24443 26877 24455 26911
rect 24397 26871 24455 26877
rect 24486 26868 24492 26920
rect 24544 26868 24550 26920
rect 23566 26800 23572 26852
rect 23624 26800 23630 26852
rect 24213 26843 24271 26849
rect 24213 26809 24225 26843
rect 24259 26840 24271 26843
rect 24688 26840 24716 27016
rect 25774 27004 25780 27016
rect 25832 27004 25838 27056
rect 25866 27004 25872 27056
rect 25924 27004 25930 27056
rect 28092 27044 28120 27084
rect 29822 27072 29828 27084
rect 29880 27072 29886 27124
rect 30834 27072 30840 27124
rect 30892 27112 30898 27124
rect 31021 27115 31079 27121
rect 31021 27112 31033 27115
rect 30892 27084 31033 27112
rect 30892 27072 30898 27084
rect 31021 27081 31033 27084
rect 31067 27081 31079 27115
rect 31021 27075 31079 27081
rect 27356 27016 28120 27044
rect 25593 26979 25651 26985
rect 25593 26945 25605 26979
rect 25639 26976 25651 26979
rect 25682 26976 25688 26988
rect 25639 26948 25688 26976
rect 25639 26945 25651 26948
rect 25593 26939 25651 26945
rect 25682 26936 25688 26948
rect 25740 26936 25746 26988
rect 25406 26868 25412 26920
rect 25464 26868 25470 26920
rect 25883 26917 25911 27004
rect 27356 26976 27384 27016
rect 28902 27004 28908 27056
rect 28960 27004 28966 27056
rect 29641 27047 29699 27053
rect 29641 27013 29653 27047
rect 29687 27013 29699 27047
rect 29641 27007 29699 27013
rect 28920 26976 28948 27004
rect 25976 26948 27384 26976
rect 27448 26948 28948 26976
rect 29089 26979 29147 26985
rect 25869 26911 25927 26917
rect 25869 26877 25881 26911
rect 25915 26877 25927 26911
rect 25869 26871 25927 26877
rect 24259 26812 24716 26840
rect 24765 26843 24823 26849
rect 24259 26809 24271 26812
rect 24213 26803 24271 26809
rect 24765 26809 24777 26843
rect 24811 26840 24823 26843
rect 24854 26840 24860 26852
rect 24811 26812 24860 26840
rect 24811 26809 24823 26812
rect 24765 26803 24823 26809
rect 24854 26800 24860 26812
rect 24912 26800 24918 26852
rect 25038 26800 25044 26852
rect 25096 26840 25102 26852
rect 25976 26840 26004 26948
rect 26053 26911 26111 26917
rect 26053 26877 26065 26911
rect 26099 26877 26111 26911
rect 27448 26894 27476 26948
rect 29089 26945 29101 26979
rect 29135 26945 29147 26979
rect 29656 26976 29684 27007
rect 30466 27004 30472 27056
rect 30524 27004 30530 27056
rect 30285 26979 30343 26985
rect 30285 26976 30297 26979
rect 29656 26948 30297 26976
rect 29089 26939 29147 26945
rect 30285 26945 30297 26948
rect 30331 26945 30343 26979
rect 30285 26939 30343 26945
rect 26053 26871 26111 26877
rect 25096 26812 26004 26840
rect 26068 26840 26096 26871
rect 27890 26868 27896 26920
rect 27948 26868 27954 26920
rect 28442 26868 28448 26920
rect 28500 26868 28506 26920
rect 28629 26911 28687 26917
rect 28629 26877 28641 26911
rect 28675 26877 28687 26911
rect 28629 26871 28687 26877
rect 28813 26911 28871 26917
rect 28813 26877 28825 26911
rect 28859 26877 28871 26911
rect 29104 26908 29132 26939
rect 30484 26908 30512 27004
rect 29104 26880 30512 26908
rect 28813 26871 28871 26877
rect 27908 26840 27936 26868
rect 28644 26840 28672 26871
rect 26068 26812 26188 26840
rect 27908 26812 28672 26840
rect 28828 26840 28856 26871
rect 30558 26868 30564 26920
rect 30616 26908 30622 26920
rect 30837 26911 30895 26917
rect 30837 26908 30849 26911
rect 30616 26880 30849 26908
rect 30616 26868 30622 26880
rect 30837 26877 30849 26880
rect 30883 26877 30895 26911
rect 30837 26871 30895 26877
rect 31757 26911 31815 26917
rect 31757 26877 31769 26911
rect 31803 26908 31815 26911
rect 33134 26908 33140 26920
rect 31803 26880 33140 26908
rect 31803 26877 31815 26880
rect 31757 26871 31815 26877
rect 33134 26868 33140 26880
rect 33192 26868 33198 26920
rect 28828 26812 29316 26840
rect 25096 26800 25102 26812
rect 26160 26784 26188 26812
rect 20180 26744 22968 26772
rect 23661 26775 23719 26781
rect 23661 26741 23673 26775
rect 23707 26772 23719 26775
rect 24486 26772 24492 26784
rect 23707 26744 24492 26772
rect 23707 26741 23719 26744
rect 23661 26735 23719 26741
rect 24486 26732 24492 26744
rect 24544 26732 24550 26784
rect 24581 26775 24639 26781
rect 24581 26741 24593 26775
rect 24627 26772 24639 26775
rect 24946 26772 24952 26784
rect 24627 26744 24952 26772
rect 24627 26741 24639 26744
rect 24581 26735 24639 26741
rect 24946 26732 24952 26744
rect 25004 26732 25010 26784
rect 25590 26732 25596 26784
rect 25648 26732 25654 26784
rect 26142 26732 26148 26784
rect 26200 26732 26206 26784
rect 26326 26732 26332 26784
rect 26384 26772 26390 26784
rect 27338 26772 27344 26784
rect 26384 26744 27344 26772
rect 26384 26732 26390 26744
rect 27338 26732 27344 26744
rect 27396 26732 27402 26784
rect 27890 26732 27896 26784
rect 27948 26732 27954 26784
rect 29288 26781 29316 26812
rect 30098 26800 30104 26852
rect 30156 26840 30162 26852
rect 30745 26843 30803 26849
rect 30745 26840 30757 26843
rect 30156 26812 30757 26840
rect 30156 26800 30162 26812
rect 30745 26809 30757 26812
rect 30791 26809 30803 26843
rect 30745 26803 30803 26809
rect 28721 26775 28779 26781
rect 28721 26741 28733 26775
rect 28767 26772 28779 26775
rect 29181 26775 29239 26781
rect 29181 26772 29193 26775
rect 28767 26744 29193 26772
rect 28767 26741 28779 26744
rect 28721 26735 28779 26741
rect 29181 26741 29193 26744
rect 29227 26741 29239 26775
rect 29181 26735 29239 26741
rect 29273 26775 29331 26781
rect 29273 26741 29285 26775
rect 29319 26772 29331 26775
rect 29362 26772 29368 26784
rect 29319 26744 29368 26772
rect 29319 26741 29331 26744
rect 29273 26735 29331 26741
rect 29362 26732 29368 26744
rect 29420 26732 29426 26784
rect 29454 26732 29460 26784
rect 29512 26772 29518 26784
rect 29733 26775 29791 26781
rect 29733 26772 29745 26775
rect 29512 26744 29745 26772
rect 29512 26732 29518 26744
rect 29733 26741 29745 26744
rect 29779 26741 29791 26775
rect 29733 26735 29791 26741
rect 30374 26732 30380 26784
rect 30432 26772 30438 26784
rect 30653 26775 30711 26781
rect 30653 26772 30665 26775
rect 30432 26744 30665 26772
rect 30432 26732 30438 26744
rect 30653 26741 30665 26744
rect 30699 26741 30711 26775
rect 30653 26735 30711 26741
rect 31386 26732 31392 26784
rect 31444 26772 31450 26784
rect 31481 26775 31539 26781
rect 31481 26772 31493 26775
rect 31444 26744 31493 26772
rect 31444 26732 31450 26744
rect 31481 26741 31493 26744
rect 31527 26741 31539 26775
rect 31481 26735 31539 26741
rect 2760 26682 32200 26704
rect 2760 26630 6946 26682
rect 6998 26630 7010 26682
rect 7062 26630 7074 26682
rect 7126 26630 7138 26682
rect 7190 26630 7202 26682
rect 7254 26630 14306 26682
rect 14358 26630 14370 26682
rect 14422 26630 14434 26682
rect 14486 26630 14498 26682
rect 14550 26630 14562 26682
rect 14614 26630 21666 26682
rect 21718 26630 21730 26682
rect 21782 26630 21794 26682
rect 21846 26630 21858 26682
rect 21910 26630 21922 26682
rect 21974 26630 29026 26682
rect 29078 26630 29090 26682
rect 29142 26630 29154 26682
rect 29206 26630 29218 26682
rect 29270 26630 29282 26682
rect 29334 26630 32200 26682
rect 2760 26608 32200 26630
rect 5629 26571 5687 26577
rect 5629 26537 5641 26571
rect 5675 26568 5687 26571
rect 6822 26568 6828 26580
rect 5675 26540 6828 26568
rect 5675 26537 5687 26540
rect 5629 26531 5687 26537
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 7742 26528 7748 26580
rect 7800 26528 7806 26580
rect 8021 26571 8079 26577
rect 8021 26537 8033 26571
rect 8067 26537 8079 26571
rect 8021 26531 8079 26537
rect 4448 26472 5856 26500
rect 4448 26441 4476 26472
rect 5828 26444 5856 26472
rect 6638 26460 6644 26512
rect 6696 26460 6702 26512
rect 7101 26503 7159 26509
rect 7101 26469 7113 26503
rect 7147 26500 7159 26503
rect 8036 26500 8064 26531
rect 8386 26528 8392 26580
rect 8444 26528 8450 26580
rect 8481 26571 8539 26577
rect 8481 26537 8493 26571
rect 8527 26568 8539 26571
rect 8754 26568 8760 26580
rect 8527 26540 8760 26568
rect 8527 26537 8539 26540
rect 8481 26531 8539 26537
rect 8754 26528 8760 26540
rect 8812 26528 8818 26580
rect 8849 26571 8907 26577
rect 8849 26537 8861 26571
rect 8895 26568 8907 26571
rect 9398 26568 9404 26580
rect 8895 26540 9404 26568
rect 8895 26537 8907 26540
rect 8849 26531 8907 26537
rect 9398 26528 9404 26540
rect 9456 26528 9462 26580
rect 10318 26528 10324 26580
rect 10376 26568 10382 26580
rect 10505 26571 10563 26577
rect 10505 26568 10517 26571
rect 10376 26540 10517 26568
rect 10376 26528 10382 26540
rect 10505 26537 10517 26540
rect 10551 26568 10563 26571
rect 10594 26568 10600 26580
rect 10551 26540 10600 26568
rect 10551 26537 10563 26540
rect 10505 26531 10563 26537
rect 10594 26528 10600 26540
rect 10652 26528 10658 26580
rect 11238 26568 11244 26580
rect 10796 26540 11244 26568
rect 7147 26472 8064 26500
rect 8772 26500 8800 26528
rect 9125 26503 9183 26509
rect 9125 26500 9137 26503
rect 8772 26472 9137 26500
rect 7147 26469 7159 26472
rect 7101 26463 7159 26469
rect 9125 26469 9137 26472
rect 9171 26469 9183 26503
rect 9125 26463 9183 26469
rect 9217 26503 9275 26509
rect 9217 26469 9229 26503
rect 9263 26500 9275 26503
rect 9306 26500 9312 26512
rect 9263 26472 9312 26500
rect 9263 26469 9275 26472
rect 9217 26463 9275 26469
rect 9306 26460 9312 26472
rect 9364 26500 9370 26512
rect 10689 26503 10747 26509
rect 10689 26500 10701 26503
rect 9364 26472 10701 26500
rect 9364 26460 9370 26472
rect 10689 26469 10701 26472
rect 10735 26469 10747 26503
rect 10689 26463 10747 26469
rect 4433 26435 4491 26441
rect 4433 26401 4445 26435
rect 4479 26401 4491 26435
rect 4433 26395 4491 26401
rect 4522 26392 4528 26444
rect 4580 26392 4586 26444
rect 5810 26392 5816 26444
rect 5868 26392 5874 26444
rect 7834 26392 7840 26444
rect 7892 26432 7898 26444
rect 7892 26404 8708 26432
rect 7892 26392 7898 26404
rect 3234 26324 3240 26376
rect 3292 26324 3298 26376
rect 7374 26324 7380 26376
rect 7432 26364 7438 26376
rect 8478 26364 8484 26376
rect 7432 26336 8484 26364
rect 7432 26324 7438 26336
rect 8478 26324 8484 26336
rect 8536 26324 8542 26376
rect 8573 26367 8631 26373
rect 8573 26333 8585 26367
rect 8619 26333 8631 26367
rect 8680 26364 8708 26404
rect 9030 26392 9036 26444
rect 9088 26392 9094 26444
rect 9401 26435 9459 26441
rect 9401 26432 9413 26435
rect 9232 26404 9413 26432
rect 9232 26364 9260 26404
rect 9401 26401 9413 26404
rect 9447 26401 9459 26435
rect 9401 26395 9459 26401
rect 10594 26392 10600 26444
rect 10652 26392 10658 26444
rect 10796 26441 10824 26540
rect 11238 26528 11244 26540
rect 11296 26568 11302 26580
rect 12253 26571 12311 26577
rect 11296 26540 12204 26568
rect 11296 26528 11302 26540
rect 12176 26512 12204 26540
rect 12253 26537 12265 26571
rect 12299 26568 12311 26571
rect 12434 26568 12440 26580
rect 12299 26540 12440 26568
rect 12299 26537 12311 26540
rect 12253 26531 12311 26537
rect 10870 26460 10876 26512
rect 10928 26500 10934 26512
rect 11517 26503 11575 26509
rect 11517 26500 11529 26503
rect 10928 26472 11529 26500
rect 10928 26460 10934 26472
rect 11517 26469 11529 26472
rect 11563 26469 11575 26503
rect 11517 26463 11575 26469
rect 12158 26460 12164 26512
rect 12216 26460 12222 26512
rect 10781 26435 10839 26441
rect 10781 26401 10793 26435
rect 10827 26401 10839 26435
rect 11333 26435 11391 26441
rect 11333 26432 11345 26435
rect 10781 26395 10839 26401
rect 10888 26404 11345 26432
rect 10888 26364 10916 26404
rect 11333 26401 11345 26404
rect 11379 26401 11391 26435
rect 11333 26395 11391 26401
rect 11422 26392 11428 26444
rect 11480 26392 11486 26444
rect 11606 26392 11612 26444
rect 11664 26392 11670 26444
rect 11701 26435 11759 26441
rect 11701 26401 11713 26435
rect 11747 26432 11759 26435
rect 12268 26432 12296 26531
rect 12434 26528 12440 26540
rect 12492 26528 12498 26580
rect 14826 26528 14832 26580
rect 14884 26568 14890 26580
rect 14921 26571 14979 26577
rect 14921 26568 14933 26571
rect 14884 26540 14933 26568
rect 14884 26528 14890 26540
rect 14921 26537 14933 26540
rect 14967 26537 14979 26571
rect 14921 26531 14979 26537
rect 15194 26528 15200 26580
rect 15252 26568 15258 26580
rect 15378 26568 15384 26580
rect 15252 26540 15384 26568
rect 15252 26528 15258 26540
rect 15378 26528 15384 26540
rect 15436 26528 15442 26580
rect 17034 26528 17040 26580
rect 17092 26528 17098 26580
rect 18141 26571 18199 26577
rect 18141 26537 18153 26571
rect 18187 26568 18199 26571
rect 19242 26568 19248 26580
rect 18187 26540 19248 26568
rect 18187 26537 18199 26540
rect 18141 26531 18199 26537
rect 19242 26528 19248 26540
rect 19300 26528 19306 26580
rect 19337 26571 19395 26577
rect 19337 26537 19349 26571
rect 19383 26568 19395 26571
rect 19518 26568 19524 26580
rect 19383 26540 19524 26568
rect 19383 26537 19395 26540
rect 19337 26531 19395 26537
rect 19518 26528 19524 26540
rect 19576 26528 19582 26580
rect 19705 26571 19763 26577
rect 19705 26537 19717 26571
rect 19751 26537 19763 26571
rect 19705 26531 19763 26537
rect 13262 26460 13268 26512
rect 13320 26500 13326 26512
rect 14734 26500 14740 26512
rect 13320 26472 14740 26500
rect 13320 26460 13326 26472
rect 14734 26460 14740 26472
rect 14792 26500 14798 26512
rect 17052 26500 17080 26528
rect 18417 26503 18475 26509
rect 18417 26500 18429 26503
rect 14792 26472 17080 26500
rect 17894 26472 18429 26500
rect 14792 26460 14798 26472
rect 11747 26404 12296 26432
rect 11747 26401 11759 26404
rect 11701 26395 11759 26401
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 16408 26441 16436 26472
rect 18417 26469 18429 26472
rect 18463 26469 18475 26503
rect 19150 26500 19156 26512
rect 18417 26463 18475 26469
rect 18984 26472 19156 26500
rect 15197 26435 15255 26441
rect 15197 26432 15209 26435
rect 12676 26404 15209 26432
rect 12676 26392 12682 26404
rect 15197 26401 15209 26404
rect 15243 26432 15255 26435
rect 15933 26435 15991 26441
rect 15933 26432 15945 26435
rect 15243 26404 15945 26432
rect 15243 26401 15255 26404
rect 15197 26395 15255 26401
rect 15933 26401 15945 26404
rect 15979 26401 15991 26435
rect 15933 26395 15991 26401
rect 16393 26435 16451 26441
rect 16393 26401 16405 26435
rect 16439 26401 16451 26435
rect 16393 26395 16451 26401
rect 18509 26435 18567 26441
rect 18509 26401 18521 26435
rect 18555 26432 18567 26435
rect 18874 26432 18880 26444
rect 18555 26404 18880 26432
rect 18555 26401 18567 26404
rect 18509 26395 18567 26401
rect 8680 26336 9168 26364
rect 8573 26327 8631 26333
rect 5166 26188 5172 26240
rect 5224 26188 5230 26240
rect 8110 26188 8116 26240
rect 8168 26228 8174 26240
rect 8588 26228 8616 26327
rect 8168 26200 8616 26228
rect 9140 26228 9168 26336
rect 9232 26336 10916 26364
rect 11149 26367 11207 26373
rect 9232 26308 9260 26336
rect 11149 26333 11161 26367
rect 11195 26364 11207 26367
rect 11440 26364 11468 26392
rect 11195 26336 11468 26364
rect 11195 26333 11207 26336
rect 11149 26327 11207 26333
rect 13354 26324 13360 26376
rect 13412 26324 13418 26376
rect 14182 26324 14188 26376
rect 14240 26364 14246 26376
rect 14277 26367 14335 26373
rect 14277 26364 14289 26367
rect 14240 26336 14289 26364
rect 14240 26324 14246 26336
rect 14277 26333 14289 26336
rect 14323 26333 14335 26367
rect 15948 26364 15976 26395
rect 18874 26392 18880 26404
rect 18932 26392 18938 26444
rect 15948 26336 16528 26364
rect 14277 26327 14335 26333
rect 9214 26256 9220 26308
rect 9272 26256 9278 26308
rect 10137 26299 10195 26305
rect 9324 26268 10088 26296
rect 9324 26228 9352 26268
rect 10060 26240 10088 26268
rect 10137 26265 10149 26299
rect 10183 26296 10195 26299
rect 14001 26299 14059 26305
rect 10183 26268 12434 26296
rect 10183 26265 10195 26268
rect 10137 26259 10195 26265
rect 9140 26200 9352 26228
rect 8168 26188 8174 26200
rect 9582 26188 9588 26240
rect 9640 26228 9646 26240
rect 9677 26231 9735 26237
rect 9677 26228 9689 26231
rect 9640 26200 9689 26228
rect 9640 26188 9646 26200
rect 9677 26197 9689 26200
rect 9723 26197 9735 26231
rect 9677 26191 9735 26197
rect 10042 26188 10048 26240
rect 10100 26188 10106 26240
rect 10502 26188 10508 26240
rect 10560 26228 10566 26240
rect 11514 26228 11520 26240
rect 10560 26200 11520 26228
rect 10560 26188 10566 26200
rect 11514 26188 11520 26200
rect 11572 26188 11578 26240
rect 11882 26188 11888 26240
rect 11940 26188 11946 26240
rect 12406 26228 12434 26268
rect 14001 26265 14013 26299
rect 14047 26296 14059 26299
rect 14642 26296 14648 26308
rect 14047 26268 14648 26296
rect 14047 26265 14059 26268
rect 14001 26259 14059 26265
rect 14642 26256 14648 26268
rect 14700 26256 14706 26308
rect 15562 26296 15568 26308
rect 15028 26268 15568 26296
rect 13446 26228 13452 26240
rect 12406 26200 13452 26228
rect 13446 26188 13452 26200
rect 13504 26228 13510 26240
rect 15028 26228 15056 26268
rect 15562 26256 15568 26268
rect 15620 26256 15626 26308
rect 13504 26200 15056 26228
rect 13504 26188 13510 26200
rect 15102 26188 15108 26240
rect 15160 26188 15166 26240
rect 15930 26188 15936 26240
rect 15988 26228 15994 26240
rect 16025 26231 16083 26237
rect 16025 26228 16037 26231
rect 15988 26200 16037 26228
rect 15988 26188 15994 26200
rect 16025 26197 16037 26200
rect 16071 26197 16083 26231
rect 16500 26228 16528 26336
rect 16666 26324 16672 26376
rect 16724 26324 16730 26376
rect 18414 26324 18420 26376
rect 18472 26364 18478 26376
rect 18984 26364 19012 26472
rect 19150 26460 19156 26472
rect 19208 26500 19214 26512
rect 19720 26500 19748 26531
rect 19794 26528 19800 26580
rect 19852 26528 19858 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 20165 26571 20223 26577
rect 20165 26568 20177 26571
rect 20128 26540 20177 26568
rect 20128 26528 20134 26540
rect 20165 26537 20177 26540
rect 20211 26568 20223 26571
rect 22186 26568 22192 26580
rect 20211 26540 21404 26568
rect 20211 26537 20223 26540
rect 20165 26531 20223 26537
rect 19208 26472 19564 26500
rect 19720 26472 20484 26500
rect 19208 26460 19214 26472
rect 19536 26432 19564 26472
rect 20257 26435 20315 26441
rect 20257 26432 20269 26435
rect 19536 26404 20269 26432
rect 20257 26401 20269 26404
rect 20303 26401 20315 26435
rect 20257 26395 20315 26401
rect 18472 26336 19012 26364
rect 19061 26367 19119 26373
rect 18472 26324 18478 26336
rect 19061 26333 19073 26367
rect 19107 26333 19119 26367
rect 19061 26327 19119 26333
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26364 19303 26367
rect 19426 26364 19432 26376
rect 19291 26336 19432 26364
rect 19291 26333 19303 26336
rect 19245 26327 19303 26333
rect 16758 26228 16764 26240
rect 16500 26200 16764 26228
rect 16025 26191 16083 26197
rect 16758 26188 16764 26200
rect 16816 26188 16822 26240
rect 18506 26188 18512 26240
rect 18564 26228 18570 26240
rect 18785 26231 18843 26237
rect 18785 26228 18797 26231
rect 18564 26200 18797 26228
rect 18564 26188 18570 26200
rect 18785 26197 18797 26200
rect 18831 26228 18843 26231
rect 19076 26228 19104 26327
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 20349 26367 20407 26373
rect 19628 26336 20116 26364
rect 19628 26228 19656 26336
rect 20088 26308 20116 26336
rect 20349 26333 20361 26367
rect 20395 26333 20407 26367
rect 20456 26364 20484 26472
rect 21177 26367 21235 26373
rect 21177 26364 21189 26367
rect 20456 26336 21189 26364
rect 20349 26327 20407 26333
rect 21177 26333 21189 26336
rect 21223 26333 21235 26367
rect 21376 26364 21404 26540
rect 21836 26540 22192 26568
rect 21836 26509 21864 26540
rect 22186 26528 22192 26540
rect 22244 26528 22250 26580
rect 23293 26571 23351 26577
rect 23293 26537 23305 26571
rect 23339 26568 23351 26571
rect 23382 26568 23388 26580
rect 23339 26540 23388 26568
rect 23339 26537 23351 26540
rect 23293 26531 23351 26537
rect 23382 26528 23388 26540
rect 23440 26528 23446 26580
rect 25038 26568 25044 26580
rect 23492 26540 25044 26568
rect 21821 26503 21879 26509
rect 21821 26469 21833 26503
rect 21867 26469 21879 26503
rect 21821 26463 21879 26469
rect 22462 26460 22468 26512
rect 22520 26460 22526 26512
rect 23492 26500 23520 26540
rect 25038 26528 25044 26540
rect 25096 26528 25102 26580
rect 25225 26571 25283 26577
rect 25225 26537 25237 26571
rect 25271 26568 25283 26571
rect 25406 26568 25412 26580
rect 25271 26540 25412 26568
rect 25271 26537 25283 26540
rect 25225 26531 25283 26537
rect 25406 26528 25412 26540
rect 25464 26528 25470 26580
rect 26237 26571 26295 26577
rect 26237 26537 26249 26571
rect 26283 26568 26295 26571
rect 26878 26568 26884 26580
rect 26283 26540 26884 26568
rect 26283 26537 26295 26540
rect 26237 26531 26295 26537
rect 26878 26528 26884 26540
rect 26936 26528 26942 26580
rect 27338 26568 27344 26580
rect 27080 26540 27344 26568
rect 25682 26500 25688 26512
rect 23400 26472 23520 26500
rect 24978 26472 25688 26500
rect 21450 26392 21456 26444
rect 21508 26432 21514 26444
rect 21545 26435 21603 26441
rect 21545 26432 21557 26435
rect 21508 26404 21557 26432
rect 21508 26392 21514 26404
rect 21545 26401 21557 26404
rect 21591 26401 21603 26435
rect 21545 26395 21603 26401
rect 23400 26364 23428 26472
rect 25682 26460 25688 26472
rect 25740 26460 25746 26512
rect 26326 26500 26332 26512
rect 25884 26472 26332 26500
rect 23474 26392 23480 26444
rect 23532 26392 23538 26444
rect 25593 26435 25651 26441
rect 25593 26401 25605 26435
rect 25639 26432 25651 26435
rect 25884 26432 25912 26472
rect 26326 26460 26332 26472
rect 26384 26460 26390 26512
rect 26510 26460 26516 26512
rect 26568 26460 26574 26512
rect 26602 26460 26608 26512
rect 26660 26460 26666 26512
rect 26786 26509 26792 26512
rect 26743 26503 26792 26509
rect 26743 26469 26755 26503
rect 26789 26469 26792 26503
rect 26743 26463 26792 26469
rect 26786 26460 26792 26463
rect 26844 26460 26850 26512
rect 25639 26404 25912 26432
rect 25961 26435 26019 26441
rect 25639 26401 25651 26404
rect 25593 26395 25651 26401
rect 25961 26401 25973 26435
rect 26007 26401 26019 26435
rect 25961 26395 26019 26401
rect 26421 26435 26479 26441
rect 26421 26401 26433 26435
rect 26467 26430 26479 26435
rect 26881 26435 26939 26441
rect 26467 26402 26648 26430
rect 26467 26401 26479 26402
rect 26421 26395 26479 26401
rect 21376 26336 23428 26364
rect 23753 26367 23811 26373
rect 21177 26327 21235 26333
rect 23753 26333 23765 26367
rect 23799 26364 23811 26367
rect 25222 26364 25228 26376
rect 23799 26336 25228 26364
rect 23799 26333 23811 26336
rect 23753 26327 23811 26333
rect 20070 26256 20076 26308
rect 20128 26296 20134 26308
rect 20364 26296 20392 26327
rect 25222 26324 25228 26336
rect 25280 26324 25286 26376
rect 25501 26367 25559 26373
rect 25501 26333 25513 26367
rect 25547 26333 25559 26367
rect 25976 26364 26004 26395
rect 26620 26364 26648 26402
rect 26881 26401 26893 26435
rect 26927 26432 26939 26435
rect 27080 26432 27108 26540
rect 27338 26528 27344 26540
rect 27396 26528 27402 26580
rect 27522 26528 27528 26580
rect 27580 26528 27586 26580
rect 27801 26571 27859 26577
rect 27801 26537 27813 26571
rect 27847 26568 27859 26571
rect 28442 26568 28448 26580
rect 27847 26540 28448 26568
rect 27847 26537 27859 26540
rect 27801 26531 27859 26537
rect 28442 26528 28448 26540
rect 28500 26528 28506 26580
rect 29454 26568 29460 26580
rect 29196 26540 29460 26568
rect 27157 26503 27215 26509
rect 27157 26469 27169 26503
rect 27203 26500 27215 26503
rect 29086 26500 29092 26512
rect 27203 26472 29092 26500
rect 27203 26469 27215 26472
rect 27157 26463 27215 26469
rect 26927 26404 27108 26432
rect 26927 26401 26939 26404
rect 26881 26395 26939 26401
rect 26970 26364 26976 26376
rect 25976 26336 26556 26364
rect 26620 26336 26976 26364
rect 25501 26327 25559 26333
rect 20128 26268 20392 26296
rect 20128 26256 20134 26268
rect 24946 26256 24952 26308
rect 25004 26296 25010 26308
rect 25516 26296 25544 26327
rect 25004 26268 25544 26296
rect 26145 26299 26203 26305
rect 25004 26256 25010 26268
rect 26145 26265 26157 26299
rect 26191 26296 26203 26299
rect 26418 26296 26424 26308
rect 26191 26268 26424 26296
rect 26191 26265 26203 26268
rect 26145 26259 26203 26265
rect 26418 26256 26424 26268
rect 26476 26256 26482 26308
rect 26528 26296 26556 26336
rect 26970 26324 26976 26336
rect 27028 26324 27034 26376
rect 27172 26296 27200 26463
rect 27433 26435 27491 26441
rect 27433 26401 27445 26435
rect 27479 26432 27491 26435
rect 27798 26432 27804 26444
rect 27479 26404 27804 26432
rect 27479 26401 27491 26404
rect 27433 26395 27491 26401
rect 27798 26392 27804 26404
rect 27856 26392 27862 26444
rect 27985 26435 28043 26441
rect 27985 26401 27997 26435
rect 28031 26401 28043 26435
rect 27985 26395 28043 26401
rect 26528 26268 27200 26296
rect 27706 26256 27712 26308
rect 27764 26296 27770 26308
rect 28000 26296 28028 26395
rect 28258 26392 28264 26444
rect 28316 26392 28322 26444
rect 28460 26441 28488 26472
rect 29086 26460 29092 26472
rect 29144 26460 29150 26512
rect 29196 26509 29224 26540
rect 29454 26528 29460 26540
rect 29512 26528 29518 26580
rect 30650 26528 30656 26580
rect 30708 26528 30714 26580
rect 29181 26503 29239 26509
rect 29181 26469 29193 26503
rect 29227 26469 29239 26503
rect 30837 26503 30895 26509
rect 30837 26500 30849 26503
rect 30406 26472 30849 26500
rect 29181 26463 29239 26469
rect 30837 26469 30849 26472
rect 30883 26469 30895 26503
rect 30837 26463 30895 26469
rect 28445 26435 28503 26441
rect 28445 26401 28457 26435
rect 28491 26401 28503 26435
rect 28445 26395 28503 26401
rect 28626 26392 28632 26444
rect 28684 26392 28690 26444
rect 28810 26392 28816 26444
rect 28868 26392 28874 26444
rect 30926 26392 30932 26444
rect 30984 26392 30990 26444
rect 28166 26324 28172 26376
rect 28224 26364 28230 26376
rect 28644 26364 28672 26392
rect 28905 26367 28963 26373
rect 28905 26364 28917 26367
rect 28224 26336 28917 26364
rect 28224 26324 28230 26336
rect 28905 26333 28917 26336
rect 28951 26333 28963 26367
rect 30944 26364 30972 26392
rect 28905 26327 28963 26333
rect 30300 26336 30972 26364
rect 30300 26308 30328 26336
rect 27764 26268 28948 26296
rect 27764 26256 27770 26268
rect 28920 26240 28948 26268
rect 30282 26256 30288 26308
rect 30340 26256 30346 26308
rect 18831 26200 19656 26228
rect 18831 26197 18843 26200
rect 18785 26191 18843 26197
rect 20622 26188 20628 26240
rect 20680 26188 20686 26240
rect 24854 26188 24860 26240
rect 24912 26228 24918 26240
rect 25869 26231 25927 26237
rect 25869 26228 25881 26231
rect 24912 26200 25881 26228
rect 24912 26188 24918 26200
rect 25869 26197 25881 26200
rect 25915 26197 25927 26231
rect 25869 26191 25927 26197
rect 28721 26231 28779 26237
rect 28721 26197 28733 26231
rect 28767 26228 28779 26231
rect 28810 26228 28816 26240
rect 28767 26200 28816 26228
rect 28767 26197 28779 26200
rect 28721 26191 28779 26197
rect 28810 26188 28816 26200
rect 28868 26188 28874 26240
rect 28902 26188 28908 26240
rect 28960 26188 28966 26240
rect 2760 26138 32200 26160
rect 2760 26086 6286 26138
rect 6338 26086 6350 26138
rect 6402 26086 6414 26138
rect 6466 26086 6478 26138
rect 6530 26086 6542 26138
rect 6594 26086 13646 26138
rect 13698 26086 13710 26138
rect 13762 26086 13774 26138
rect 13826 26086 13838 26138
rect 13890 26086 13902 26138
rect 13954 26086 21006 26138
rect 21058 26086 21070 26138
rect 21122 26086 21134 26138
rect 21186 26086 21198 26138
rect 21250 26086 21262 26138
rect 21314 26086 28366 26138
rect 28418 26086 28430 26138
rect 28482 26086 28494 26138
rect 28546 26086 28558 26138
rect 28610 26086 28622 26138
rect 28674 26086 32200 26138
rect 2760 26064 32200 26086
rect 3513 26027 3571 26033
rect 3513 25993 3525 26027
rect 3559 26024 3571 26027
rect 4522 26024 4528 26036
rect 3559 25996 4528 26024
rect 3559 25993 3571 25996
rect 3513 25987 3571 25993
rect 4522 25984 4528 25996
rect 4580 25984 4586 26036
rect 9030 25984 9036 26036
rect 9088 26024 9094 26036
rect 9582 26024 9588 26036
rect 9088 25996 9588 26024
rect 9088 25984 9094 25996
rect 9582 25984 9588 25996
rect 9640 25984 9646 26036
rect 10318 25984 10324 26036
rect 10376 25984 10382 26036
rect 10870 25984 10876 26036
rect 10928 25984 10934 26036
rect 11606 25984 11612 26036
rect 11664 26024 11670 26036
rect 12161 26027 12219 26033
rect 12161 26024 12173 26027
rect 11664 25996 12173 26024
rect 11664 25984 11670 25996
rect 12161 25993 12173 25996
rect 12207 26024 12219 26027
rect 12207 25996 16574 26024
rect 12207 25993 12219 25996
rect 12161 25987 12219 25993
rect 4246 25848 4252 25900
rect 4304 25888 4310 25900
rect 5261 25891 5319 25897
rect 5261 25888 5273 25891
rect 4304 25860 5273 25888
rect 4304 25848 4310 25860
rect 5261 25857 5273 25860
rect 5307 25857 5319 25891
rect 5261 25851 5319 25857
rect 5810 25848 5816 25900
rect 5868 25888 5874 25900
rect 6733 25891 6791 25897
rect 6733 25888 6745 25891
rect 5868 25860 6745 25888
rect 5868 25848 5874 25860
rect 6733 25857 6745 25860
rect 6779 25888 6791 25891
rect 9861 25891 9919 25897
rect 9861 25888 9873 25891
rect 6779 25860 9873 25888
rect 6779 25857 6791 25860
rect 6733 25851 6791 25857
rect 9861 25857 9873 25860
rect 9907 25857 9919 25891
rect 9861 25851 9919 25857
rect 8478 25780 8484 25832
rect 8536 25780 8542 25832
rect 9217 25823 9275 25829
rect 9217 25789 9229 25823
rect 9263 25820 9275 25823
rect 9398 25820 9404 25832
rect 9263 25792 9404 25820
rect 9263 25789 9275 25792
rect 9217 25783 9275 25789
rect 9398 25780 9404 25792
rect 9456 25780 9462 25832
rect 4554 25724 4936 25752
rect 4908 25684 4936 25724
rect 4982 25712 4988 25764
rect 5040 25712 5046 25764
rect 7742 25712 7748 25764
rect 7800 25712 7806 25764
rect 8202 25712 8208 25764
rect 8260 25712 8266 25764
rect 5258 25684 5264 25696
rect 4908 25656 5264 25684
rect 5258 25644 5264 25656
rect 5316 25644 5322 25696
rect 5626 25644 5632 25696
rect 5684 25644 5690 25696
rect 6178 25644 6184 25696
rect 6236 25644 6242 25696
rect 7282 25644 7288 25696
rect 7340 25684 7346 25696
rect 7834 25684 7840 25696
rect 7340 25656 7840 25684
rect 7340 25644 7346 25656
rect 7834 25644 7840 25656
rect 7892 25644 7898 25696
rect 8570 25644 8576 25696
rect 8628 25644 8634 25696
rect 9306 25644 9312 25696
rect 9364 25644 9370 25696
rect 9582 25644 9588 25696
rect 9640 25684 9646 25696
rect 10336 25684 10364 25984
rect 10962 25916 10968 25968
rect 11020 25916 11026 25968
rect 16546 25956 16574 25996
rect 17310 25984 17316 26036
rect 17368 26024 17374 26036
rect 17773 26027 17831 26033
rect 17773 26024 17785 26027
rect 17368 25996 17785 26024
rect 17368 25984 17374 25996
rect 17773 25993 17785 25996
rect 17819 25993 17831 26027
rect 17773 25987 17831 25993
rect 18785 26027 18843 26033
rect 18785 25993 18797 26027
rect 18831 26024 18843 26027
rect 19702 26024 19708 26036
rect 18831 25996 19708 26024
rect 18831 25993 18843 25996
rect 18785 25987 18843 25993
rect 19702 25984 19708 25996
rect 19760 25984 19766 26036
rect 21450 25984 21456 26036
rect 21508 25984 21514 26036
rect 25222 25984 25228 26036
rect 25280 25984 25286 26036
rect 29362 25984 29368 26036
rect 29420 26024 29426 26036
rect 30101 26027 30159 26033
rect 30101 26024 30113 26027
rect 29420 25996 30113 26024
rect 29420 25984 29426 25996
rect 30101 25993 30113 25996
rect 30147 25993 30159 26027
rect 30101 25987 30159 25993
rect 20901 25959 20959 25965
rect 20901 25956 20913 25959
rect 16546 25928 19104 25956
rect 10980 25888 11008 25916
rect 10888 25860 11008 25888
rect 10594 25780 10600 25832
rect 10652 25820 10658 25832
rect 10689 25823 10747 25829
rect 10689 25820 10701 25823
rect 10652 25792 10701 25820
rect 10652 25780 10658 25792
rect 10689 25789 10701 25792
rect 10735 25820 10747 25823
rect 10778 25820 10784 25832
rect 10735 25792 10784 25820
rect 10735 25789 10747 25792
rect 10689 25783 10747 25789
rect 10778 25780 10784 25792
rect 10836 25780 10842 25832
rect 10888 25829 10916 25860
rect 11330 25848 11336 25900
rect 11388 25848 11394 25900
rect 12897 25891 12955 25897
rect 12897 25857 12909 25891
rect 12943 25888 12955 25891
rect 13262 25888 13268 25900
rect 12943 25860 13268 25888
rect 12943 25857 12955 25860
rect 12897 25851 12955 25857
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 14645 25891 14703 25897
rect 14645 25857 14657 25891
rect 14691 25888 14703 25891
rect 15286 25888 15292 25900
rect 14691 25860 15292 25888
rect 14691 25857 14703 25860
rect 14645 25851 14703 25857
rect 15286 25848 15292 25860
rect 15344 25848 15350 25900
rect 17034 25848 17040 25900
rect 17092 25848 17098 25900
rect 18414 25888 18420 25900
rect 17512 25860 18420 25888
rect 10873 25823 10931 25829
rect 10873 25789 10885 25823
rect 10919 25789 10931 25823
rect 10873 25783 10931 25789
rect 10965 25823 11023 25829
rect 10965 25789 10977 25823
rect 11011 25789 11023 25823
rect 11348 25820 11376 25848
rect 11609 25823 11667 25829
rect 11609 25820 11621 25823
rect 11348 25792 11621 25820
rect 10965 25783 11023 25789
rect 11609 25789 11621 25792
rect 11655 25789 11667 25823
rect 11609 25783 11667 25789
rect 9640 25656 10364 25684
rect 9640 25644 9646 25656
rect 10502 25644 10508 25696
rect 10560 25684 10566 25696
rect 10980 25684 11008 25783
rect 12802 25780 12808 25832
rect 12860 25780 12866 25832
rect 14734 25780 14740 25832
rect 14792 25780 14798 25832
rect 16298 25780 16304 25832
rect 16356 25780 16362 25832
rect 17218 25780 17224 25832
rect 17276 25780 17282 25832
rect 17512 25829 17540 25860
rect 18414 25848 18420 25860
rect 18472 25848 18478 25900
rect 19076 25888 19104 25928
rect 20456 25928 20913 25956
rect 19610 25888 19616 25900
rect 19076 25860 19616 25888
rect 19610 25848 19616 25860
rect 19668 25848 19674 25900
rect 19886 25848 19892 25900
rect 19944 25888 19950 25900
rect 20456 25888 20484 25928
rect 20901 25925 20913 25928
rect 20947 25925 20959 25959
rect 21468 25956 21496 25984
rect 21468 25928 22140 25956
rect 20901 25919 20959 25925
rect 22112 25897 22140 25928
rect 28902 25916 28908 25968
rect 28960 25956 28966 25968
rect 28960 25928 30328 25956
rect 28960 25916 28966 25928
rect 19944 25860 20484 25888
rect 22097 25891 22155 25897
rect 19944 25848 19950 25860
rect 22097 25857 22109 25891
rect 22143 25857 22155 25891
rect 22097 25851 22155 25857
rect 24765 25891 24823 25897
rect 24765 25857 24777 25891
rect 24811 25857 24823 25891
rect 27525 25891 27583 25897
rect 24765 25851 24823 25857
rect 25148 25860 26372 25888
rect 17497 25823 17555 25829
rect 17497 25789 17509 25823
rect 17543 25789 17555 25823
rect 17497 25783 17555 25789
rect 17589 25823 17647 25829
rect 17589 25789 17601 25823
rect 17635 25789 17647 25823
rect 17589 25783 17647 25789
rect 13170 25712 13176 25764
rect 13228 25712 13234 25764
rect 15102 25752 15108 25764
rect 14398 25724 15108 25752
rect 15102 25712 15108 25724
rect 15160 25712 15166 25764
rect 17405 25755 17463 25761
rect 17405 25752 17417 25755
rect 15212 25724 17417 25752
rect 10560 25656 11008 25684
rect 10560 25644 10566 25656
rect 11422 25644 11428 25696
rect 11480 25684 11486 25696
rect 11885 25687 11943 25693
rect 11885 25684 11897 25687
rect 11480 25656 11897 25684
rect 11480 25644 11486 25656
rect 11885 25653 11897 25656
rect 11931 25653 11943 25687
rect 11885 25647 11943 25653
rect 14090 25644 14096 25696
rect 14148 25684 14154 25696
rect 15212 25684 15240 25724
rect 17405 25721 17417 25724
rect 17451 25721 17463 25755
rect 17405 25715 17463 25721
rect 14148 25656 15240 25684
rect 14148 25644 14154 25656
rect 15470 25644 15476 25696
rect 15528 25684 15534 25696
rect 15749 25687 15807 25693
rect 15749 25684 15761 25687
rect 15528 25656 15761 25684
rect 15528 25644 15534 25656
rect 15749 25653 15761 25656
rect 15795 25653 15807 25687
rect 15749 25647 15807 25653
rect 16482 25644 16488 25696
rect 16540 25644 16546 25696
rect 17494 25644 17500 25696
rect 17552 25684 17558 25696
rect 17604 25684 17632 25783
rect 20530 25780 20536 25832
rect 20588 25780 20594 25832
rect 21450 25780 21456 25832
rect 21508 25780 21514 25832
rect 21821 25823 21879 25829
rect 21821 25789 21833 25823
rect 21867 25820 21879 25823
rect 21867 25792 22048 25820
rect 21867 25789 21879 25792
rect 21821 25783 21879 25789
rect 22020 25764 22048 25792
rect 20257 25755 20315 25761
rect 19826 25724 20208 25752
rect 18049 25687 18107 25693
rect 18049 25684 18061 25687
rect 17552 25656 18061 25684
rect 17552 25644 17558 25656
rect 18049 25653 18061 25656
rect 18095 25653 18107 25687
rect 18049 25647 18107 25653
rect 18506 25644 18512 25696
rect 18564 25644 18570 25696
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 19886 25684 19892 25696
rect 19484 25656 19892 25684
rect 19484 25644 19490 25656
rect 19886 25644 19892 25656
rect 19944 25644 19950 25696
rect 20180 25684 20208 25724
rect 20257 25721 20269 25755
rect 20303 25752 20315 25755
rect 20622 25752 20628 25764
rect 20303 25724 20628 25752
rect 20303 25721 20315 25724
rect 20257 25715 20315 25721
rect 20622 25712 20628 25724
rect 20680 25712 20686 25764
rect 21729 25755 21787 25761
rect 21729 25752 21741 25755
rect 20732 25724 21741 25752
rect 20732 25684 20760 25724
rect 21729 25721 21741 25724
rect 21775 25721 21787 25755
rect 21729 25715 21787 25721
rect 22002 25712 22008 25764
rect 22060 25712 22066 25764
rect 22112 25752 22140 25851
rect 23474 25780 23480 25832
rect 23532 25780 23538 25832
rect 22278 25752 22284 25764
rect 22112 25724 22284 25752
rect 22278 25712 22284 25724
rect 22336 25712 22342 25764
rect 22370 25712 22376 25764
rect 22428 25712 22434 25764
rect 24780 25752 24808 25851
rect 25148 25832 25176 25860
rect 26344 25832 26372 25860
rect 27525 25857 27537 25891
rect 27571 25888 27583 25891
rect 28166 25888 28172 25900
rect 27571 25860 28172 25888
rect 27571 25857 27583 25860
rect 27525 25851 27583 25857
rect 28166 25848 28172 25860
rect 28224 25848 28230 25900
rect 29273 25891 29331 25897
rect 29273 25857 29285 25891
rect 29319 25888 29331 25891
rect 29319 25860 29408 25888
rect 29319 25857 29331 25860
rect 29273 25851 29331 25857
rect 25130 25780 25136 25832
rect 25188 25780 25194 25832
rect 25314 25780 25320 25832
rect 25372 25820 25378 25832
rect 25777 25823 25835 25829
rect 25777 25820 25789 25823
rect 25372 25792 25789 25820
rect 25372 25780 25378 25792
rect 25777 25789 25789 25792
rect 25823 25789 25835 25823
rect 25777 25783 25835 25789
rect 25866 25780 25872 25832
rect 25924 25820 25930 25832
rect 25924 25792 26188 25820
rect 25924 25780 25930 25792
rect 26160 25761 26188 25792
rect 26326 25780 26332 25832
rect 26384 25780 26390 25832
rect 28810 25780 28816 25832
rect 28868 25820 28874 25832
rect 29380 25829 29408 25860
rect 30300 25829 30328 25928
rect 29365 25823 29423 25829
rect 28868 25792 28934 25820
rect 28868 25780 28874 25792
rect 29365 25789 29377 25823
rect 29411 25789 29423 25823
rect 29365 25783 29423 25789
rect 30285 25823 30343 25829
rect 30285 25789 30297 25823
rect 30331 25789 30343 25823
rect 30285 25783 30343 25789
rect 30374 25780 30380 25832
rect 30432 25780 30438 25832
rect 26145 25755 26203 25761
rect 24780 25724 25544 25752
rect 25516 25696 25544 25724
rect 26145 25721 26157 25755
rect 26191 25721 26203 25755
rect 26145 25715 26203 25721
rect 27801 25755 27859 25761
rect 27801 25721 27813 25755
rect 27847 25752 27859 25755
rect 27890 25752 27896 25764
rect 27847 25724 27896 25752
rect 27847 25721 27859 25724
rect 27801 25715 27859 25721
rect 27890 25712 27896 25724
rect 27948 25712 27954 25764
rect 30098 25712 30104 25764
rect 30156 25712 30162 25764
rect 20180 25656 20760 25684
rect 23842 25644 23848 25696
rect 23900 25644 23906 25696
rect 25498 25644 25504 25696
rect 25556 25644 25562 25696
rect 26237 25687 26295 25693
rect 26237 25653 26249 25687
rect 26283 25684 26295 25687
rect 26602 25684 26608 25696
rect 26283 25656 26608 25684
rect 26283 25653 26295 25656
rect 26237 25647 26295 25653
rect 26602 25644 26608 25656
rect 26660 25644 26666 25696
rect 29086 25644 29092 25696
rect 29144 25684 29150 25696
rect 29549 25687 29607 25693
rect 29549 25684 29561 25687
rect 29144 25656 29561 25684
rect 29144 25644 29150 25656
rect 29549 25653 29561 25656
rect 29595 25684 29607 25687
rect 30116 25684 30144 25712
rect 29595 25656 30144 25684
rect 29595 25653 29607 25656
rect 29549 25647 29607 25653
rect 2760 25594 32200 25616
rect 2760 25542 6946 25594
rect 6998 25542 7010 25594
rect 7062 25542 7074 25594
rect 7126 25542 7138 25594
rect 7190 25542 7202 25594
rect 7254 25542 14306 25594
rect 14358 25542 14370 25594
rect 14422 25542 14434 25594
rect 14486 25542 14498 25594
rect 14550 25542 14562 25594
rect 14614 25542 21666 25594
rect 21718 25542 21730 25594
rect 21782 25542 21794 25594
rect 21846 25542 21858 25594
rect 21910 25542 21922 25594
rect 21974 25542 29026 25594
rect 29078 25542 29090 25594
rect 29142 25542 29154 25594
rect 29206 25542 29218 25594
rect 29270 25542 29282 25594
rect 29334 25542 32200 25594
rect 2760 25520 32200 25542
rect 4709 25483 4767 25489
rect 4709 25449 4721 25483
rect 4755 25480 4767 25483
rect 4982 25480 4988 25492
rect 4755 25452 4988 25480
rect 4755 25449 4767 25452
rect 4709 25443 4767 25449
rect 4982 25440 4988 25452
rect 5040 25440 5046 25492
rect 5077 25483 5135 25489
rect 5077 25449 5089 25483
rect 5123 25480 5135 25483
rect 5166 25480 5172 25492
rect 5123 25452 5172 25480
rect 5123 25449 5135 25452
rect 5077 25443 5135 25449
rect 5166 25440 5172 25452
rect 5224 25440 5230 25492
rect 5258 25440 5264 25492
rect 5316 25480 5322 25492
rect 6273 25483 6331 25489
rect 6273 25480 6285 25483
rect 5316 25452 6285 25480
rect 5316 25440 5322 25452
rect 6273 25449 6285 25452
rect 6319 25449 6331 25483
rect 6273 25443 6331 25449
rect 7101 25483 7159 25489
rect 7101 25449 7113 25483
rect 7147 25480 7159 25483
rect 7147 25452 7696 25480
rect 7147 25449 7159 25452
rect 7101 25443 7159 25449
rect 5810 25412 5816 25424
rect 5184 25384 5816 25412
rect 5184 25353 5212 25384
rect 5810 25372 5816 25384
rect 5868 25372 5874 25424
rect 5905 25415 5963 25421
rect 5905 25381 5917 25415
rect 5951 25412 5963 25415
rect 6178 25412 6184 25424
rect 5951 25384 6184 25412
rect 5951 25381 5963 25384
rect 5905 25375 5963 25381
rect 6178 25372 6184 25384
rect 6236 25412 6242 25424
rect 7668 25412 7696 25452
rect 7742 25440 7748 25492
rect 7800 25440 7806 25492
rect 8021 25483 8079 25489
rect 8021 25449 8033 25483
rect 8067 25480 8079 25483
rect 8202 25480 8208 25492
rect 8067 25452 8208 25480
rect 8067 25449 8079 25452
rect 8021 25443 8079 25449
rect 8202 25440 8208 25452
rect 8260 25440 8266 25492
rect 8389 25483 8447 25489
rect 8389 25449 8401 25483
rect 8435 25480 8447 25483
rect 9306 25480 9312 25492
rect 8435 25452 9312 25480
rect 8435 25449 8447 25452
rect 8389 25443 8447 25449
rect 9306 25440 9312 25452
rect 9364 25440 9370 25492
rect 10597 25483 10655 25489
rect 10597 25449 10609 25483
rect 10643 25480 10655 25483
rect 10962 25480 10968 25492
rect 10643 25452 10968 25480
rect 10643 25449 10655 25452
rect 10597 25443 10655 25449
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 11606 25480 11612 25492
rect 11072 25452 11612 25480
rect 11072 25412 11100 25452
rect 11606 25440 11612 25452
rect 11664 25440 11670 25492
rect 11882 25440 11888 25492
rect 11940 25440 11946 25492
rect 12802 25440 12808 25492
rect 12860 25480 12866 25492
rect 12989 25483 13047 25489
rect 12989 25480 13001 25483
rect 12860 25452 13001 25480
rect 12860 25440 12866 25452
rect 12989 25449 13001 25452
rect 13035 25449 13047 25483
rect 12989 25443 13047 25449
rect 13170 25440 13176 25492
rect 13228 25480 13234 25492
rect 13449 25483 13507 25489
rect 13449 25480 13461 25483
rect 13228 25452 13461 25480
rect 13228 25440 13234 25452
rect 13449 25449 13461 25452
rect 13495 25449 13507 25483
rect 13449 25443 13507 25449
rect 13817 25483 13875 25489
rect 13817 25449 13829 25483
rect 13863 25480 13875 25483
rect 14734 25480 14740 25492
rect 13863 25452 14740 25480
rect 13863 25449 13875 25452
rect 13817 25443 13875 25449
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 15470 25480 15476 25492
rect 15212 25452 15476 25480
rect 11422 25412 11428 25424
rect 6236 25384 7512 25412
rect 6236 25372 6242 25384
rect 7484 25356 7512 25384
rect 7668 25384 11100 25412
rect 11164 25384 11428 25412
rect 5169 25347 5227 25353
rect 5169 25313 5181 25347
rect 5215 25313 5227 25347
rect 5169 25307 5227 25313
rect 5721 25347 5779 25353
rect 5721 25313 5733 25347
rect 5767 25313 5779 25347
rect 5721 25307 5779 25313
rect 6089 25347 6147 25353
rect 6089 25313 6101 25347
rect 6135 25313 6147 25347
rect 6089 25307 6147 25313
rect 3418 25236 3424 25288
rect 3476 25236 3482 25288
rect 5353 25279 5411 25285
rect 5353 25245 5365 25279
rect 5399 25245 5411 25279
rect 5353 25239 5411 25245
rect 5368 25208 5396 25239
rect 5368 25180 5672 25208
rect 5644 25152 5672 25180
rect 4065 25143 4123 25149
rect 4065 25109 4077 25143
rect 4111 25140 4123 25143
rect 4522 25140 4528 25152
rect 4111 25112 4528 25140
rect 4111 25109 4123 25112
rect 4065 25103 4123 25109
rect 4522 25100 4528 25112
rect 4580 25100 4586 25152
rect 5534 25100 5540 25152
rect 5592 25100 5598 25152
rect 5626 25100 5632 25152
rect 5684 25100 5690 25152
rect 5736 25140 5764 25307
rect 5902 25236 5908 25288
rect 5960 25236 5966 25288
rect 6104 25276 6132 25307
rect 6270 25304 6276 25356
rect 6328 25344 6334 25356
rect 6365 25347 6423 25353
rect 6365 25344 6377 25347
rect 6328 25316 6377 25344
rect 6328 25304 6334 25316
rect 6365 25313 6377 25316
rect 6411 25344 6423 25347
rect 7282 25344 7288 25356
rect 6411 25316 7288 25344
rect 6411 25313 6423 25316
rect 6365 25307 6423 25313
rect 7282 25304 7288 25316
rect 7340 25304 7346 25356
rect 7466 25304 7472 25356
rect 7524 25304 7530 25356
rect 7668 25276 7696 25384
rect 7834 25304 7840 25356
rect 7892 25304 7898 25356
rect 8481 25347 8539 25353
rect 8481 25313 8493 25347
rect 8527 25344 8539 25347
rect 9674 25344 9680 25356
rect 8527 25316 9680 25344
rect 8527 25313 8539 25316
rect 8481 25307 8539 25313
rect 9674 25304 9680 25316
rect 9732 25344 9738 25356
rect 9953 25347 10011 25353
rect 9953 25344 9965 25347
rect 9732 25316 9965 25344
rect 9732 25304 9738 25316
rect 9953 25313 9965 25316
rect 9999 25313 10011 25347
rect 9953 25307 10011 25313
rect 10042 25304 10048 25356
rect 10100 25344 10106 25356
rect 10229 25347 10287 25353
rect 10229 25344 10241 25347
rect 10100 25316 10241 25344
rect 10100 25304 10106 25316
rect 10229 25313 10241 25316
rect 10275 25313 10287 25347
rect 10229 25307 10287 25313
rect 10318 25304 10324 25356
rect 10376 25304 10382 25356
rect 10505 25347 10563 25353
rect 10505 25313 10517 25347
rect 10551 25344 10563 25347
rect 10778 25344 10784 25356
rect 10551 25316 10784 25344
rect 10551 25313 10563 25316
rect 10505 25307 10563 25313
rect 10778 25304 10784 25316
rect 10836 25304 10842 25356
rect 11164 25353 11192 25384
rect 11422 25372 11428 25384
rect 11480 25372 11486 25424
rect 11517 25415 11575 25421
rect 11517 25381 11529 25415
rect 11563 25412 11575 25415
rect 11900 25412 11928 25440
rect 13265 25415 13323 25421
rect 13265 25412 13277 25415
rect 11563 25384 11928 25412
rect 12742 25384 13277 25412
rect 11563 25381 11575 25384
rect 11517 25375 11575 25381
rect 13265 25381 13277 25384
rect 13311 25381 13323 25415
rect 13538 25412 13544 25424
rect 13265 25375 13323 25381
rect 13372 25384 13544 25412
rect 13372 25353 13400 25384
rect 13538 25372 13544 25384
rect 13596 25412 13602 25424
rect 15212 25421 15240 25452
rect 15470 25440 15476 25452
rect 15528 25440 15534 25492
rect 16669 25483 16727 25489
rect 16669 25449 16681 25483
rect 16715 25480 16727 25483
rect 17034 25480 17040 25492
rect 16715 25452 17040 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 20530 25480 20536 25492
rect 18708 25452 20536 25480
rect 15197 25415 15255 25421
rect 13596 25384 14780 25412
rect 13596 25372 13602 25384
rect 14752 25356 14780 25384
rect 15197 25381 15209 25415
rect 15243 25381 15255 25415
rect 15197 25375 15255 25381
rect 15930 25372 15936 25424
rect 15988 25372 15994 25424
rect 16758 25372 16764 25424
rect 16816 25412 16822 25424
rect 16945 25415 17003 25421
rect 16945 25412 16957 25415
rect 16816 25384 16957 25412
rect 16816 25372 16822 25384
rect 16945 25381 16957 25384
rect 16991 25381 17003 25415
rect 16945 25375 17003 25381
rect 11149 25347 11207 25353
rect 11149 25313 11161 25347
rect 11195 25313 11207 25347
rect 11149 25307 11207 25313
rect 13357 25347 13415 25353
rect 13357 25313 13369 25347
rect 13403 25313 13415 25347
rect 13357 25307 13415 25313
rect 13446 25304 13452 25356
rect 13504 25304 13510 25356
rect 13909 25347 13967 25353
rect 13909 25313 13921 25347
rect 13955 25344 13967 25347
rect 14277 25347 14335 25353
rect 13955 25316 14136 25344
rect 13955 25313 13967 25316
rect 13909 25307 13967 25313
rect 6104 25248 7696 25276
rect 8573 25279 8631 25285
rect 8573 25245 8585 25279
rect 8619 25245 8631 25279
rect 8573 25239 8631 25245
rect 5920 25208 5948 25236
rect 8110 25208 8116 25220
rect 5920 25180 8116 25208
rect 8110 25168 8116 25180
rect 8168 25208 8174 25220
rect 8588 25208 8616 25239
rect 9306 25236 9312 25288
rect 9364 25236 9370 25288
rect 10873 25279 10931 25285
rect 10873 25245 10885 25279
rect 10919 25276 10931 25279
rect 11054 25276 11060 25288
rect 10919 25248 11060 25276
rect 10919 25245 10931 25248
rect 10873 25239 10931 25245
rect 11054 25236 11060 25248
rect 11112 25236 11118 25288
rect 11241 25279 11299 25285
rect 11241 25276 11253 25279
rect 11164 25248 11253 25276
rect 11164 25220 11192 25248
rect 11241 25245 11253 25248
rect 11287 25245 11299 25279
rect 11241 25239 11299 25245
rect 11514 25236 11520 25288
rect 11572 25276 11578 25288
rect 13464 25276 13492 25304
rect 14108 25288 14136 25316
rect 14277 25313 14289 25347
rect 14323 25313 14335 25347
rect 14277 25307 14335 25313
rect 14001 25279 14059 25285
rect 14001 25276 14013 25279
rect 11572 25248 13400 25276
rect 13464 25248 14013 25276
rect 11572 25236 11578 25248
rect 9033 25211 9091 25217
rect 9033 25208 9045 25211
rect 8168 25180 9045 25208
rect 8168 25168 8174 25180
rect 9033 25177 9045 25180
rect 9079 25177 9091 25211
rect 9033 25171 9091 25177
rect 10336 25180 11100 25208
rect 6733 25143 6791 25149
rect 6733 25140 6745 25143
rect 5736 25112 6745 25140
rect 6733 25109 6745 25112
rect 6779 25140 6791 25143
rect 9582 25140 9588 25152
rect 6779 25112 9588 25140
rect 6779 25109 6791 25112
rect 6733 25103 6791 25109
rect 9582 25100 9588 25112
rect 9640 25100 9646 25152
rect 10134 25100 10140 25152
rect 10192 25100 10198 25152
rect 10336 25149 10364 25180
rect 10321 25143 10379 25149
rect 10321 25109 10333 25143
rect 10367 25109 10379 25143
rect 10321 25103 10379 25109
rect 10870 25100 10876 25152
rect 10928 25100 10934 25152
rect 11072 25140 11100 25180
rect 11146 25168 11152 25220
rect 11204 25168 11210 25220
rect 13372 25208 13400 25248
rect 14001 25245 14013 25248
rect 14047 25245 14059 25279
rect 14001 25239 14059 25245
rect 14090 25236 14096 25288
rect 14148 25236 14154 25288
rect 14292 25208 14320 25307
rect 14734 25304 14740 25356
rect 14792 25304 14798 25356
rect 17586 25304 17592 25356
rect 17644 25344 17650 25356
rect 18708 25353 18736 25452
rect 20530 25440 20536 25452
rect 20588 25440 20594 25492
rect 22370 25440 22376 25492
rect 22428 25480 22434 25492
rect 22649 25483 22707 25489
rect 22649 25480 22661 25483
rect 22428 25452 22661 25480
rect 22428 25440 22434 25452
rect 22649 25449 22661 25452
rect 22695 25449 22707 25483
rect 22649 25443 22707 25449
rect 23842 25440 23848 25492
rect 23900 25440 23906 25492
rect 24857 25483 24915 25489
rect 24857 25480 24869 25483
rect 24780 25452 24869 25480
rect 21453 25415 21511 25421
rect 21453 25412 21465 25415
rect 20194 25384 21465 25412
rect 21453 25381 21465 25384
rect 21499 25381 21511 25415
rect 21453 25375 21511 25381
rect 22462 25372 22468 25424
rect 22520 25372 22526 25424
rect 23860 25412 23888 25440
rect 23584 25384 23796 25412
rect 23860 25384 24256 25412
rect 17773 25347 17831 25353
rect 17773 25344 17785 25347
rect 17644 25316 17785 25344
rect 17644 25304 17650 25316
rect 17773 25313 17785 25316
rect 17819 25344 17831 25347
rect 18693 25347 18751 25353
rect 17819 25316 18552 25344
rect 17819 25313 17831 25316
rect 17773 25307 17831 25313
rect 14458 25236 14464 25288
rect 14516 25276 14522 25288
rect 14553 25279 14611 25285
rect 14553 25276 14565 25279
rect 14516 25248 14565 25276
rect 14516 25236 14522 25248
rect 14553 25245 14565 25248
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 14642 25236 14648 25288
rect 14700 25276 14706 25288
rect 14921 25279 14979 25285
rect 14921 25276 14933 25279
rect 14700 25248 14933 25276
rect 14700 25236 14706 25248
rect 14921 25245 14933 25248
rect 14967 25245 14979 25279
rect 18414 25276 18420 25288
rect 14921 25239 14979 25245
rect 15028 25248 18420 25276
rect 15028 25208 15056 25248
rect 18414 25236 18420 25248
rect 18472 25236 18478 25288
rect 13372 25180 15056 25208
rect 13998 25140 14004 25152
rect 11072 25112 14004 25140
rect 13998 25100 14004 25112
rect 14056 25100 14062 25152
rect 14550 25100 14556 25152
rect 14608 25100 14614 25152
rect 14829 25143 14887 25149
rect 14829 25109 14841 25143
rect 14875 25140 14887 25143
rect 15378 25140 15384 25152
rect 14875 25112 15384 25140
rect 14875 25109 14887 25112
rect 14829 25103 14887 25109
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 18141 25143 18199 25149
rect 18141 25109 18153 25143
rect 18187 25140 18199 25143
rect 18322 25140 18328 25152
rect 18187 25112 18328 25140
rect 18187 25109 18199 25112
rect 18141 25103 18199 25109
rect 18322 25100 18328 25112
rect 18380 25140 18386 25152
rect 18524 25140 18552 25316
rect 18693 25313 18705 25347
rect 18739 25313 18751 25347
rect 18693 25307 18751 25313
rect 21545 25347 21603 25353
rect 21545 25313 21557 25347
rect 21591 25344 21603 25347
rect 22002 25344 22008 25356
rect 21591 25316 22008 25344
rect 21591 25313 21603 25316
rect 21545 25307 21603 25313
rect 22002 25304 22008 25316
rect 22060 25344 22066 25356
rect 22373 25347 22431 25353
rect 22373 25344 22385 25347
rect 22060 25316 22385 25344
rect 22060 25304 22066 25316
rect 22373 25313 22385 25316
rect 22419 25313 22431 25347
rect 22373 25307 22431 25313
rect 18969 25279 19027 25285
rect 18969 25245 18981 25279
rect 19015 25276 19027 25279
rect 19518 25276 19524 25288
rect 19015 25248 19524 25276
rect 19015 25245 19027 25248
rect 18969 25239 19027 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 21269 25279 21327 25285
rect 21269 25245 21281 25279
rect 21315 25245 21327 25279
rect 22388 25276 22416 25307
rect 22738 25276 22744 25288
rect 22388 25248 22744 25276
rect 21269 25239 21327 25245
rect 20441 25211 20499 25217
rect 20441 25177 20453 25211
rect 20487 25208 20499 25211
rect 21284 25208 21312 25239
rect 22738 25236 22744 25248
rect 22796 25236 22802 25288
rect 23293 25279 23351 25285
rect 23293 25245 23305 25279
rect 23339 25276 23351 25279
rect 23477 25279 23535 25285
rect 23477 25276 23489 25279
rect 23339 25248 23489 25276
rect 23339 25245 23351 25248
rect 23293 25239 23351 25245
rect 23477 25245 23489 25248
rect 23523 25245 23535 25279
rect 23477 25239 23535 25245
rect 23584 25208 23612 25384
rect 23661 25347 23719 25353
rect 23661 25313 23673 25347
rect 23707 25313 23719 25347
rect 23661 25307 23719 25313
rect 20487 25180 23612 25208
rect 20487 25177 20499 25180
rect 20441 25171 20499 25177
rect 19058 25140 19064 25152
rect 18380 25112 19064 25140
rect 18380 25100 18386 25112
rect 19058 25100 19064 25112
rect 19116 25100 19122 25152
rect 20622 25100 20628 25152
rect 20680 25100 20686 25152
rect 23676 25140 23704 25307
rect 23768 25208 23796 25384
rect 23934 25304 23940 25356
rect 23992 25304 23998 25356
rect 24228 25353 24256 25384
rect 24121 25347 24179 25353
rect 24121 25313 24133 25347
rect 24167 25313 24179 25347
rect 24121 25307 24179 25313
rect 24213 25347 24271 25353
rect 24213 25313 24225 25347
rect 24259 25313 24271 25347
rect 24213 25307 24271 25313
rect 24136 25276 24164 25307
rect 24780 25276 24808 25452
rect 24857 25449 24869 25452
rect 24903 25449 24915 25483
rect 24857 25443 24915 25449
rect 24949 25483 25007 25489
rect 24949 25449 24961 25483
rect 24995 25480 25007 25483
rect 25314 25480 25320 25492
rect 24995 25452 25320 25480
rect 24995 25449 25007 25452
rect 24949 25443 25007 25449
rect 25314 25440 25320 25452
rect 25372 25440 25378 25492
rect 25590 25440 25596 25492
rect 25648 25440 25654 25492
rect 25682 25440 25688 25492
rect 25740 25440 25746 25492
rect 25958 25440 25964 25492
rect 26016 25480 26022 25492
rect 26605 25483 26663 25489
rect 26605 25480 26617 25483
rect 26016 25452 26617 25480
rect 26016 25440 26022 25452
rect 26605 25449 26617 25452
rect 26651 25480 26663 25483
rect 26694 25480 26700 25492
rect 26651 25452 26700 25480
rect 26651 25449 26663 25452
rect 26605 25443 26663 25449
rect 26694 25440 26700 25452
rect 26752 25440 26758 25492
rect 27890 25440 27896 25492
rect 27948 25480 27954 25492
rect 30742 25480 30748 25492
rect 27948 25452 30748 25480
rect 27948 25440 27954 25452
rect 30742 25440 30748 25452
rect 30800 25480 30806 25492
rect 31386 25480 31392 25492
rect 30800 25452 31392 25480
rect 30800 25440 30806 25452
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 25608 25412 25636 25440
rect 25424 25384 25636 25412
rect 25700 25384 30512 25412
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 25133 25347 25191 25353
rect 25133 25344 25145 25347
rect 24912 25316 25145 25344
rect 24912 25304 24918 25316
rect 25133 25313 25145 25316
rect 25179 25313 25191 25347
rect 25133 25307 25191 25313
rect 25222 25304 25228 25356
rect 25280 25304 25286 25356
rect 25424 25353 25452 25384
rect 25409 25347 25467 25353
rect 25409 25313 25421 25347
rect 25455 25313 25467 25347
rect 25409 25307 25467 25313
rect 25498 25304 25504 25356
rect 25556 25344 25562 25356
rect 25593 25347 25651 25353
rect 25593 25344 25605 25347
rect 25556 25316 25605 25344
rect 25556 25304 25562 25316
rect 25593 25313 25605 25316
rect 25639 25313 25651 25347
rect 25593 25307 25651 25313
rect 24946 25276 24952 25288
rect 24136 25248 24952 25276
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25700 25276 25728 25384
rect 26050 25304 26056 25356
rect 26108 25304 26114 25356
rect 28445 25347 28503 25353
rect 28445 25313 28457 25347
rect 28491 25344 28503 25347
rect 29362 25344 29368 25356
rect 28491 25316 29368 25344
rect 28491 25313 28503 25316
rect 28445 25307 28503 25313
rect 29362 25304 29368 25316
rect 29420 25304 29426 25356
rect 29641 25347 29699 25353
rect 29641 25313 29653 25347
rect 29687 25344 29699 25347
rect 29730 25344 29736 25356
rect 29687 25316 29736 25344
rect 29687 25313 29699 25316
rect 29641 25307 29699 25313
rect 29730 25304 29736 25316
rect 29788 25304 29794 25356
rect 30484 25353 30512 25384
rect 30469 25347 30527 25353
rect 30469 25313 30481 25347
rect 30515 25313 30527 25347
rect 30469 25307 30527 25313
rect 25240 25248 25728 25276
rect 25240 25208 25268 25248
rect 26326 25236 26332 25288
rect 26384 25276 26390 25288
rect 31294 25276 31300 25288
rect 26384 25248 31300 25276
rect 26384 25236 26390 25248
rect 31294 25236 31300 25248
rect 31352 25236 31358 25288
rect 31665 25279 31723 25285
rect 31665 25245 31677 25279
rect 31711 25276 31723 25279
rect 33134 25276 33140 25288
rect 31711 25248 33140 25276
rect 31711 25245 31723 25248
rect 31665 25239 31723 25245
rect 33134 25236 33140 25248
rect 33192 25236 33198 25288
rect 23768 25180 25268 25208
rect 25317 25211 25375 25217
rect 25317 25177 25329 25211
rect 25363 25208 25375 25211
rect 25406 25208 25412 25220
rect 25363 25180 25412 25208
rect 25363 25177 25375 25180
rect 25317 25171 25375 25177
rect 25332 25140 25360 25171
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 28166 25168 28172 25220
rect 28224 25168 28230 25220
rect 23676 25112 25360 25140
rect 27982 25100 27988 25152
rect 28040 25100 28046 25152
rect 28997 25143 29055 25149
rect 28997 25109 29009 25143
rect 29043 25140 29055 25143
rect 29178 25140 29184 25152
rect 29043 25112 29184 25140
rect 29043 25109 29055 25112
rect 28997 25103 29055 25109
rect 29178 25100 29184 25112
rect 29236 25140 29242 25152
rect 30374 25140 30380 25152
rect 29236 25112 30380 25140
rect 29236 25100 29242 25112
rect 30374 25100 30380 25112
rect 30432 25100 30438 25152
rect 2760 25050 32200 25072
rect 2760 24998 6286 25050
rect 6338 24998 6350 25050
rect 6402 24998 6414 25050
rect 6466 24998 6478 25050
rect 6530 24998 6542 25050
rect 6594 24998 13646 25050
rect 13698 24998 13710 25050
rect 13762 24998 13774 25050
rect 13826 24998 13838 25050
rect 13890 24998 13902 25050
rect 13954 24998 21006 25050
rect 21058 24998 21070 25050
rect 21122 24998 21134 25050
rect 21186 24998 21198 25050
rect 21250 24998 21262 25050
rect 21314 24998 28366 25050
rect 28418 24998 28430 25050
rect 28482 24998 28494 25050
rect 28546 24998 28558 25050
rect 28610 24998 28622 25050
rect 28674 24998 32200 25050
rect 2760 24976 32200 24998
rect 5810 24896 5816 24948
rect 5868 24936 5874 24948
rect 5905 24939 5963 24945
rect 5905 24936 5917 24939
rect 5868 24908 5917 24936
rect 5868 24896 5874 24908
rect 5905 24905 5917 24908
rect 5951 24905 5963 24939
rect 5905 24899 5963 24905
rect 7824 24939 7882 24945
rect 7824 24905 7836 24939
rect 7870 24936 7882 24939
rect 8570 24936 8576 24948
rect 7870 24908 8576 24936
rect 7870 24905 7882 24908
rect 7824 24899 7882 24905
rect 8570 24896 8576 24908
rect 8628 24896 8634 24948
rect 9306 24896 9312 24948
rect 9364 24896 9370 24948
rect 9398 24896 9404 24948
rect 9456 24896 9462 24948
rect 10042 24896 10048 24948
rect 10100 24896 10106 24948
rect 10870 24896 10876 24948
rect 10928 24936 10934 24948
rect 11698 24936 11704 24948
rect 10928 24908 11704 24936
rect 10928 24896 10934 24908
rect 11698 24896 11704 24908
rect 11756 24896 11762 24948
rect 14274 24936 14280 24948
rect 12544 24908 14280 24936
rect 10060 24868 10088 24896
rect 10321 24871 10379 24877
rect 10060 24840 10272 24868
rect 1302 24760 1308 24812
rect 1360 24800 1366 24812
rect 3513 24803 3571 24809
rect 3513 24800 3525 24803
rect 1360 24772 3525 24800
rect 1360 24760 1366 24772
rect 3513 24769 3525 24772
rect 3559 24769 3571 24803
rect 3513 24763 3571 24769
rect 4246 24760 4252 24812
rect 4304 24800 4310 24812
rect 7374 24800 7380 24812
rect 4304 24772 7380 24800
rect 4304 24760 4310 24772
rect 7374 24760 7380 24772
rect 7432 24800 7438 24812
rect 7561 24803 7619 24809
rect 7561 24800 7573 24803
rect 7432 24772 7573 24800
rect 7432 24760 7438 24772
rect 7561 24769 7573 24772
rect 7607 24769 7619 24803
rect 7561 24763 7619 24769
rect 8956 24772 10180 24800
rect 3234 24692 3240 24744
rect 3292 24692 3298 24744
rect 5261 24735 5319 24741
rect 5261 24701 5273 24735
rect 5307 24732 5319 24735
rect 5534 24732 5540 24744
rect 5307 24704 5540 24732
rect 5307 24701 5319 24704
rect 5261 24695 5319 24701
rect 5534 24692 5540 24704
rect 5592 24692 5598 24744
rect 5813 24735 5871 24741
rect 5813 24701 5825 24735
rect 5859 24732 5871 24735
rect 6178 24732 6184 24744
rect 5859 24704 6184 24732
rect 5859 24701 5871 24704
rect 5813 24695 5871 24701
rect 6178 24692 6184 24704
rect 6236 24692 6242 24744
rect 6454 24692 6460 24744
rect 6512 24692 6518 24744
rect 7282 24692 7288 24744
rect 7340 24692 7346 24744
rect 8956 24718 8984 24772
rect 10152 24744 10180 24772
rect 9582 24692 9588 24744
rect 9640 24692 9646 24744
rect 9674 24692 9680 24744
rect 9732 24692 9738 24744
rect 9950 24692 9956 24744
rect 10008 24692 10014 24744
rect 10134 24692 10140 24744
rect 10192 24692 10198 24744
rect 10244 24741 10272 24840
rect 10321 24837 10333 24871
rect 10367 24868 10379 24871
rect 10686 24868 10692 24880
rect 10367 24840 10692 24868
rect 10367 24837 10379 24840
rect 10321 24831 10379 24837
rect 10686 24828 10692 24840
rect 10744 24828 10750 24880
rect 10778 24828 10784 24880
rect 10836 24868 10842 24880
rect 11882 24868 11888 24880
rect 10836 24840 11888 24868
rect 10836 24828 10842 24840
rect 11882 24828 11888 24840
rect 11940 24828 11946 24880
rect 11977 24803 12035 24809
rect 11977 24800 11989 24803
rect 10336 24772 11989 24800
rect 10229 24735 10287 24741
rect 10229 24701 10241 24735
rect 10275 24701 10287 24735
rect 10229 24695 10287 24701
rect 3878 24624 3884 24676
rect 3936 24664 3942 24676
rect 3936 24636 6684 24664
rect 3936 24624 3942 24636
rect 4614 24556 4620 24608
rect 4672 24556 4678 24608
rect 5258 24556 5264 24608
rect 5316 24596 5322 24608
rect 5442 24596 5448 24608
rect 5316 24568 5448 24596
rect 5316 24556 5322 24568
rect 5442 24556 5448 24568
rect 5500 24556 5506 24608
rect 5626 24556 5632 24608
rect 5684 24596 5690 24608
rect 6656 24605 6684 24636
rect 9122 24624 9128 24676
rect 9180 24664 9186 24676
rect 9769 24667 9827 24673
rect 9769 24664 9781 24667
rect 9180 24636 9781 24664
rect 9180 24624 9186 24636
rect 9769 24633 9781 24636
rect 9815 24664 9827 24667
rect 10336 24664 10364 24772
rect 11977 24769 11989 24772
rect 12023 24769 12035 24803
rect 12544 24800 12572 24908
rect 14274 24896 14280 24908
rect 14332 24896 14338 24948
rect 14550 24896 14556 24948
rect 14608 24936 14614 24948
rect 14918 24936 14924 24948
rect 14608 24908 14924 24936
rect 14608 24896 14614 24908
rect 14918 24896 14924 24908
rect 14976 24896 14982 24948
rect 15562 24896 15568 24948
rect 15620 24896 15626 24948
rect 15749 24939 15807 24945
rect 15749 24905 15761 24939
rect 15795 24936 15807 24939
rect 16298 24936 16304 24948
rect 15795 24908 16304 24936
rect 15795 24905 15807 24908
rect 15749 24899 15807 24905
rect 16298 24896 16304 24908
rect 16356 24896 16362 24948
rect 18506 24936 18512 24948
rect 16546 24908 18512 24936
rect 14458 24868 14464 24880
rect 13924 24840 14464 24868
rect 11977 24763 12035 24769
rect 12084 24772 12572 24800
rect 12621 24803 12679 24809
rect 10778 24692 10784 24744
rect 10836 24692 10842 24744
rect 10962 24692 10968 24744
rect 11020 24692 11026 24744
rect 11149 24735 11207 24741
rect 11149 24701 11161 24735
rect 11195 24732 11207 24735
rect 11422 24732 11428 24744
rect 11195 24704 11428 24732
rect 11195 24701 11207 24704
rect 11149 24695 11207 24701
rect 11422 24692 11428 24704
rect 11480 24692 11486 24744
rect 11514 24692 11520 24744
rect 11572 24692 11578 24744
rect 11793 24735 11851 24741
rect 11793 24701 11805 24735
rect 11839 24701 11851 24735
rect 11793 24695 11851 24701
rect 10873 24667 10931 24673
rect 10873 24664 10885 24667
rect 9815 24636 10364 24664
rect 10428 24636 10885 24664
rect 9815 24633 9827 24636
rect 9769 24627 9827 24633
rect 5721 24599 5779 24605
rect 5721 24596 5733 24599
rect 5684 24568 5733 24596
rect 5684 24556 5690 24568
rect 5721 24565 5733 24568
rect 5767 24565 5779 24599
rect 5721 24559 5779 24565
rect 6641 24599 6699 24605
rect 6641 24565 6653 24599
rect 6687 24596 6699 24599
rect 10428 24596 10456 24636
rect 10873 24633 10885 24636
rect 10919 24633 10931 24667
rect 10873 24627 10931 24633
rect 11054 24624 11060 24676
rect 11112 24664 11118 24676
rect 11532 24664 11560 24692
rect 11112 24636 11560 24664
rect 11112 24624 11118 24636
rect 11808 24608 11836 24695
rect 11882 24692 11888 24744
rect 11940 24692 11946 24744
rect 12084 24741 12112 24772
rect 12621 24769 12633 24803
rect 12667 24800 12679 24803
rect 13262 24800 13268 24812
rect 12667 24772 13268 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 13262 24760 13268 24772
rect 13320 24760 13326 24812
rect 13924 24744 13952 24840
rect 14458 24828 14464 24840
rect 14516 24868 14522 24880
rect 15102 24868 15108 24880
rect 14516 24840 15108 24868
rect 14516 24828 14522 24840
rect 15102 24828 15108 24840
rect 15160 24828 15166 24880
rect 14090 24760 14096 24812
rect 14148 24760 14154 24812
rect 14369 24803 14427 24809
rect 14369 24769 14381 24803
rect 14415 24800 14427 24803
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 14415 24772 15025 24800
rect 14415 24769 14427 24772
rect 14369 24763 14427 24769
rect 15013 24769 15025 24772
rect 15059 24769 15071 24803
rect 15580 24800 15608 24896
rect 16546 24868 16574 24908
rect 18506 24896 18512 24908
rect 18564 24936 18570 24948
rect 18564 24908 19012 24936
rect 18564 24896 18570 24908
rect 18984 24880 19012 24908
rect 19518 24896 19524 24948
rect 19576 24896 19582 24948
rect 27890 24936 27896 24948
rect 19628 24908 27896 24936
rect 16316 24840 16574 24868
rect 16316 24809 16344 24840
rect 18966 24828 18972 24880
rect 19024 24828 19030 24880
rect 19058 24828 19064 24880
rect 19116 24868 19122 24880
rect 19628 24868 19656 24908
rect 27890 24896 27896 24908
rect 27948 24896 27954 24948
rect 27982 24896 27988 24948
rect 28040 24896 28046 24948
rect 28166 24896 28172 24948
rect 28224 24896 28230 24948
rect 29730 24896 29736 24948
rect 29788 24936 29794 24948
rect 30009 24939 30067 24945
rect 30009 24936 30021 24939
rect 29788 24908 30021 24936
rect 29788 24896 29794 24908
rect 30009 24905 30021 24908
rect 30055 24905 30067 24939
rect 30009 24899 30067 24905
rect 19116 24840 19656 24868
rect 19116 24828 19122 24840
rect 23474 24828 23480 24880
rect 23532 24828 23538 24880
rect 25498 24828 25504 24880
rect 25556 24828 25562 24880
rect 28000 24868 28028 24896
rect 28000 24840 28396 24868
rect 16301 24803 16359 24809
rect 16301 24800 16313 24803
rect 15580 24772 16313 24800
rect 15013 24763 15071 24769
rect 16301 24769 16313 24772
rect 16347 24769 16359 24803
rect 16301 24763 16359 24769
rect 17126 24760 17132 24812
rect 17184 24800 17190 24812
rect 17681 24803 17739 24809
rect 17681 24800 17693 24803
rect 17184 24772 17693 24800
rect 17184 24760 17190 24772
rect 17681 24769 17693 24772
rect 17727 24769 17739 24803
rect 17681 24763 17739 24769
rect 19610 24760 19616 24812
rect 19668 24800 19674 24812
rect 19981 24803 20039 24809
rect 19981 24800 19993 24803
rect 19668 24772 19993 24800
rect 19668 24760 19674 24772
rect 19981 24769 19993 24772
rect 20027 24769 20039 24803
rect 19981 24763 20039 24769
rect 20070 24760 20076 24812
rect 20128 24760 20134 24812
rect 23293 24803 23351 24809
rect 23293 24769 23305 24803
rect 23339 24800 23351 24803
rect 23492 24800 23520 24828
rect 23339 24772 23520 24800
rect 23339 24769 23351 24772
rect 23293 24763 23351 24769
rect 12069 24735 12127 24741
rect 12069 24701 12081 24735
rect 12115 24701 12127 24735
rect 12345 24735 12403 24741
rect 12345 24732 12357 24735
rect 12069 24695 12127 24701
rect 12176 24704 12357 24732
rect 11900 24664 11928 24692
rect 12176 24664 12204 24704
rect 12345 24701 12357 24704
rect 12391 24701 12403 24735
rect 12345 24695 12403 24701
rect 12529 24735 12587 24741
rect 12529 24701 12541 24735
rect 12575 24701 12587 24735
rect 12529 24695 12587 24701
rect 11900 24636 12204 24664
rect 12250 24624 12256 24676
rect 12308 24624 12314 24676
rect 6687 24568 10456 24596
rect 6687 24565 6699 24568
rect 6641 24559 6699 24565
rect 10594 24556 10600 24608
rect 10652 24556 10658 24608
rect 11238 24556 11244 24608
rect 11296 24556 11302 24608
rect 11790 24556 11796 24608
rect 11848 24556 11854 24608
rect 12268 24596 12296 24624
rect 12437 24599 12495 24605
rect 12437 24596 12449 24599
rect 12268 24568 12449 24596
rect 12437 24565 12449 24568
rect 12483 24565 12495 24599
rect 12544 24596 12572 24695
rect 13906 24692 13912 24744
rect 13964 24692 13970 24744
rect 13998 24692 14004 24744
rect 14056 24692 14062 24744
rect 14108 24732 14136 24760
rect 14461 24735 14519 24741
rect 14461 24732 14473 24735
rect 14108 24704 14473 24732
rect 14461 24701 14473 24704
rect 14507 24701 14519 24735
rect 14461 24695 14519 24701
rect 16117 24735 16175 24741
rect 16117 24701 16129 24735
rect 16163 24732 16175 24735
rect 16482 24732 16488 24744
rect 16163 24704 16488 24732
rect 16163 24701 16175 24704
rect 16117 24695 16175 24701
rect 16482 24692 16488 24704
rect 16540 24692 16546 24744
rect 19058 24692 19064 24744
rect 19116 24692 19122 24744
rect 19889 24735 19947 24741
rect 19889 24701 19901 24735
rect 19935 24732 19947 24735
rect 20622 24732 20628 24744
rect 19935 24704 20628 24732
rect 19935 24701 19947 24704
rect 19889 24695 19947 24701
rect 20622 24692 20628 24704
rect 20680 24692 20686 24744
rect 21450 24692 21456 24744
rect 21508 24692 21514 24744
rect 22557 24735 22615 24741
rect 22557 24701 22569 24735
rect 22603 24732 22615 24735
rect 22646 24732 22652 24744
rect 22603 24704 22652 24732
rect 22603 24701 22615 24704
rect 22557 24695 22615 24701
rect 22646 24692 22652 24704
rect 22704 24692 22710 24744
rect 22738 24692 22744 24744
rect 22796 24732 22802 24744
rect 23385 24735 23443 24741
rect 23385 24732 23397 24735
rect 22796 24704 23397 24732
rect 22796 24692 22802 24704
rect 23385 24701 23397 24704
rect 23431 24732 23443 24735
rect 25516 24732 25544 24828
rect 27706 24760 27712 24812
rect 27764 24760 27770 24812
rect 28258 24760 28264 24812
rect 28316 24760 28322 24812
rect 28368 24800 28396 24840
rect 28537 24803 28595 24809
rect 28537 24800 28549 24803
rect 28368 24772 28549 24800
rect 28537 24769 28549 24772
rect 28583 24769 28595 24803
rect 28537 24763 28595 24769
rect 23431 24704 25544 24732
rect 27801 24735 27859 24741
rect 23431 24701 23443 24704
rect 23385 24695 23443 24701
rect 27801 24701 27813 24735
rect 27847 24701 27859 24735
rect 27801 24695 27859 24701
rect 12897 24667 12955 24673
rect 12897 24633 12909 24667
rect 12943 24664 12955 24667
rect 12986 24664 12992 24676
rect 12943 24636 12992 24664
rect 12943 24633 12955 24636
rect 12897 24627 12955 24633
rect 12986 24624 12992 24636
rect 13044 24624 13050 24676
rect 16132 24636 16574 24664
rect 16132 24608 16160 24636
rect 14826 24596 14832 24608
rect 12544 24568 14832 24596
rect 12437 24559 12495 24565
rect 14826 24556 14832 24568
rect 14884 24556 14890 24608
rect 16114 24556 16120 24608
rect 16172 24556 16178 24608
rect 16206 24556 16212 24608
rect 16264 24556 16270 24608
rect 16546 24596 16574 24636
rect 16776 24636 17908 24664
rect 16776 24605 16804 24636
rect 16761 24599 16819 24605
rect 16761 24596 16773 24599
rect 16546 24568 16773 24596
rect 16761 24565 16773 24568
rect 16807 24565 16819 24599
rect 16761 24559 16819 24565
rect 17126 24556 17132 24608
rect 17184 24556 17190 24608
rect 17494 24556 17500 24608
rect 17552 24556 17558 24608
rect 17880 24596 17908 24636
rect 17954 24624 17960 24676
rect 18012 24624 18018 24676
rect 21468 24664 21496 24692
rect 19444 24636 21496 24664
rect 19334 24596 19340 24608
rect 17880 24568 19340 24596
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 19444 24605 19472 24636
rect 19429 24599 19487 24605
rect 19429 24565 19441 24599
rect 19475 24565 19487 24599
rect 19429 24559 19487 24565
rect 22830 24556 22836 24608
rect 22888 24596 22894 24608
rect 23109 24599 23167 24605
rect 23109 24596 23121 24599
rect 22888 24568 23121 24596
rect 22888 24556 22894 24568
rect 23109 24565 23121 24568
rect 23155 24565 23167 24599
rect 23109 24559 23167 24565
rect 24670 24556 24676 24608
rect 24728 24596 24734 24608
rect 25774 24596 25780 24608
rect 24728 24568 25780 24596
rect 24728 24556 24734 24568
rect 25774 24556 25780 24568
rect 25832 24556 25838 24608
rect 27816 24596 27844 24695
rect 27890 24692 27896 24744
rect 27948 24692 27954 24744
rect 27982 24692 27988 24744
rect 28040 24692 28046 24744
rect 30282 24692 30288 24744
rect 30340 24692 30346 24744
rect 30193 24667 30251 24673
rect 30193 24664 30205 24667
rect 29762 24636 30205 24664
rect 30193 24633 30205 24636
rect 30239 24633 30251 24667
rect 30193 24627 30251 24633
rect 29178 24596 29184 24608
rect 27816 24568 29184 24596
rect 29178 24556 29184 24568
rect 29236 24556 29242 24608
rect 2760 24506 32200 24528
rect 2760 24454 6946 24506
rect 6998 24454 7010 24506
rect 7062 24454 7074 24506
rect 7126 24454 7138 24506
rect 7190 24454 7202 24506
rect 7254 24454 14306 24506
rect 14358 24454 14370 24506
rect 14422 24454 14434 24506
rect 14486 24454 14498 24506
rect 14550 24454 14562 24506
rect 14614 24454 21666 24506
rect 21718 24454 21730 24506
rect 21782 24454 21794 24506
rect 21846 24454 21858 24506
rect 21910 24454 21922 24506
rect 21974 24454 29026 24506
rect 29078 24454 29090 24506
rect 29142 24454 29154 24506
rect 29206 24454 29218 24506
rect 29270 24454 29282 24506
rect 29334 24454 32200 24506
rect 2760 24432 32200 24454
rect 3418 24352 3424 24404
rect 3476 24352 3482 24404
rect 3878 24352 3884 24404
rect 3936 24352 3942 24404
rect 4614 24352 4620 24404
rect 4672 24352 4678 24404
rect 5997 24395 6055 24401
rect 5997 24361 6009 24395
rect 6043 24392 6055 24395
rect 6454 24392 6460 24404
rect 6043 24364 6460 24392
rect 6043 24361 6055 24364
rect 5997 24355 6055 24361
rect 6454 24352 6460 24364
rect 6512 24352 6518 24404
rect 7282 24352 7288 24404
rect 7340 24352 7346 24404
rect 7742 24352 7748 24404
rect 7800 24392 7806 24404
rect 8665 24395 8723 24401
rect 8665 24392 8677 24395
rect 7800 24364 8677 24392
rect 7800 24352 7806 24364
rect 8665 24361 8677 24364
rect 8711 24392 8723 24395
rect 8938 24392 8944 24404
rect 8711 24364 8944 24392
rect 8711 24361 8723 24364
rect 8665 24355 8723 24361
rect 8938 24352 8944 24364
rect 8996 24392 9002 24404
rect 10686 24392 10692 24404
rect 8996 24364 9352 24392
rect 8996 24352 9002 24364
rect 4525 24327 4583 24333
rect 4525 24293 4537 24327
rect 4571 24324 4583 24327
rect 4632 24324 4660 24352
rect 4571 24296 4660 24324
rect 4571 24293 4583 24296
rect 4525 24287 4583 24293
rect 3234 24216 3240 24268
rect 3292 24256 3298 24268
rect 3789 24259 3847 24265
rect 3789 24256 3801 24259
rect 3292 24228 3801 24256
rect 3292 24216 3298 24228
rect 3789 24225 3801 24228
rect 3835 24225 3847 24259
rect 3789 24219 3847 24225
rect 4246 24216 4252 24268
rect 4304 24216 4310 24268
rect 5626 24216 5632 24268
rect 5684 24216 5690 24268
rect 3329 24191 3387 24197
rect 3329 24157 3341 24191
rect 3375 24188 3387 24191
rect 4065 24191 4123 24197
rect 4065 24188 4077 24191
rect 3375 24160 4077 24188
rect 3375 24157 3387 24160
rect 3329 24151 3387 24157
rect 4065 24157 4077 24160
rect 4111 24188 4123 24191
rect 4111 24160 4292 24188
rect 4111 24157 4123 24160
rect 4065 24151 4123 24157
rect 4264 24132 4292 24160
rect 4246 24080 4252 24132
rect 4304 24080 4310 24132
rect 7300 24120 7328 24352
rect 9122 24284 9128 24336
rect 9180 24284 9186 24336
rect 7650 24216 7656 24268
rect 7708 24256 7714 24268
rect 8941 24259 8999 24265
rect 8941 24256 8953 24259
rect 7708 24228 8953 24256
rect 7708 24216 7714 24228
rect 8941 24225 8953 24228
rect 8987 24225 8999 24259
rect 8941 24219 8999 24225
rect 8956 24188 8984 24219
rect 9030 24216 9036 24268
rect 9088 24216 9094 24268
rect 9324 24265 9352 24364
rect 10520 24364 10692 24392
rect 10520 24324 10548 24364
rect 10686 24352 10692 24364
rect 10744 24352 10750 24404
rect 10778 24352 10784 24404
rect 10836 24392 10842 24404
rect 12434 24392 12440 24404
rect 10836 24364 12440 24392
rect 10836 24352 10842 24364
rect 12434 24352 12440 24364
rect 12492 24352 12498 24404
rect 12989 24395 13047 24401
rect 12989 24361 13001 24395
rect 13035 24392 13047 24395
rect 13354 24392 13360 24404
rect 13035 24364 13360 24392
rect 13035 24361 13047 24364
rect 12989 24355 13047 24361
rect 13354 24352 13360 24364
rect 13412 24352 13418 24404
rect 21361 24395 21419 24401
rect 21361 24392 21373 24395
rect 14384 24364 21373 24392
rect 14384 24336 14412 24364
rect 21361 24361 21373 24364
rect 21407 24392 21419 24395
rect 21726 24392 21732 24404
rect 21407 24364 21732 24392
rect 21407 24361 21419 24364
rect 21361 24355 21419 24361
rect 21726 24352 21732 24364
rect 21784 24352 21790 24404
rect 22646 24352 22652 24404
rect 22704 24352 22710 24404
rect 26694 24352 26700 24404
rect 26752 24392 26758 24404
rect 26752 24364 27016 24392
rect 26752 24352 26758 24364
rect 10442 24296 10548 24324
rect 10594 24284 10600 24336
rect 10652 24324 10658 24336
rect 10873 24327 10931 24333
rect 10873 24324 10885 24327
rect 10652 24296 10885 24324
rect 10652 24284 10658 24296
rect 10873 24293 10885 24296
rect 10919 24293 10931 24327
rect 10873 24287 10931 24293
rect 13262 24284 13268 24336
rect 13320 24324 13326 24336
rect 13541 24327 13599 24333
rect 13541 24324 13553 24327
rect 13320 24296 13553 24324
rect 13320 24284 13326 24296
rect 13541 24293 13553 24296
rect 13587 24293 13599 24327
rect 13541 24287 13599 24293
rect 14366 24284 14372 24336
rect 14424 24284 14430 24336
rect 14734 24284 14740 24336
rect 14792 24284 14798 24336
rect 18138 24284 18144 24336
rect 18196 24324 18202 24336
rect 18693 24327 18751 24333
rect 18693 24324 18705 24327
rect 18196 24296 18705 24324
rect 18196 24284 18202 24296
rect 18693 24293 18705 24296
rect 18739 24293 18751 24327
rect 18693 24287 18751 24293
rect 19058 24284 19064 24336
rect 19116 24284 19122 24336
rect 19889 24327 19947 24333
rect 19889 24293 19901 24327
rect 19935 24324 19947 24327
rect 20070 24324 20076 24336
rect 19935 24296 20076 24324
rect 19935 24293 19947 24296
rect 19889 24287 19947 24293
rect 20070 24284 20076 24296
rect 20128 24284 20134 24336
rect 26988 24333 27016 24364
rect 26973 24327 27031 24333
rect 26252 24296 26832 24324
rect 26252 24268 26280 24296
rect 9309 24259 9367 24265
rect 9309 24225 9321 24259
rect 9355 24225 9367 24259
rect 9309 24219 9367 24225
rect 11146 24216 11152 24268
rect 11204 24216 11210 24268
rect 11238 24216 11244 24268
rect 11296 24256 11302 24268
rect 11514 24256 11520 24268
rect 11296 24228 11520 24256
rect 11296 24216 11302 24228
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 12437 24259 12495 24265
rect 12437 24256 12449 24259
rect 11655 24228 12449 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 12437 24225 12449 24228
rect 12483 24256 12495 24259
rect 12618 24256 12624 24268
rect 12483 24228 12624 24256
rect 12483 24225 12495 24228
rect 12437 24219 12495 24225
rect 12618 24216 12624 24228
rect 12676 24216 12682 24268
rect 15838 24216 15844 24268
rect 15896 24216 15902 24268
rect 17037 24259 17095 24265
rect 17037 24225 17049 24259
rect 17083 24256 17095 24259
rect 17126 24256 17132 24268
rect 17083 24228 17132 24256
rect 17083 24225 17095 24228
rect 17037 24219 17095 24225
rect 10778 24188 10784 24200
rect 8956 24160 10784 24188
rect 10778 24148 10784 24160
rect 10836 24148 10842 24200
rect 11532 24188 11560 24216
rect 12713 24191 12771 24197
rect 12713 24188 12725 24191
rect 11532 24160 12725 24188
rect 12713 24157 12725 24160
rect 12759 24188 12771 24191
rect 13906 24188 13912 24200
rect 12759 24160 13912 24188
rect 12759 24157 12771 24160
rect 12713 24151 12771 24157
rect 13906 24148 13912 24160
rect 13964 24148 13970 24200
rect 14458 24148 14464 24200
rect 14516 24148 14522 24200
rect 16209 24191 16267 24197
rect 16209 24157 16221 24191
rect 16255 24188 16267 24191
rect 16853 24191 16911 24197
rect 16853 24188 16865 24191
rect 16255 24160 16865 24188
rect 16255 24157 16267 24160
rect 16209 24151 16267 24157
rect 16853 24157 16865 24160
rect 16899 24157 16911 24191
rect 16853 24151 16911 24157
rect 7300 24092 8892 24120
rect 5902 24012 5908 24064
rect 5960 24052 5966 24064
rect 6641 24055 6699 24061
rect 6641 24052 6653 24055
rect 5960 24024 6653 24052
rect 5960 24012 5966 24024
rect 6641 24021 6653 24024
rect 6687 24021 6699 24055
rect 6641 24015 6699 24021
rect 8754 24012 8760 24064
rect 8812 24012 8818 24064
rect 8864 24052 8892 24092
rect 11900 24092 12848 24120
rect 9401 24055 9459 24061
rect 9401 24052 9413 24055
rect 8864 24024 9413 24052
rect 9401 24021 9413 24024
rect 9447 24021 9459 24055
rect 9401 24015 9459 24021
rect 11514 24012 11520 24064
rect 11572 24052 11578 24064
rect 11900 24061 11928 24092
rect 11885 24055 11943 24061
rect 11885 24052 11897 24055
rect 11572 24024 11897 24052
rect 11572 24012 11578 24024
rect 11885 24021 11897 24024
rect 11931 24021 11943 24055
rect 11885 24015 11943 24021
rect 12250 24012 12256 24064
rect 12308 24012 12314 24064
rect 12820 24061 12848 24092
rect 16022 24080 16028 24132
rect 16080 24120 16086 24132
rect 17052 24120 17080 24219
rect 17126 24216 17132 24228
rect 17184 24216 17190 24268
rect 18509 24259 18567 24265
rect 18509 24256 18521 24259
rect 17512 24228 18521 24256
rect 17512 24200 17540 24228
rect 18509 24225 18521 24228
rect 18555 24225 18567 24259
rect 18509 24219 18567 24225
rect 18601 24259 18659 24265
rect 18601 24225 18613 24259
rect 18647 24225 18659 24259
rect 18601 24219 18659 24225
rect 17221 24191 17279 24197
rect 17221 24157 17233 24191
rect 17267 24188 17279 24191
rect 17494 24188 17500 24200
rect 17267 24160 17500 24188
rect 17267 24157 17279 24160
rect 17221 24151 17279 24157
rect 16080 24092 17080 24120
rect 16080 24080 16086 24092
rect 12805 24055 12863 24061
rect 12805 24021 12817 24055
rect 12851 24052 12863 24055
rect 14918 24052 14924 24064
rect 12851 24024 14924 24052
rect 12851 24021 12863 24024
rect 12805 24015 12863 24021
rect 14918 24012 14924 24024
rect 14976 24012 14982 24064
rect 15286 24012 15292 24064
rect 15344 24052 15350 24064
rect 16206 24052 16212 24064
rect 15344 24024 16212 24052
rect 15344 24012 15350 24024
rect 16206 24012 16212 24024
rect 16264 24052 16270 24064
rect 16301 24055 16359 24061
rect 16301 24052 16313 24055
rect 16264 24024 16313 24052
rect 16264 24012 16270 24024
rect 16301 24021 16313 24024
rect 16347 24021 16359 24055
rect 16301 24015 16359 24021
rect 16942 24012 16948 24064
rect 17000 24052 17006 24064
rect 17236 24052 17264 24151
rect 17494 24148 17500 24160
rect 17552 24148 17558 24200
rect 18616 24188 18644 24219
rect 18874 24216 18880 24268
rect 18932 24216 18938 24268
rect 19150 24216 19156 24268
rect 19208 24216 19214 24268
rect 21545 24259 21603 24265
rect 21545 24225 21557 24259
rect 21591 24256 21603 24259
rect 22281 24259 22339 24265
rect 21591 24228 21772 24256
rect 21591 24225 21603 24228
rect 21545 24219 21603 24225
rect 19426 24188 19432 24200
rect 18616 24160 19432 24188
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 17954 24080 17960 24132
rect 18012 24120 18018 24132
rect 18325 24123 18383 24129
rect 18325 24120 18337 24123
rect 18012 24092 18337 24120
rect 18012 24080 18018 24092
rect 18325 24089 18337 24092
rect 18371 24089 18383 24123
rect 18325 24083 18383 24089
rect 17000 24024 17264 24052
rect 17000 24012 17006 24024
rect 18874 24012 18880 24064
rect 18932 24052 18938 24064
rect 19429 24055 19487 24061
rect 19429 24052 19441 24055
rect 18932 24024 19441 24052
rect 18932 24012 18938 24024
rect 19429 24021 19441 24024
rect 19475 24021 19487 24055
rect 19429 24015 19487 24021
rect 21450 24012 21456 24064
rect 21508 24052 21514 24064
rect 21637 24055 21695 24061
rect 21637 24052 21649 24055
rect 21508 24024 21649 24052
rect 21508 24012 21514 24024
rect 21637 24021 21649 24024
rect 21683 24021 21695 24055
rect 21744 24052 21772 24228
rect 22281 24225 22293 24259
rect 22327 24256 22339 24259
rect 24118 24256 24124 24268
rect 22327 24228 24124 24256
rect 22327 24225 22339 24228
rect 22281 24219 22339 24225
rect 24118 24216 24124 24228
rect 24176 24216 24182 24268
rect 25130 24216 25136 24268
rect 25188 24265 25194 24268
rect 25188 24256 25199 24265
rect 25188 24228 25233 24256
rect 25188 24219 25199 24228
rect 25188 24216 25194 24219
rect 25406 24216 25412 24268
rect 25464 24216 25470 24268
rect 25590 24216 25596 24268
rect 25648 24216 25654 24268
rect 25866 24216 25872 24268
rect 25924 24256 25930 24268
rect 26234 24256 26240 24268
rect 25924 24228 26240 24256
rect 25924 24216 25930 24228
rect 26234 24216 26240 24228
rect 26292 24216 26298 24268
rect 26513 24259 26571 24265
rect 26513 24225 26525 24259
rect 26559 24225 26571 24259
rect 26513 24219 26571 24225
rect 22097 24191 22155 24197
rect 22097 24157 22109 24191
rect 22143 24157 22155 24191
rect 22097 24151 22155 24157
rect 22112 24120 22140 24151
rect 22186 24148 22192 24200
rect 22244 24148 22250 24200
rect 24302 24148 24308 24200
rect 24360 24148 24366 24200
rect 26528 24188 26556 24219
rect 26602 24216 26608 24268
rect 26660 24216 26666 24268
rect 26804 24265 26832 24296
rect 26973 24293 26985 24327
rect 27019 24324 27031 24327
rect 27890 24324 27896 24336
rect 27019 24296 27896 24324
rect 27019 24293 27031 24296
rect 26973 24287 27031 24293
rect 27890 24284 27896 24296
rect 27948 24284 27954 24336
rect 26789 24259 26847 24265
rect 26789 24225 26801 24259
rect 26835 24225 26847 24259
rect 26789 24219 26847 24225
rect 28629 24191 28687 24197
rect 28629 24188 28641 24191
rect 26528 24160 28641 24188
rect 28629 24157 28641 24160
rect 28675 24157 28687 24191
rect 28629 24151 28687 24157
rect 29273 24191 29331 24197
rect 29273 24157 29285 24191
rect 29319 24188 29331 24191
rect 30374 24188 30380 24200
rect 29319 24160 30380 24188
rect 29319 24157 29331 24160
rect 29273 24151 29331 24157
rect 24210 24120 24216 24132
rect 22112 24092 24216 24120
rect 24210 24080 24216 24092
rect 24268 24120 24274 24132
rect 25777 24123 25835 24129
rect 25777 24120 25789 24123
rect 24268 24092 25789 24120
rect 24268 24080 24274 24092
rect 25777 24089 25789 24092
rect 25823 24089 25835 24123
rect 28644 24120 28672 24151
rect 30374 24148 30380 24160
rect 30432 24148 30438 24200
rect 31570 24148 31576 24200
rect 31628 24148 31634 24200
rect 31849 24191 31907 24197
rect 31849 24157 31861 24191
rect 31895 24188 31907 24191
rect 33134 24188 33140 24200
rect 31895 24160 33140 24188
rect 31895 24157 31907 24160
rect 31849 24151 31907 24157
rect 33134 24148 33140 24160
rect 33192 24148 33198 24200
rect 29454 24120 29460 24132
rect 28644 24092 29460 24120
rect 25777 24083 25835 24089
rect 29454 24080 29460 24092
rect 29512 24080 29518 24132
rect 22094 24052 22100 24064
rect 21744 24024 22100 24052
rect 21637 24015 21695 24021
rect 22094 24012 22100 24024
rect 22152 24012 22158 24064
rect 23934 24012 23940 24064
rect 23992 24052 23998 24064
rect 24854 24052 24860 24064
rect 23992 24024 24860 24052
rect 23992 24012 23998 24024
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 24946 24012 24952 24064
rect 25004 24052 25010 24064
rect 25041 24055 25099 24061
rect 25041 24052 25053 24055
rect 25004 24024 25053 24052
rect 25004 24012 25010 24024
rect 25041 24021 25053 24024
rect 25087 24021 25099 24055
rect 25041 24015 25099 24021
rect 25130 24012 25136 24064
rect 25188 24052 25194 24064
rect 28074 24052 28080 24064
rect 25188 24024 28080 24052
rect 25188 24012 25194 24024
rect 28074 24012 28080 24024
rect 28132 24012 28138 24064
rect 2760 23962 32200 23984
rect 2760 23910 6286 23962
rect 6338 23910 6350 23962
rect 6402 23910 6414 23962
rect 6466 23910 6478 23962
rect 6530 23910 6542 23962
rect 6594 23910 13646 23962
rect 13698 23910 13710 23962
rect 13762 23910 13774 23962
rect 13826 23910 13838 23962
rect 13890 23910 13902 23962
rect 13954 23910 21006 23962
rect 21058 23910 21070 23962
rect 21122 23910 21134 23962
rect 21186 23910 21198 23962
rect 21250 23910 21262 23962
rect 21314 23910 28366 23962
rect 28418 23910 28430 23962
rect 28482 23910 28494 23962
rect 28546 23910 28558 23962
rect 28610 23910 28622 23962
rect 28674 23910 32200 23962
rect 2760 23888 32200 23910
rect 3145 23851 3203 23857
rect 3145 23817 3157 23851
rect 3191 23848 3203 23851
rect 3234 23848 3240 23860
rect 3191 23820 3240 23848
rect 3191 23817 3203 23820
rect 3145 23811 3203 23817
rect 3234 23808 3240 23820
rect 3292 23808 3298 23860
rect 4154 23808 4160 23860
rect 4212 23848 4218 23860
rect 7653 23851 7711 23857
rect 4212 23820 5856 23848
rect 4212 23808 4218 23820
rect 4522 23672 4528 23724
rect 4580 23712 4586 23724
rect 4617 23715 4675 23721
rect 4617 23712 4629 23715
rect 4580 23684 4629 23712
rect 4580 23672 4586 23684
rect 4617 23681 4629 23684
rect 4663 23681 4675 23715
rect 4617 23675 4675 23681
rect 4893 23715 4951 23721
rect 4893 23681 4905 23715
rect 4939 23712 4951 23715
rect 5718 23712 5724 23724
rect 4939 23684 5724 23712
rect 4939 23681 4951 23684
rect 4893 23675 4951 23681
rect 5718 23672 5724 23684
rect 5776 23672 5782 23724
rect 5828 23712 5856 23820
rect 7653 23817 7665 23851
rect 7699 23848 7711 23851
rect 7742 23848 7748 23860
rect 7699 23820 7748 23848
rect 7699 23817 7711 23820
rect 7653 23811 7711 23817
rect 7742 23808 7748 23820
rect 7800 23808 7806 23860
rect 7834 23808 7840 23860
rect 7892 23848 7898 23860
rect 11054 23848 11060 23860
rect 7892 23820 11060 23848
rect 7892 23808 7898 23820
rect 11054 23808 11060 23820
rect 11112 23808 11118 23860
rect 11146 23808 11152 23860
rect 11204 23848 11210 23860
rect 11330 23848 11336 23860
rect 11204 23820 11336 23848
rect 11204 23808 11210 23820
rect 11330 23808 11336 23820
rect 11388 23808 11394 23860
rect 11422 23808 11428 23860
rect 11480 23848 11486 23860
rect 11480 23820 12434 23848
rect 11480 23808 11486 23820
rect 7009 23715 7067 23721
rect 7009 23712 7021 23715
rect 5828 23684 7021 23712
rect 7009 23681 7021 23684
rect 7055 23681 7067 23715
rect 7760 23712 7788 23808
rect 12406 23780 12434 23820
rect 12986 23808 12992 23860
rect 13044 23808 13050 23860
rect 13998 23808 14004 23860
rect 14056 23808 14062 23860
rect 14366 23808 14372 23860
rect 14424 23808 14430 23860
rect 15838 23808 15844 23860
rect 15896 23848 15902 23860
rect 16577 23851 16635 23857
rect 16577 23848 16589 23851
rect 15896 23820 16589 23848
rect 15896 23808 15902 23820
rect 16577 23817 16589 23820
rect 16623 23817 16635 23851
rect 16577 23811 16635 23817
rect 17862 23808 17868 23860
rect 17920 23848 17926 23860
rect 18322 23848 18328 23860
rect 17920 23820 18328 23848
rect 17920 23808 17926 23820
rect 18322 23808 18328 23820
rect 18380 23808 18386 23860
rect 18414 23808 18420 23860
rect 18472 23808 18478 23860
rect 25314 23808 25320 23860
rect 25372 23848 25378 23860
rect 25777 23851 25835 23857
rect 25777 23848 25789 23851
rect 25372 23820 25789 23848
rect 25372 23808 25378 23820
rect 25777 23817 25789 23820
rect 25823 23817 25835 23851
rect 26694 23848 26700 23860
rect 25777 23811 25835 23817
rect 26252 23820 26700 23848
rect 13906 23780 13912 23792
rect 12406 23752 13912 23780
rect 13906 23740 13912 23752
rect 13964 23740 13970 23792
rect 7760 23684 8340 23712
rect 7009 23675 7067 23681
rect 5169 23647 5227 23653
rect 5169 23613 5181 23647
rect 5215 23613 5227 23647
rect 5169 23607 5227 23613
rect 6365 23647 6423 23653
rect 6365 23613 6377 23647
rect 6411 23644 6423 23647
rect 6546 23644 6552 23656
rect 6411 23616 6552 23644
rect 6411 23613 6423 23616
rect 6365 23607 6423 23613
rect 5077 23579 5135 23585
rect 4186 23548 4292 23576
rect 4264 23508 4292 23548
rect 5077 23545 5089 23579
rect 5123 23545 5135 23579
rect 5077 23539 5135 23545
rect 5092 23508 5120 23539
rect 5184 23520 5212 23607
rect 6546 23604 6552 23616
rect 6604 23604 6610 23656
rect 7742 23604 7748 23656
rect 7800 23644 7806 23656
rect 8312 23653 8340 23684
rect 8386 23672 8392 23724
rect 8444 23672 8450 23724
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23712 8723 23715
rect 8754 23712 8760 23724
rect 8711 23684 8760 23712
rect 8711 23681 8723 23684
rect 8665 23675 8723 23681
rect 8754 23672 8760 23684
rect 8812 23672 8818 23724
rect 11330 23672 11336 23724
rect 11388 23712 11394 23724
rect 12250 23712 12256 23724
rect 11388 23684 12256 23712
rect 11388 23672 11394 23684
rect 12250 23672 12256 23684
rect 12308 23712 12314 23724
rect 12897 23715 12955 23721
rect 12897 23712 12909 23715
rect 12308 23684 12909 23712
rect 12308 23672 12314 23684
rect 12897 23681 12909 23684
rect 12943 23712 12955 23715
rect 14384 23712 14412 23808
rect 15194 23740 15200 23792
rect 15252 23780 15258 23792
rect 15654 23780 15660 23792
rect 15252 23752 15660 23780
rect 15252 23740 15258 23752
rect 15654 23740 15660 23752
rect 15712 23780 15718 23792
rect 16117 23783 16175 23789
rect 16117 23780 16129 23783
rect 15712 23752 16129 23780
rect 15712 23740 15718 23752
rect 16117 23749 16129 23752
rect 16163 23749 16175 23783
rect 16117 23743 16175 23749
rect 14826 23712 14832 23724
rect 12943 23684 14412 23712
rect 14476 23684 14832 23712
rect 12943 23681 12955 23684
rect 12897 23675 12955 23681
rect 7929 23647 7987 23653
rect 7929 23644 7941 23647
rect 7800 23616 7941 23644
rect 7800 23604 7806 23616
rect 7929 23613 7941 23616
rect 7975 23613 7987 23647
rect 7929 23607 7987 23613
rect 8297 23647 8355 23653
rect 8297 23613 8309 23647
rect 8343 23613 8355 23647
rect 8297 23607 8355 23613
rect 10413 23647 10471 23653
rect 10413 23613 10425 23647
rect 10459 23644 10471 23647
rect 11974 23644 11980 23656
rect 10459 23616 11980 23644
rect 10459 23613 10471 23616
rect 10413 23607 10471 23613
rect 11974 23604 11980 23616
rect 12032 23604 12038 23656
rect 13538 23604 13544 23656
rect 13596 23604 13602 23656
rect 14292 23653 14320 23684
rect 14093 23647 14151 23653
rect 14093 23613 14105 23647
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23613 14335 23647
rect 14476 23644 14504 23684
rect 14826 23672 14832 23684
rect 14884 23712 14890 23724
rect 14884 23684 16574 23712
rect 14884 23672 14890 23684
rect 14277 23607 14335 23613
rect 14384 23616 14504 23644
rect 7650 23536 7656 23588
rect 7708 23576 7714 23588
rect 8021 23579 8079 23585
rect 8021 23576 8033 23579
rect 7708 23548 8033 23576
rect 7708 23536 7714 23548
rect 8021 23545 8033 23548
rect 8067 23545 8079 23579
rect 8021 23539 8079 23545
rect 8110 23536 8116 23588
rect 8168 23536 8174 23588
rect 10321 23579 10379 23585
rect 10321 23576 10333 23579
rect 9890 23548 10333 23576
rect 10321 23545 10333 23548
rect 10367 23545 10379 23579
rect 10321 23539 10379 23545
rect 11882 23536 11888 23588
rect 11940 23576 11946 23588
rect 14108 23576 14136 23607
rect 14384 23576 14412 23616
rect 14642 23604 14648 23656
rect 14700 23644 14706 23656
rect 15289 23647 15347 23653
rect 15289 23644 15301 23647
rect 14700 23616 15301 23644
rect 14700 23604 14706 23616
rect 15289 23613 15301 23616
rect 15335 23613 15347 23647
rect 15289 23607 15347 23613
rect 15378 23604 15384 23656
rect 15436 23644 15442 23656
rect 15473 23647 15531 23653
rect 15473 23644 15485 23647
rect 15436 23616 15485 23644
rect 15436 23604 15442 23616
rect 15473 23613 15485 23616
rect 15519 23613 15531 23647
rect 15473 23607 15531 23613
rect 16114 23604 16120 23656
rect 16172 23644 16178 23656
rect 16301 23647 16359 23653
rect 16301 23644 16313 23647
rect 16172 23616 16313 23644
rect 16172 23604 16178 23616
rect 16301 23613 16313 23616
rect 16347 23613 16359 23647
rect 16546 23644 16574 23684
rect 22278 23672 22284 23724
rect 22336 23712 22342 23724
rect 22557 23715 22615 23721
rect 22557 23712 22569 23715
rect 22336 23684 22569 23712
rect 22336 23672 22342 23684
rect 22557 23681 22569 23684
rect 22603 23712 22615 23715
rect 23106 23712 23112 23724
rect 22603 23684 23112 23712
rect 22603 23681 22615 23684
rect 22557 23675 22615 23681
rect 23106 23672 23112 23684
rect 23164 23672 23170 23724
rect 25317 23715 25375 23721
rect 25317 23681 25329 23715
rect 25363 23712 25375 23715
rect 25498 23712 25504 23724
rect 25363 23684 25504 23712
rect 25363 23681 25375 23684
rect 25317 23675 25375 23681
rect 25498 23672 25504 23684
rect 25556 23672 25562 23724
rect 25682 23672 25688 23724
rect 25740 23712 25746 23724
rect 25740 23684 26096 23712
rect 25740 23672 25746 23684
rect 16669 23647 16727 23653
rect 16669 23644 16681 23647
rect 16546 23616 16681 23644
rect 16301 23607 16359 23613
rect 16669 23613 16681 23616
rect 16715 23613 16727 23647
rect 16669 23607 16727 23613
rect 17586 23604 17592 23656
rect 17644 23604 17650 23656
rect 18601 23647 18659 23653
rect 18601 23644 18613 23647
rect 18340 23616 18613 23644
rect 11940 23548 14044 23576
rect 14108 23548 14412 23576
rect 11940 23536 11946 23548
rect 4264 23480 5120 23508
rect 5166 23468 5172 23520
rect 5224 23468 5230 23520
rect 5534 23468 5540 23520
rect 5592 23508 5598 23520
rect 5721 23511 5779 23517
rect 5721 23508 5733 23511
rect 5592 23480 5733 23508
rect 5592 23468 5598 23480
rect 5721 23477 5733 23480
rect 5767 23477 5779 23511
rect 5721 23471 5779 23477
rect 6454 23468 6460 23520
rect 6512 23468 6518 23520
rect 7742 23468 7748 23520
rect 7800 23468 7806 23520
rect 10137 23511 10195 23517
rect 10137 23477 10149 23511
rect 10183 23508 10195 23511
rect 10686 23508 10692 23520
rect 10183 23480 10692 23508
rect 10183 23477 10195 23480
rect 10137 23471 10195 23477
rect 10686 23468 10692 23480
rect 10744 23468 10750 23520
rect 12529 23511 12587 23517
rect 12529 23477 12541 23511
rect 12575 23508 12587 23511
rect 13446 23508 13452 23520
rect 12575 23480 13452 23508
rect 12575 23477 12587 23480
rect 12529 23471 12587 23477
rect 13446 23468 13452 23480
rect 13504 23468 13510 23520
rect 14016 23508 14044 23548
rect 14458 23536 14464 23588
rect 14516 23576 14522 23588
rect 15105 23579 15163 23585
rect 15105 23576 15117 23579
rect 14516 23548 15117 23576
rect 14516 23536 14522 23548
rect 15105 23545 15117 23548
rect 15151 23576 15163 23579
rect 15746 23576 15752 23588
rect 15151 23548 15752 23576
rect 15151 23545 15163 23548
rect 15105 23539 15163 23545
rect 15746 23536 15752 23548
rect 15804 23536 15810 23588
rect 18340 23520 18368 23616
rect 18601 23613 18613 23616
rect 18647 23613 18659 23647
rect 18601 23607 18659 23613
rect 18690 23604 18696 23656
rect 18748 23604 18754 23656
rect 19702 23604 19708 23656
rect 19760 23604 19766 23656
rect 20441 23647 20499 23653
rect 20441 23613 20453 23647
rect 20487 23613 20499 23647
rect 20441 23607 20499 23613
rect 20456 23576 20484 23607
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 21545 23647 21603 23653
rect 21545 23644 21557 23647
rect 20956 23616 21557 23644
rect 20956 23604 20962 23616
rect 21545 23613 21557 23616
rect 21591 23613 21603 23647
rect 21545 23607 21603 23613
rect 21726 23604 21732 23656
rect 21784 23644 21790 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 21784 23616 21833 23644
rect 21784 23604 21790 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 22094 23644 22100 23656
rect 21821 23607 21879 23613
rect 22066 23604 22100 23644
rect 22152 23644 22158 23656
rect 26068 23653 26096 23684
rect 26252 23653 26280 23820
rect 26694 23808 26700 23820
rect 26752 23808 26758 23860
rect 27617 23851 27675 23857
rect 27617 23817 27629 23851
rect 27663 23848 27675 23851
rect 27982 23848 27988 23860
rect 27663 23820 27988 23848
rect 27663 23817 27675 23820
rect 27617 23811 27675 23817
rect 26418 23740 26424 23792
rect 26476 23740 26482 23792
rect 27632 23780 27660 23811
rect 27982 23808 27988 23820
rect 28040 23808 28046 23860
rect 29181 23783 29239 23789
rect 29181 23780 29193 23783
rect 26528 23752 27660 23780
rect 27723 23752 29193 23780
rect 23017 23647 23075 23653
rect 23017 23644 23029 23647
rect 22152 23616 23029 23644
rect 22152 23604 22158 23616
rect 23017 23613 23029 23616
rect 23063 23644 23075 23647
rect 25593 23647 25651 23653
rect 25593 23644 25605 23647
rect 23063 23616 23428 23644
rect 23063 23613 23075 23616
rect 23017 23607 23075 23613
rect 20530 23576 20536 23588
rect 20456 23548 20536 23576
rect 20530 23536 20536 23548
rect 20588 23576 20594 23588
rect 22066 23576 22094 23604
rect 23400 23588 23428 23616
rect 25332 23616 25605 23644
rect 20588 23548 22094 23576
rect 20588 23536 20594 23548
rect 23382 23536 23388 23588
rect 23440 23536 23446 23588
rect 24946 23576 24952 23588
rect 24610 23548 24952 23576
rect 24946 23536 24952 23548
rect 25004 23536 25010 23588
rect 25041 23579 25099 23585
rect 25041 23545 25053 23579
rect 25087 23576 25099 23579
rect 25130 23576 25136 23588
rect 25087 23548 25136 23576
rect 25087 23545 25099 23548
rect 25041 23539 25099 23545
rect 25130 23536 25136 23548
rect 25188 23536 25194 23588
rect 14642 23508 14648 23520
rect 14016 23480 14648 23508
rect 14642 23468 14648 23480
rect 14700 23468 14706 23520
rect 15381 23511 15439 23517
rect 15381 23477 15393 23511
rect 15427 23508 15439 23511
rect 15470 23508 15476 23520
rect 15427 23480 15476 23508
rect 15427 23477 15439 23480
rect 15381 23471 15439 23477
rect 15470 23468 15476 23480
rect 15528 23468 15534 23520
rect 15562 23468 15568 23520
rect 15620 23508 15626 23520
rect 15933 23511 15991 23517
rect 15933 23508 15945 23511
rect 15620 23480 15945 23508
rect 15620 23468 15626 23480
rect 15933 23477 15945 23480
rect 15979 23508 15991 23511
rect 16022 23508 16028 23520
rect 15979 23480 16028 23508
rect 15979 23477 15991 23480
rect 15933 23471 15991 23477
rect 16022 23468 16028 23480
rect 16080 23468 16086 23520
rect 16945 23511 17003 23517
rect 16945 23477 16957 23511
rect 16991 23508 17003 23511
rect 17034 23508 17040 23520
rect 16991 23480 17040 23508
rect 16991 23477 17003 23480
rect 16945 23471 17003 23477
rect 17034 23468 17040 23480
rect 17092 23468 17098 23520
rect 17957 23511 18015 23517
rect 17957 23477 17969 23511
rect 18003 23508 18015 23511
rect 18322 23508 18328 23520
rect 18003 23480 18328 23508
rect 18003 23477 18015 23480
rect 17957 23471 18015 23477
rect 18322 23468 18328 23480
rect 18380 23468 18386 23520
rect 18874 23468 18880 23520
rect 18932 23468 18938 23520
rect 19058 23468 19064 23520
rect 19116 23468 19122 23520
rect 20346 23468 20352 23520
rect 20404 23468 20410 23520
rect 20990 23468 20996 23520
rect 21048 23468 21054 23520
rect 23109 23511 23167 23517
rect 23109 23477 23121 23511
rect 23155 23508 23167 23511
rect 23474 23508 23480 23520
rect 23155 23480 23480 23508
rect 23155 23477 23167 23480
rect 23109 23471 23167 23477
rect 23474 23468 23480 23480
rect 23532 23468 23538 23520
rect 23569 23511 23627 23517
rect 23569 23477 23581 23511
rect 23615 23508 23627 23511
rect 24394 23508 24400 23520
rect 23615 23480 24400 23508
rect 23615 23477 23627 23480
rect 23569 23471 23627 23477
rect 24394 23468 24400 23480
rect 24452 23468 24458 23520
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 25332 23508 25360 23616
rect 25593 23613 25605 23616
rect 25639 23613 25651 23647
rect 25593 23607 25651 23613
rect 25869 23647 25927 23653
rect 25869 23613 25881 23647
rect 25915 23613 25927 23647
rect 25869 23607 25927 23613
rect 26053 23647 26111 23653
rect 26053 23613 26065 23647
rect 26099 23613 26111 23647
rect 26053 23607 26111 23613
rect 26237 23647 26295 23653
rect 26237 23613 26249 23647
rect 26283 23613 26295 23647
rect 26237 23607 26295 23613
rect 24912 23480 25360 23508
rect 25409 23511 25467 23517
rect 24912 23468 24918 23480
rect 25409 23477 25421 23511
rect 25455 23508 25467 23511
rect 25774 23508 25780 23520
rect 25455 23480 25780 23508
rect 25455 23477 25467 23480
rect 25409 23471 25467 23477
rect 25774 23468 25780 23480
rect 25832 23468 25838 23520
rect 25884 23508 25912 23607
rect 26068 23576 26096 23607
rect 26326 23604 26332 23656
rect 26384 23604 26390 23656
rect 26418 23604 26424 23656
rect 26476 23604 26482 23656
rect 26528 23646 26556 23752
rect 26605 23657 26663 23663
rect 26605 23646 26617 23657
rect 26528 23623 26617 23646
rect 26651 23623 26663 23657
rect 26528 23618 26663 23623
rect 26528 23576 26556 23618
rect 26605 23617 26663 23618
rect 26694 23604 26700 23656
rect 26752 23604 26758 23656
rect 26878 23604 26884 23656
rect 26936 23604 26942 23656
rect 27723 23653 27751 23752
rect 29181 23749 29193 23752
rect 29227 23780 29239 23783
rect 29638 23780 29644 23792
rect 29227 23752 29644 23780
rect 29227 23749 29239 23752
rect 29181 23743 29239 23749
rect 29638 23740 29644 23752
rect 29696 23740 29702 23792
rect 27708 23647 27766 23653
rect 27708 23613 27720 23647
rect 27754 23613 27766 23647
rect 27708 23607 27766 23613
rect 27798 23604 27804 23656
rect 27856 23644 27862 23656
rect 28810 23644 28816 23656
rect 27856 23616 28816 23644
rect 27856 23604 27862 23616
rect 28810 23604 28816 23616
rect 28868 23604 28874 23656
rect 26068 23548 26556 23576
rect 27982 23536 27988 23588
rect 28040 23576 28046 23588
rect 28905 23579 28963 23585
rect 28905 23576 28917 23579
rect 28040 23548 28917 23576
rect 28040 23536 28046 23548
rect 28905 23545 28917 23548
rect 28951 23545 28963 23579
rect 28905 23539 28963 23545
rect 26050 23508 26056 23520
rect 25884 23480 26056 23508
rect 26050 23468 26056 23480
rect 26108 23468 26114 23520
rect 27065 23511 27123 23517
rect 27065 23477 27077 23511
rect 27111 23508 27123 23511
rect 27338 23508 27344 23520
rect 27111 23480 27344 23508
rect 27111 23477 27123 23480
rect 27065 23471 27123 23477
rect 27338 23468 27344 23480
rect 27396 23468 27402 23520
rect 29362 23468 29368 23520
rect 29420 23468 29426 23520
rect 2760 23418 32200 23440
rect 2760 23366 6946 23418
rect 6998 23366 7010 23418
rect 7062 23366 7074 23418
rect 7126 23366 7138 23418
rect 7190 23366 7202 23418
rect 7254 23366 14306 23418
rect 14358 23366 14370 23418
rect 14422 23366 14434 23418
rect 14486 23366 14498 23418
rect 14550 23366 14562 23418
rect 14614 23366 21666 23418
rect 21718 23366 21730 23418
rect 21782 23366 21794 23418
rect 21846 23366 21858 23418
rect 21910 23366 21922 23418
rect 21974 23366 29026 23418
rect 29078 23366 29090 23418
rect 29142 23366 29154 23418
rect 29206 23366 29218 23418
rect 29270 23366 29282 23418
rect 29334 23366 32200 23418
rect 2760 23344 32200 23366
rect 3973 23307 4031 23313
rect 3973 23273 3985 23307
rect 4019 23304 4031 23307
rect 4154 23304 4160 23316
rect 4019 23276 4160 23304
rect 4019 23273 4031 23276
rect 3973 23267 4031 23273
rect 4154 23264 4160 23276
rect 4212 23264 4218 23316
rect 4430 23264 4436 23316
rect 4488 23304 4494 23316
rect 5258 23304 5264 23316
rect 4488 23276 5264 23304
rect 4488 23264 4494 23276
rect 5258 23264 5264 23276
rect 5316 23304 5322 23316
rect 6181 23307 6239 23313
rect 5316 23276 6132 23304
rect 5316 23264 5322 23276
rect 4982 23196 4988 23248
rect 5040 23196 5046 23248
rect 5445 23239 5503 23245
rect 5445 23205 5457 23239
rect 5491 23236 5503 23239
rect 5534 23236 5540 23248
rect 5491 23208 5540 23236
rect 5491 23205 5503 23208
rect 5445 23199 5503 23205
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 6104 23236 6132 23276
rect 6181 23273 6193 23307
rect 6227 23304 6239 23307
rect 6454 23304 6460 23316
rect 6227 23276 6460 23304
rect 6227 23273 6239 23276
rect 6181 23267 6239 23273
rect 6454 23264 6460 23276
rect 6512 23264 6518 23316
rect 6546 23264 6552 23316
rect 6604 23264 6610 23316
rect 9674 23264 9680 23316
rect 9732 23304 9738 23316
rect 11054 23304 11060 23316
rect 9732 23276 11060 23304
rect 9732 23264 9738 23276
rect 11054 23264 11060 23276
rect 11112 23304 11118 23316
rect 12897 23307 12955 23313
rect 12897 23304 12909 23307
rect 11112 23276 12909 23304
rect 11112 23264 11118 23276
rect 7009 23239 7067 23245
rect 7009 23236 7021 23239
rect 6104 23208 7021 23236
rect 7009 23205 7021 23208
rect 7055 23236 7067 23239
rect 7098 23236 7104 23248
rect 7055 23208 7104 23236
rect 7055 23205 7067 23208
rect 7009 23199 7067 23205
rect 7098 23196 7104 23208
rect 7156 23236 7162 23248
rect 8202 23236 8208 23248
rect 7156 23208 8208 23236
rect 7156 23196 7162 23208
rect 8202 23196 8208 23208
rect 8260 23196 8266 23248
rect 8757 23239 8815 23245
rect 8757 23205 8769 23239
rect 8803 23236 8815 23239
rect 10689 23239 10747 23245
rect 10689 23236 10701 23239
rect 8803 23208 10701 23236
rect 8803 23205 8815 23208
rect 8757 23199 8815 23205
rect 10689 23205 10701 23208
rect 10735 23236 10747 23239
rect 10965 23239 11023 23245
rect 10965 23236 10977 23239
rect 10735 23208 10977 23236
rect 10735 23205 10747 23208
rect 10689 23199 10747 23205
rect 10965 23205 10977 23208
rect 11011 23236 11023 23239
rect 11330 23236 11336 23248
rect 11011 23208 11336 23236
rect 11011 23205 11023 23208
rect 10965 23199 11023 23205
rect 11330 23196 11336 23208
rect 11388 23196 11394 23248
rect 5718 23128 5724 23180
rect 5776 23128 5782 23180
rect 7742 23128 7748 23180
rect 7800 23128 7806 23180
rect 9493 23171 9551 23177
rect 9493 23168 9505 23171
rect 8404 23140 9505 23168
rect 8404 23112 8432 23140
rect 9493 23137 9505 23140
rect 9539 23137 9551 23171
rect 12544 23168 12572 23276
rect 12897 23273 12909 23276
rect 12943 23273 12955 23307
rect 12897 23267 12955 23273
rect 13173 23307 13231 23313
rect 13173 23273 13185 23307
rect 13219 23304 13231 23307
rect 13538 23304 13544 23316
rect 13219 23276 13544 23304
rect 13219 23273 13231 23276
rect 13173 23267 13231 23273
rect 13538 23264 13544 23276
rect 13596 23264 13602 23316
rect 14734 23264 14740 23316
rect 14792 23304 14798 23316
rect 15013 23307 15071 23313
rect 15013 23304 15025 23307
rect 14792 23276 15025 23304
rect 14792 23264 14798 23276
rect 15013 23273 15025 23276
rect 15059 23273 15071 23307
rect 15013 23267 15071 23273
rect 17586 23264 17592 23316
rect 17644 23264 17650 23316
rect 18509 23307 18567 23313
rect 18509 23273 18521 23307
rect 18555 23304 18567 23307
rect 18690 23304 18696 23316
rect 18555 23276 18696 23304
rect 18555 23273 18567 23276
rect 18509 23267 18567 23273
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 25222 23264 25228 23316
rect 25280 23304 25286 23316
rect 25590 23304 25596 23316
rect 25280 23276 25596 23304
rect 25280 23264 25286 23276
rect 25590 23264 25596 23276
rect 25648 23264 25654 23316
rect 26234 23264 26240 23316
rect 26292 23304 26298 23316
rect 26292 23276 27660 23304
rect 26292 23264 26298 23276
rect 13457 23239 13515 23245
rect 13457 23205 13469 23239
rect 13503 23236 13515 23239
rect 14090 23236 14096 23248
rect 13503 23208 14096 23236
rect 13503 23205 13515 23208
rect 13457 23199 13515 23205
rect 14090 23196 14096 23208
rect 14148 23196 14154 23248
rect 14645 23239 14703 23245
rect 14645 23205 14657 23239
rect 14691 23236 14703 23239
rect 15286 23236 15292 23248
rect 14691 23208 15292 23236
rect 14691 23205 14703 23208
rect 14645 23199 14703 23205
rect 15286 23196 15292 23208
rect 15344 23196 15350 23248
rect 15838 23196 15844 23248
rect 15896 23236 15902 23248
rect 19245 23239 19303 23245
rect 15896 23208 16606 23236
rect 15896 23196 15902 23208
rect 19245 23205 19257 23239
rect 19291 23236 19303 23239
rect 19334 23236 19340 23248
rect 19291 23208 19340 23236
rect 19291 23205 19303 23208
rect 19245 23199 19303 23205
rect 19334 23196 19340 23208
rect 19392 23196 19398 23248
rect 20346 23196 20352 23248
rect 20404 23196 20410 23248
rect 20990 23196 20996 23248
rect 21048 23196 21054 23248
rect 21450 23196 21456 23248
rect 21508 23236 21514 23248
rect 25498 23236 25504 23248
rect 21508 23208 21666 23236
rect 24412 23208 25504 23236
rect 21508 23196 21514 23208
rect 13311 23171 13369 23177
rect 13311 23168 13323 23171
rect 12544 23140 13323 23168
rect 9493 23131 9551 23137
rect 13311 23137 13323 23140
rect 13357 23137 13369 23171
rect 13311 23131 13369 23137
rect 13538 23128 13544 23180
rect 13596 23128 13602 23180
rect 13725 23171 13783 23177
rect 13725 23137 13737 23171
rect 13771 23168 13783 23171
rect 14274 23168 14280 23180
rect 13771 23140 14280 23168
rect 13771 23137 13783 23140
rect 13725 23131 13783 23137
rect 5902 23100 5908 23112
rect 5644 23072 5908 23100
rect 5644 22976 5672 23072
rect 5902 23060 5908 23072
rect 5960 23060 5966 23112
rect 6089 23103 6147 23109
rect 6089 23069 6101 23103
rect 6135 23100 6147 23103
rect 6730 23100 6736 23112
rect 6135 23072 6736 23100
rect 6135 23069 6147 23072
rect 6089 23063 6147 23069
rect 6730 23060 6736 23072
rect 6788 23060 6794 23112
rect 8386 23060 8392 23112
rect 8444 23060 8450 23112
rect 8662 23060 8668 23112
rect 8720 23060 8726 23112
rect 9953 23103 10011 23109
rect 9953 23069 9965 23103
rect 9999 23100 10011 23103
rect 10962 23100 10968 23112
rect 9999 23072 10968 23100
rect 9999 23069 10011 23072
rect 9953 23063 10011 23069
rect 10962 23060 10968 23072
rect 11020 23060 11026 23112
rect 12253 23103 12311 23109
rect 12253 23069 12265 23103
rect 12299 23100 12311 23103
rect 12526 23100 12532 23112
rect 12299 23072 12532 23100
rect 12299 23069 12311 23072
rect 12253 23063 12311 23069
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 12618 23060 12624 23112
rect 12676 23100 12682 23112
rect 13740 23100 13768 23131
rect 14274 23128 14280 23140
rect 14332 23128 14338 23180
rect 14366 23128 14372 23180
rect 14424 23177 14430 23180
rect 14424 23171 14447 23177
rect 14435 23137 14447 23171
rect 14424 23131 14447 23137
rect 14553 23171 14611 23177
rect 14553 23137 14565 23171
rect 14599 23137 14611 23171
rect 14553 23131 14611 23137
rect 14737 23171 14795 23177
rect 14737 23137 14749 23171
rect 14783 23168 14795 23171
rect 14918 23168 14924 23180
rect 14783 23140 14924 23168
rect 14783 23137 14795 23140
rect 14737 23131 14795 23137
rect 14424 23128 14430 23131
rect 12676 23072 13768 23100
rect 12676 23060 12682 23072
rect 8110 22992 8116 23044
rect 8168 23032 8174 23044
rect 13262 23032 13268 23044
rect 8168 23004 13268 23032
rect 8168 22992 8174 23004
rect 13262 22992 13268 23004
rect 13320 22992 13326 23044
rect 13446 22992 13452 23044
rect 13504 23032 13510 23044
rect 14568 23032 14596 23131
rect 14918 23128 14924 23140
rect 14976 23128 14982 23180
rect 17681 23171 17739 23177
rect 17681 23137 17693 23171
rect 17727 23168 17739 23171
rect 17862 23168 17868 23180
rect 17727 23140 17868 23168
rect 17727 23137 17739 23140
rect 17681 23131 17739 23137
rect 17862 23128 17868 23140
rect 17920 23128 17926 23180
rect 24412 23177 24440 23208
rect 25498 23196 25504 23208
rect 25556 23196 25562 23248
rect 26050 23236 26056 23248
rect 25608 23208 26056 23236
rect 24213 23171 24271 23177
rect 24213 23137 24225 23171
rect 24259 23137 24271 23171
rect 24213 23131 24271 23137
rect 24397 23171 24455 23177
rect 24397 23137 24409 23171
rect 24443 23137 24455 23171
rect 24397 23131 24455 23137
rect 15565 23103 15623 23109
rect 15565 23069 15577 23103
rect 15611 23069 15623 23103
rect 15565 23063 15623 23069
rect 14734 23032 14740 23044
rect 13504 23004 14740 23032
rect 13504 22992 13510 23004
rect 14734 22992 14740 23004
rect 14792 22992 14798 23044
rect 14921 23035 14979 23041
rect 14921 23001 14933 23035
rect 14967 23032 14979 23035
rect 15580 23032 15608 23063
rect 15746 23060 15752 23112
rect 15804 23100 15810 23112
rect 15841 23103 15899 23109
rect 15841 23100 15853 23103
rect 15804 23072 15853 23100
rect 15804 23060 15810 23072
rect 15841 23069 15853 23072
rect 15887 23069 15899 23103
rect 15841 23063 15899 23069
rect 16114 23060 16120 23112
rect 16172 23060 16178 23112
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23100 18015 23103
rect 18046 23100 18052 23112
rect 18003 23072 18052 23100
rect 18003 23069 18015 23072
rect 17957 23063 18015 23069
rect 18046 23060 18052 23072
rect 18104 23060 18110 23112
rect 18966 23060 18972 23112
rect 19024 23100 19030 23112
rect 19061 23103 19119 23109
rect 19061 23100 19073 23103
rect 19024 23072 19073 23100
rect 19024 23060 19030 23072
rect 19061 23069 19073 23072
rect 19107 23069 19119 23103
rect 19061 23063 19119 23069
rect 21269 23103 21327 23109
rect 21269 23069 21281 23103
rect 21315 23100 21327 23103
rect 22094 23100 22100 23112
rect 21315 23072 22100 23100
rect 21315 23069 21327 23072
rect 21269 23063 21327 23069
rect 22094 23060 22100 23072
rect 22152 23060 22158 23112
rect 22830 23060 22836 23112
rect 22888 23060 22894 23112
rect 23106 23060 23112 23112
rect 23164 23060 23170 23112
rect 24026 23060 24032 23112
rect 24084 23060 24090 23112
rect 14967 23004 15608 23032
rect 24228 23032 24256 23131
rect 24670 23128 24676 23180
rect 24728 23128 24734 23180
rect 25041 23171 25099 23177
rect 25041 23137 25053 23171
rect 25087 23168 25099 23171
rect 25608 23168 25636 23208
rect 26050 23196 26056 23208
rect 26108 23196 26114 23248
rect 26160 23208 27476 23236
rect 25866 23177 25872 23180
rect 25715 23171 25773 23177
rect 25715 23168 25727 23171
rect 25087 23140 25727 23168
rect 25087 23137 25099 23140
rect 25041 23131 25099 23137
rect 25715 23137 25727 23140
rect 25761 23137 25773 23171
rect 25715 23131 25773 23137
rect 25823 23171 25872 23177
rect 25823 23137 25835 23171
rect 25869 23137 25872 23171
rect 25823 23131 25872 23137
rect 25866 23128 25872 23131
rect 25924 23168 25930 23180
rect 26160 23168 26188 23208
rect 26329 23171 26387 23177
rect 26329 23168 26341 23171
rect 25924 23140 26188 23168
rect 26252 23140 26341 23168
rect 25924 23128 25930 23140
rect 24581 23103 24639 23109
rect 24581 23069 24593 23103
rect 24627 23100 24639 23103
rect 24627 23072 24900 23100
rect 24627 23069 24639 23072
rect 24581 23063 24639 23069
rect 24762 23032 24768 23044
rect 24228 23004 24768 23032
rect 14967 23001 14979 23004
rect 14921 22995 14979 23001
rect 24762 22992 24768 23004
rect 24820 22992 24826 23044
rect 24872 23032 24900 23072
rect 24946 23060 24952 23112
rect 25004 23100 25010 23112
rect 25317 23103 25375 23109
rect 25317 23100 25329 23103
rect 25004 23072 25329 23100
rect 25004 23060 25010 23072
rect 25317 23069 25329 23072
rect 25363 23069 25375 23103
rect 26252 23100 26280 23140
rect 26329 23137 26341 23140
rect 26375 23168 26387 23171
rect 26602 23168 26608 23180
rect 26375 23140 26608 23168
rect 26375 23137 26387 23140
rect 26329 23131 26387 23137
rect 26602 23128 26608 23140
rect 26660 23128 26666 23180
rect 26694 23128 26700 23180
rect 26752 23128 26758 23180
rect 26789 23171 26847 23177
rect 26789 23137 26801 23171
rect 26835 23168 26847 23171
rect 26878 23168 26884 23180
rect 26835 23140 26884 23168
rect 26835 23137 26847 23140
rect 26789 23131 26847 23137
rect 26804 23100 26832 23131
rect 26878 23128 26884 23140
rect 26936 23168 26942 23180
rect 27448 23177 27476 23208
rect 27249 23171 27307 23177
rect 27249 23168 27261 23171
rect 26936 23140 27261 23168
rect 26936 23128 26942 23140
rect 27249 23137 27261 23140
rect 27295 23137 27307 23171
rect 27249 23131 27307 23137
rect 27433 23171 27491 23177
rect 27433 23137 27445 23171
rect 27479 23137 27491 23171
rect 27433 23131 27491 23137
rect 25317 23063 25375 23069
rect 25792 23072 26280 23100
rect 26344 23072 26832 23100
rect 27448 23100 27476 23131
rect 27522 23100 27528 23112
rect 27448 23072 27528 23100
rect 25792 23032 25820 23072
rect 26344 23044 26372 23072
rect 27522 23060 27528 23072
rect 27580 23060 27586 23112
rect 27632 23109 27660 23276
rect 30374 23264 30380 23316
rect 30432 23264 30438 23316
rect 29914 23196 29920 23248
rect 29972 23196 29978 23248
rect 28258 23128 28264 23180
rect 28316 23168 28322 23180
rect 28629 23171 28687 23177
rect 28629 23168 28641 23171
rect 28316 23140 28641 23168
rect 28316 23128 28322 23140
rect 28629 23137 28641 23140
rect 28675 23137 28687 23171
rect 28629 23131 28687 23137
rect 31294 23128 31300 23180
rect 31352 23128 31358 23180
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23069 27675 23103
rect 27617 23063 27675 23069
rect 24872 23004 25820 23032
rect 25869 23035 25927 23041
rect 25869 23001 25881 23035
rect 25915 23032 25927 23035
rect 25958 23032 25964 23044
rect 25915 23004 25964 23032
rect 25915 23001 25927 23004
rect 25869 22995 25927 23001
rect 25958 22992 25964 23004
rect 26016 22992 26022 23044
rect 26234 22992 26240 23044
rect 26292 22992 26298 23044
rect 26326 22992 26332 23044
rect 26384 22992 26390 23044
rect 26786 22992 26792 23044
rect 26844 23032 26850 23044
rect 28276 23032 28304 23128
rect 28902 23060 28908 23112
rect 28960 23060 28966 23112
rect 30282 23060 30288 23112
rect 30340 23100 30346 23112
rect 30653 23103 30711 23109
rect 30653 23100 30665 23103
rect 30340 23072 30665 23100
rect 30340 23060 30346 23072
rect 30653 23069 30665 23072
rect 30699 23069 30711 23103
rect 30653 23063 30711 23069
rect 26844 23004 28304 23032
rect 26844 22992 26850 23004
rect 5626 22924 5632 22976
rect 5684 22924 5690 22976
rect 7190 22924 7196 22976
rect 7248 22924 7254 22976
rect 7650 22924 7656 22976
rect 7708 22964 7714 22976
rect 8021 22967 8079 22973
rect 8021 22964 8033 22967
rect 7708 22936 8033 22964
rect 7708 22924 7714 22936
rect 8021 22933 8033 22936
rect 8067 22933 8079 22967
rect 8021 22927 8079 22933
rect 13538 22924 13544 22976
rect 13596 22964 13602 22976
rect 14001 22967 14059 22973
rect 14001 22964 14013 22967
rect 13596 22936 14013 22964
rect 13596 22924 13602 22936
rect 14001 22933 14013 22936
rect 14047 22933 14059 22967
rect 14001 22927 14059 22933
rect 14274 22924 14280 22976
rect 14332 22964 14338 22976
rect 14826 22964 14832 22976
rect 14332 22936 14832 22964
rect 14332 22924 14338 22936
rect 14826 22924 14832 22936
rect 14884 22924 14890 22976
rect 15378 22924 15384 22976
rect 15436 22964 15442 22976
rect 18874 22964 18880 22976
rect 15436 22936 18880 22964
rect 15436 22924 15442 22936
rect 18874 22924 18880 22936
rect 18932 22924 18938 22976
rect 21358 22924 21364 22976
rect 21416 22924 21422 22976
rect 23198 22924 23204 22976
rect 23256 22964 23262 22976
rect 23477 22967 23535 22973
rect 23477 22964 23489 22967
rect 23256 22936 23489 22964
rect 23256 22924 23262 22936
rect 23477 22933 23489 22936
rect 23523 22933 23535 22967
rect 23477 22927 23535 22933
rect 24397 22967 24455 22973
rect 24397 22933 24409 22967
rect 24443 22964 24455 22967
rect 24854 22964 24860 22976
rect 24443 22936 24860 22964
rect 24443 22933 24455 22936
rect 24397 22927 24455 22933
rect 24854 22924 24860 22936
rect 24912 22924 24918 22976
rect 25041 22967 25099 22973
rect 25041 22933 25053 22967
rect 25087 22964 25099 22967
rect 25774 22964 25780 22976
rect 25087 22936 25780 22964
rect 25087 22933 25099 22936
rect 25041 22927 25099 22933
rect 25774 22924 25780 22936
rect 25832 22924 25838 22976
rect 28718 22924 28724 22976
rect 28776 22964 28782 22976
rect 31294 22964 31300 22976
rect 28776 22936 31300 22964
rect 28776 22924 28782 22936
rect 31294 22924 31300 22936
rect 31352 22924 31358 22976
rect 2760 22874 32200 22896
rect 2760 22822 6286 22874
rect 6338 22822 6350 22874
rect 6402 22822 6414 22874
rect 6466 22822 6478 22874
rect 6530 22822 6542 22874
rect 6594 22822 13646 22874
rect 13698 22822 13710 22874
rect 13762 22822 13774 22874
rect 13826 22822 13838 22874
rect 13890 22822 13902 22874
rect 13954 22822 21006 22874
rect 21058 22822 21070 22874
rect 21122 22822 21134 22874
rect 21186 22822 21198 22874
rect 21250 22822 21262 22874
rect 21314 22822 28366 22874
rect 28418 22822 28430 22874
rect 28482 22822 28494 22874
rect 28546 22822 28558 22874
rect 28610 22822 28622 22874
rect 28674 22822 32200 22874
rect 2760 22800 32200 22822
rect 4982 22720 4988 22772
rect 5040 22760 5046 22772
rect 5077 22763 5135 22769
rect 5077 22760 5089 22763
rect 5040 22732 5089 22760
rect 5040 22720 5046 22732
rect 5077 22729 5089 22732
rect 5123 22729 5135 22763
rect 5077 22723 5135 22729
rect 5718 22720 5724 22772
rect 5776 22760 5782 22772
rect 5776 22732 7052 22760
rect 5776 22720 5782 22732
rect 5192 22596 6408 22624
rect 5192 22568 5220 22596
rect 4433 22559 4491 22565
rect 4433 22525 4445 22559
rect 4479 22525 4491 22559
rect 4433 22519 4491 22525
rect 1302 22448 1308 22500
rect 1360 22488 1366 22500
rect 3237 22491 3295 22497
rect 3237 22488 3249 22491
rect 1360 22460 3249 22488
rect 1360 22448 1366 22460
rect 3237 22457 3249 22460
rect 3283 22457 3295 22491
rect 4448 22488 4476 22519
rect 5166 22516 5172 22568
rect 5224 22516 5230 22568
rect 6086 22516 6092 22568
rect 6144 22516 6150 22568
rect 6380 22565 6408 22596
rect 6365 22559 6423 22565
rect 6365 22525 6377 22559
rect 6411 22556 6423 22559
rect 7024 22556 7052 22732
rect 7190 22720 7196 22772
rect 7248 22760 7254 22772
rect 7634 22763 7692 22769
rect 7634 22760 7646 22763
rect 7248 22732 7646 22760
rect 7248 22720 7254 22732
rect 7634 22729 7646 22732
rect 7680 22729 7692 22763
rect 7634 22723 7692 22729
rect 8662 22720 8668 22772
rect 8720 22760 8726 22772
rect 9125 22763 9183 22769
rect 9125 22760 9137 22763
rect 8720 22732 9137 22760
rect 8720 22720 8726 22732
rect 9125 22729 9137 22732
rect 9171 22729 9183 22763
rect 9125 22723 9183 22729
rect 14182 22720 14188 22772
rect 14240 22760 14246 22772
rect 14277 22763 14335 22769
rect 14277 22760 14289 22763
rect 14240 22732 14289 22760
rect 14240 22720 14246 22732
rect 14277 22729 14289 22732
rect 14323 22729 14335 22763
rect 14277 22723 14335 22729
rect 14458 22720 14464 22772
rect 14516 22720 14522 22772
rect 14734 22720 14740 22772
rect 14792 22720 14798 22772
rect 14936 22732 15148 22760
rect 14366 22652 14372 22704
rect 14424 22692 14430 22704
rect 14936 22692 14964 22732
rect 14424 22664 14964 22692
rect 14424 22652 14430 22664
rect 15010 22652 15016 22704
rect 15068 22652 15074 22704
rect 7098 22584 7104 22636
rect 7156 22584 7162 22636
rect 8386 22624 8392 22636
rect 7392 22596 8392 22624
rect 7392 22565 7420 22596
rect 8386 22584 8392 22596
rect 8444 22584 8450 22636
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 12529 22627 12587 22633
rect 12529 22624 12541 22627
rect 12492 22596 12541 22624
rect 12492 22584 12498 22596
rect 12529 22593 12541 22596
rect 12575 22593 12587 22627
rect 15028 22624 15056 22652
rect 12529 22587 12587 22593
rect 12636 22596 15056 22624
rect 7377 22559 7435 22565
rect 7377 22556 7389 22559
rect 6411 22528 6868 22556
rect 7024 22528 7389 22556
rect 6411 22525 6423 22528
rect 6365 22519 6423 22525
rect 6638 22488 6644 22500
rect 4448 22460 6644 22488
rect 3237 22451 3295 22457
rect 6638 22448 6644 22460
rect 6696 22448 6702 22500
rect 6840 22432 6868 22528
rect 7377 22525 7389 22528
rect 7423 22525 7435 22559
rect 7377 22519 7435 22525
rect 9766 22516 9772 22568
rect 9824 22516 9830 22568
rect 10137 22559 10195 22565
rect 10137 22525 10149 22559
rect 10183 22556 10195 22559
rect 10689 22559 10747 22565
rect 10689 22556 10701 22559
rect 10183 22528 10701 22556
rect 10183 22525 10195 22528
rect 10137 22519 10195 22525
rect 10689 22525 10701 22528
rect 10735 22525 10747 22559
rect 10689 22519 10747 22525
rect 6917 22491 6975 22497
rect 6917 22457 6929 22491
rect 6963 22488 6975 22491
rect 10045 22491 10103 22497
rect 10045 22488 10057 22491
rect 6963 22460 8064 22488
rect 8878 22460 10057 22488
rect 6963 22457 6975 22460
rect 6917 22451 6975 22457
rect 5442 22380 5448 22432
rect 5500 22380 5506 22432
rect 6270 22380 6276 22432
rect 6328 22380 6334 22432
rect 6546 22380 6552 22432
rect 6604 22380 6610 22432
rect 6822 22380 6828 22432
rect 6880 22380 6886 22432
rect 7009 22423 7067 22429
rect 7009 22389 7021 22423
rect 7055 22420 7067 22423
rect 7650 22420 7656 22432
rect 7055 22392 7656 22420
rect 7055 22389 7067 22392
rect 7009 22383 7067 22389
rect 7650 22380 7656 22392
rect 7708 22380 7714 22432
rect 8036 22420 8064 22460
rect 10045 22457 10057 22460
rect 10091 22457 10103 22491
rect 10045 22451 10103 22457
rect 10152 22432 10180 22519
rect 11606 22516 11612 22568
rect 11664 22516 11670 22568
rect 11698 22516 11704 22568
rect 11756 22556 11762 22568
rect 12636 22556 12664 22596
rect 11756 22528 12664 22556
rect 11756 22516 11762 22528
rect 12802 22516 12808 22568
rect 12860 22516 12866 22568
rect 13354 22516 13360 22568
rect 13412 22556 13418 22568
rect 14093 22559 14151 22565
rect 14093 22556 14105 22559
rect 13412 22528 14105 22556
rect 13412 22516 13418 22528
rect 14093 22525 14105 22528
rect 14139 22525 14151 22559
rect 14461 22559 14519 22565
rect 14461 22556 14473 22559
rect 14093 22519 14151 22525
rect 14200 22528 14473 22556
rect 12437 22491 12495 22497
rect 12437 22457 12449 22491
rect 12483 22488 12495 22491
rect 12618 22488 12624 22500
rect 12483 22460 12624 22488
rect 12483 22457 12495 22460
rect 12437 22451 12495 22457
rect 12618 22448 12624 22460
rect 12676 22488 12682 22500
rect 13541 22491 13599 22497
rect 13541 22488 13553 22491
rect 12676 22460 13553 22488
rect 12676 22448 12682 22460
rect 13541 22457 13553 22460
rect 13587 22457 13599 22491
rect 13541 22451 13599 22457
rect 14200 22432 14228 22528
rect 14461 22525 14473 22528
rect 14507 22525 14519 22559
rect 14461 22519 14519 22525
rect 14550 22516 14556 22568
rect 14608 22516 14614 22568
rect 14660 22565 14688 22596
rect 15120 22568 15148 22732
rect 15304 22732 15976 22760
rect 14645 22559 14703 22565
rect 14645 22525 14657 22559
rect 14691 22525 14703 22559
rect 14645 22519 14703 22525
rect 14734 22516 14740 22568
rect 14792 22516 14798 22568
rect 14921 22559 14979 22565
rect 14921 22525 14933 22559
rect 14967 22525 14979 22559
rect 14921 22519 14979 22525
rect 15013 22559 15071 22565
rect 15013 22525 15025 22559
rect 15059 22556 15071 22559
rect 15102 22556 15108 22568
rect 15059 22528 15108 22556
rect 15059 22525 15071 22528
rect 15013 22519 15071 22525
rect 14568 22488 14596 22516
rect 14936 22488 14964 22519
rect 15102 22516 15108 22528
rect 15160 22516 15166 22568
rect 15304 22565 15332 22732
rect 15565 22695 15623 22701
rect 15565 22661 15577 22695
rect 15611 22661 15623 22695
rect 15565 22655 15623 22661
rect 15580 22624 15608 22655
rect 15838 22652 15844 22704
rect 15896 22652 15902 22704
rect 15948 22692 15976 22732
rect 16114 22720 16120 22772
rect 16172 22760 16178 22772
rect 16669 22763 16727 22769
rect 16669 22760 16681 22763
rect 16172 22732 16681 22760
rect 16172 22720 16178 22732
rect 16669 22729 16681 22732
rect 16715 22729 16727 22763
rect 16669 22723 16727 22729
rect 17034 22720 17040 22772
rect 17092 22760 17098 22772
rect 17092 22732 19012 22760
rect 17092 22720 17098 22732
rect 17052 22692 17080 22720
rect 15948 22664 17080 22692
rect 18877 22695 18935 22701
rect 18877 22661 18889 22695
rect 18923 22661 18935 22695
rect 18877 22655 18935 22661
rect 16025 22627 16083 22633
rect 16025 22624 16037 22627
rect 15580 22596 16037 22624
rect 16025 22593 16037 22596
rect 16071 22593 16083 22627
rect 16945 22627 17003 22633
rect 16945 22624 16957 22627
rect 16025 22587 16083 22593
rect 16546 22596 16957 22624
rect 15289 22559 15347 22565
rect 15289 22525 15301 22559
rect 15335 22525 15347 22559
rect 15289 22519 15347 22525
rect 15381 22559 15439 22565
rect 15381 22525 15393 22559
rect 15427 22556 15439 22559
rect 15562 22556 15568 22568
rect 15427 22528 15568 22556
rect 15427 22525 15439 22528
rect 15381 22519 15439 22525
rect 15562 22516 15568 22528
rect 15620 22516 15626 22568
rect 15749 22559 15807 22565
rect 15749 22525 15761 22559
rect 15795 22525 15807 22559
rect 15749 22519 15807 22525
rect 14568 22460 14964 22488
rect 15197 22491 15255 22497
rect 15197 22457 15209 22491
rect 15243 22488 15255 22491
rect 15470 22488 15476 22500
rect 15243 22460 15476 22488
rect 15243 22457 15255 22460
rect 15197 22451 15255 22457
rect 15470 22448 15476 22460
rect 15528 22448 15534 22500
rect 9217 22423 9275 22429
rect 9217 22420 9229 22423
rect 8036 22392 9229 22420
rect 9217 22389 9229 22392
rect 9263 22389 9275 22423
rect 9217 22383 9275 22389
rect 10134 22380 10140 22432
rect 10192 22380 10198 22432
rect 10778 22380 10784 22432
rect 10836 22380 10842 22432
rect 11054 22380 11060 22432
rect 11112 22380 11118 22432
rect 11974 22380 11980 22432
rect 12032 22380 12038 22432
rect 12345 22423 12403 22429
rect 12345 22389 12357 22423
rect 12391 22420 12403 22423
rect 12526 22420 12532 22432
rect 12391 22392 12532 22420
rect 12391 22389 12403 22392
rect 12345 22383 12403 22389
rect 12526 22380 12532 22392
rect 12584 22420 12590 22432
rect 13262 22420 13268 22432
rect 12584 22392 13268 22420
rect 12584 22380 12590 22392
rect 13262 22380 13268 22392
rect 13320 22380 13326 22432
rect 13446 22380 13452 22432
rect 13504 22380 13510 22432
rect 14182 22380 14188 22432
rect 14240 22380 14246 22432
rect 14642 22380 14648 22432
rect 14700 22420 14706 22432
rect 15764 22420 15792 22519
rect 14700 22392 15792 22420
rect 14700 22380 14706 22392
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16546 22420 16574 22596
rect 16945 22593 16957 22596
rect 16991 22593 17003 22627
rect 16945 22587 17003 22593
rect 17221 22627 17279 22633
rect 17221 22593 17233 22627
rect 17267 22624 17279 22627
rect 18892 22624 18920 22655
rect 17267 22596 18920 22624
rect 18984 22624 19012 22732
rect 20898 22720 20904 22772
rect 20956 22720 20962 22772
rect 21358 22720 21364 22772
rect 21416 22720 21422 22772
rect 22186 22720 22192 22772
rect 22244 22760 22250 22772
rect 22373 22763 22431 22769
rect 22373 22760 22385 22763
rect 22244 22732 22385 22760
rect 22244 22720 22250 22732
rect 22373 22729 22385 22732
rect 22419 22729 22431 22763
rect 22373 22723 22431 22729
rect 22820 22763 22878 22769
rect 22820 22729 22832 22763
rect 22866 22760 22878 22763
rect 23198 22760 23204 22772
rect 22866 22732 23204 22760
rect 22866 22729 22878 22732
rect 22820 22723 22878 22729
rect 23198 22720 23204 22732
rect 23256 22720 23262 22772
rect 24302 22720 24308 22772
rect 24360 22720 24366 22772
rect 24670 22720 24676 22772
rect 24728 22720 24734 22772
rect 26050 22720 26056 22772
rect 26108 22760 26114 22772
rect 27617 22763 27675 22769
rect 27617 22760 27629 22763
rect 26108 22732 27629 22760
rect 26108 22720 26114 22732
rect 27617 22729 27629 22732
rect 27663 22729 27675 22763
rect 27617 22723 27675 22729
rect 28721 22763 28779 22769
rect 28721 22729 28733 22763
rect 28767 22760 28779 22763
rect 28902 22760 28908 22772
rect 28767 22732 28908 22760
rect 28767 22729 28779 22732
rect 28721 22723 28779 22729
rect 28902 22720 28908 22732
rect 28960 22720 28966 22772
rect 29089 22763 29147 22769
rect 29089 22729 29101 22763
rect 29135 22760 29147 22763
rect 29362 22760 29368 22772
rect 29135 22732 29368 22760
rect 29135 22729 29147 22732
rect 29089 22723 29147 22729
rect 29362 22720 29368 22732
rect 29420 22720 29426 22772
rect 29825 22763 29883 22769
rect 29825 22729 29837 22763
rect 29871 22760 29883 22763
rect 29914 22760 29920 22772
rect 29871 22732 29920 22760
rect 29871 22729 29883 22732
rect 29825 22723 29883 22729
rect 29914 22720 29920 22732
rect 29972 22720 29978 22772
rect 19150 22652 19156 22704
rect 19208 22692 19214 22704
rect 19208 22664 19472 22692
rect 19208 22652 19214 22664
rect 19444 22633 19472 22664
rect 19337 22627 19395 22633
rect 19337 22624 19349 22627
rect 18984 22596 19349 22624
rect 17267 22593 17279 22596
rect 17221 22587 17279 22593
rect 19337 22593 19349 22596
rect 19383 22593 19395 22627
rect 19337 22587 19395 22593
rect 19429 22627 19487 22633
rect 19429 22593 19441 22627
rect 19475 22593 19487 22627
rect 19429 22587 19487 22593
rect 19058 22516 19064 22568
rect 19116 22556 19122 22568
rect 19245 22559 19303 22565
rect 19245 22556 19257 22559
rect 19116 22528 19257 22556
rect 19116 22516 19122 22528
rect 19245 22525 19257 22528
rect 19291 22525 19303 22559
rect 19245 22519 19303 22525
rect 19889 22559 19947 22565
rect 19889 22525 19901 22559
rect 19935 22556 19947 22559
rect 20530 22556 20536 22568
rect 19935 22528 20536 22556
rect 19935 22525 19947 22528
rect 19889 22519 19947 22525
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 20714 22516 20720 22568
rect 20772 22516 20778 22568
rect 21376 22556 21404 22720
rect 21634 22692 21640 22704
rect 21468 22664 21640 22692
rect 21468 22636 21496 22664
rect 21634 22652 21640 22664
rect 21692 22652 21698 22704
rect 24688 22692 24716 22720
rect 27890 22692 27896 22704
rect 24688 22664 25636 22692
rect 21450 22584 21456 22636
rect 21508 22584 21514 22636
rect 21729 22559 21787 22565
rect 21729 22556 21741 22559
rect 21376 22528 21741 22556
rect 21729 22525 21741 22528
rect 21775 22525 21787 22559
rect 21729 22519 21787 22525
rect 22094 22516 22100 22568
rect 22152 22556 22158 22568
rect 22557 22559 22615 22565
rect 22557 22556 22569 22559
rect 22152 22528 22569 22556
rect 22152 22516 22158 22528
rect 22557 22525 22569 22528
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 24394 22516 24400 22568
rect 24452 22516 24458 22568
rect 25406 22565 25412 22568
rect 25404 22556 25412 22565
rect 25367 22528 25412 22556
rect 25404 22519 25412 22528
rect 25406 22516 25412 22519
rect 25464 22516 25470 22568
rect 25501 22559 25559 22565
rect 25501 22525 25513 22559
rect 25547 22556 25559 22559
rect 25608 22556 25636 22664
rect 25838 22664 27896 22692
rect 25838 22624 25866 22664
rect 27890 22652 27896 22664
rect 27948 22652 27954 22704
rect 28810 22652 28816 22704
rect 28868 22692 28874 22704
rect 29457 22695 29515 22701
rect 28868 22664 28994 22692
rect 28868 22652 28874 22664
rect 28169 22627 28227 22633
rect 28169 22624 28181 22627
rect 25792 22596 25866 22624
rect 26068 22596 28181 22624
rect 25547 22528 25636 22556
rect 25547 22525 25559 22528
rect 25501 22519 25559 22525
rect 25682 22516 25688 22568
rect 25740 22516 25746 22568
rect 25792 22565 25820 22596
rect 26068 22568 26096 22596
rect 28169 22593 28181 22596
rect 28215 22593 28227 22627
rect 28966 22624 28994 22664
rect 29457 22661 29469 22695
rect 29503 22661 29515 22695
rect 29457 22655 29515 22661
rect 29181 22627 29239 22633
rect 29181 22624 29193 22627
rect 28966 22596 29193 22624
rect 28169 22587 28227 22593
rect 29181 22593 29193 22596
rect 29227 22624 29239 22627
rect 29472 22624 29500 22655
rect 30282 22624 30288 22636
rect 29227 22596 29500 22624
rect 29932 22596 30288 22624
rect 29227 22593 29239 22596
rect 29181 22587 29239 22593
rect 25776 22559 25834 22565
rect 25776 22525 25788 22559
rect 25822 22525 25834 22559
rect 25776 22519 25834 22525
rect 25869 22559 25927 22565
rect 25869 22525 25881 22559
rect 25915 22525 25927 22559
rect 25869 22519 25927 22525
rect 17954 22448 17960 22500
rect 18012 22448 18018 22500
rect 19334 22448 19340 22500
rect 19392 22488 19398 22500
rect 21269 22491 21327 22497
rect 19392 22460 20208 22488
rect 19392 22448 19398 22460
rect 15896 22392 16574 22420
rect 18693 22423 18751 22429
rect 15896 22380 15902 22392
rect 18693 22389 18705 22423
rect 18739 22420 18751 22423
rect 19702 22420 19708 22432
rect 18739 22392 19708 22420
rect 18739 22389 18751 22392
rect 18693 22383 18751 22389
rect 19702 22380 19708 22392
rect 19760 22380 19766 22432
rect 19794 22380 19800 22432
rect 19852 22380 19858 22432
rect 20070 22380 20076 22432
rect 20128 22380 20134 22432
rect 20180 22420 20208 22460
rect 21269 22457 21281 22491
rect 21315 22488 21327 22491
rect 22186 22488 22192 22500
rect 21315 22460 22192 22488
rect 21315 22457 21327 22460
rect 21269 22451 21327 22457
rect 22186 22448 22192 22460
rect 22244 22448 22250 22500
rect 23474 22448 23480 22500
rect 23532 22448 23538 22500
rect 25041 22491 25099 22497
rect 25041 22457 25053 22491
rect 25087 22488 25099 22491
rect 25593 22491 25651 22497
rect 25087 22460 25452 22488
rect 25087 22457 25099 22460
rect 25041 22451 25099 22457
rect 21358 22420 21364 22432
rect 20180 22392 21364 22420
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 25222 22380 25228 22432
rect 25280 22380 25286 22432
rect 25424 22420 25452 22460
rect 25593 22457 25605 22491
rect 25639 22488 25651 22491
rect 25700 22488 25728 22516
rect 25639 22460 25728 22488
rect 25884 22488 25912 22519
rect 26050 22516 26056 22568
rect 26108 22516 26114 22568
rect 26418 22516 26424 22568
rect 26476 22556 26482 22568
rect 26786 22556 26792 22568
rect 26476 22528 26792 22556
rect 26476 22516 26482 22528
rect 26786 22516 26792 22528
rect 26844 22516 26850 22568
rect 27065 22559 27123 22565
rect 27065 22525 27077 22559
rect 27111 22525 27123 22559
rect 27433 22559 27491 22565
rect 27433 22556 27445 22559
rect 27065 22519 27123 22525
rect 27172 22528 27445 22556
rect 26326 22488 26332 22500
rect 25884 22460 26332 22488
rect 25639 22457 25651 22460
rect 25593 22451 25651 22457
rect 26326 22448 26332 22460
rect 26384 22448 26390 22500
rect 27080 22420 27108 22519
rect 27172 22432 27200 22528
rect 27433 22525 27445 22528
rect 27479 22525 27491 22559
rect 27433 22519 27491 22525
rect 27522 22516 27528 22568
rect 27580 22516 27586 22568
rect 27614 22516 27620 22568
rect 27672 22516 27678 22568
rect 27706 22516 27712 22568
rect 27764 22516 27770 22568
rect 27890 22516 27896 22568
rect 27948 22516 27954 22568
rect 28905 22559 28963 22565
rect 28905 22525 28917 22559
rect 28951 22525 28963 22559
rect 28905 22519 28963 22525
rect 29273 22559 29331 22565
rect 29273 22525 29285 22559
rect 29319 22556 29331 22559
rect 29454 22556 29460 22568
rect 29319 22528 29460 22556
rect 29319 22525 29331 22528
rect 29273 22519 29331 22525
rect 27540 22488 27568 22516
rect 28920 22488 28948 22519
rect 29454 22516 29460 22528
rect 29512 22516 29518 22568
rect 29932 22565 29960 22596
rect 30282 22584 30288 22596
rect 30340 22584 30346 22636
rect 29917 22559 29975 22565
rect 29917 22525 29929 22559
rect 29963 22525 29975 22559
rect 29917 22519 29975 22525
rect 29730 22488 29736 22500
rect 27540 22460 29736 22488
rect 29730 22448 29736 22460
rect 29788 22448 29794 22500
rect 25424 22392 27108 22420
rect 27154 22380 27160 22432
rect 27212 22380 27218 22432
rect 27246 22380 27252 22432
rect 27304 22420 27310 22432
rect 27522 22420 27528 22432
rect 27304 22392 27528 22420
rect 27304 22380 27310 22392
rect 27522 22380 27528 22392
rect 27580 22380 27586 22432
rect 27798 22380 27804 22432
rect 27856 22380 27862 22432
rect 2760 22330 32200 22352
rect 2760 22278 6946 22330
rect 6998 22278 7010 22330
rect 7062 22278 7074 22330
rect 7126 22278 7138 22330
rect 7190 22278 7202 22330
rect 7254 22278 14306 22330
rect 14358 22278 14370 22330
rect 14422 22278 14434 22330
rect 14486 22278 14498 22330
rect 14550 22278 14562 22330
rect 14614 22278 21666 22330
rect 21718 22278 21730 22330
rect 21782 22278 21794 22330
rect 21846 22278 21858 22330
rect 21910 22278 21922 22330
rect 21974 22278 29026 22330
rect 29078 22278 29090 22330
rect 29142 22278 29154 22330
rect 29206 22278 29218 22330
rect 29270 22278 29282 22330
rect 29334 22278 32200 22330
rect 2760 22256 32200 22278
rect 5442 22216 5448 22228
rect 4540 22188 5448 22216
rect 4540 22157 4568 22188
rect 5442 22176 5448 22188
rect 5500 22176 5506 22228
rect 6270 22176 6276 22228
rect 6328 22176 6334 22228
rect 6546 22216 6552 22228
rect 6380 22188 6552 22216
rect 4525 22151 4583 22157
rect 4525 22117 4537 22151
rect 4571 22117 4583 22151
rect 6288 22148 6316 22176
rect 6380 22157 6408 22188
rect 6546 22176 6552 22188
rect 6604 22176 6610 22228
rect 6638 22176 6644 22228
rect 6696 22216 6702 22228
rect 7837 22219 7895 22225
rect 7837 22216 7849 22219
rect 6696 22188 7849 22216
rect 6696 22176 6702 22188
rect 7837 22185 7849 22188
rect 7883 22216 7895 22219
rect 9766 22216 9772 22228
rect 7883 22188 9772 22216
rect 7883 22185 7895 22188
rect 7837 22179 7895 22185
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 10410 22176 10416 22228
rect 10468 22216 10474 22228
rect 10505 22219 10563 22225
rect 10505 22216 10517 22219
rect 10468 22188 10517 22216
rect 10468 22176 10474 22188
rect 10505 22185 10517 22188
rect 10551 22185 10563 22219
rect 10505 22179 10563 22185
rect 11054 22176 11060 22228
rect 11112 22176 11118 22228
rect 11974 22216 11980 22228
rect 11256 22188 11980 22216
rect 5750 22120 6316 22148
rect 6365 22151 6423 22157
rect 4525 22111 4583 22117
rect 6365 22117 6377 22151
rect 6411 22117 6423 22151
rect 11072 22148 11100 22176
rect 11256 22157 11284 22188
rect 11974 22176 11980 22188
rect 12032 22176 12038 22228
rect 12713 22219 12771 22225
rect 12713 22185 12725 22219
rect 12759 22216 12771 22219
rect 13354 22216 13360 22228
rect 12759 22188 13360 22216
rect 12759 22185 12771 22188
rect 12713 22179 12771 22185
rect 13354 22176 13360 22188
rect 13412 22176 13418 22228
rect 13446 22176 13452 22228
rect 13504 22176 13510 22228
rect 13538 22176 13544 22228
rect 13596 22216 13602 22228
rect 13596 22188 15332 22216
rect 13596 22176 13602 22188
rect 6365 22111 6423 22117
rect 10980 22120 11100 22148
rect 11241 22151 11299 22157
rect 7466 22040 7472 22092
rect 7524 22040 7530 22092
rect 8665 22083 8723 22089
rect 8665 22080 8677 22083
rect 7576 22052 8677 22080
rect 3234 21972 3240 22024
rect 3292 22012 3298 22024
rect 3513 22015 3571 22021
rect 3513 22012 3525 22015
rect 3292 21984 3525 22012
rect 3292 21972 3298 21984
rect 3513 21981 3525 21984
rect 3559 21981 3571 22015
rect 3513 21975 3571 21981
rect 4249 22015 4307 22021
rect 4249 21981 4261 22015
rect 4295 22012 4307 22015
rect 6086 22012 6092 22024
rect 4295 21984 6092 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 6086 21972 6092 21984
rect 6144 21972 6150 22024
rect 6454 21972 6460 22024
rect 6512 22012 6518 22024
rect 7576 22012 7604 22052
rect 8665 22049 8677 22052
rect 8711 22080 8723 22083
rect 9033 22083 9091 22089
rect 9033 22080 9045 22083
rect 8711 22052 9045 22080
rect 8711 22049 8723 22052
rect 8665 22043 8723 22049
rect 9033 22049 9045 22052
rect 9079 22049 9091 22083
rect 9033 22043 9091 22049
rect 10045 22083 10103 22089
rect 10045 22049 10057 22083
rect 10091 22049 10103 22083
rect 10045 22043 10103 22049
rect 10597 22083 10655 22089
rect 10597 22049 10609 22083
rect 10643 22080 10655 22083
rect 10980 22080 11008 22120
rect 11241 22117 11253 22151
rect 11287 22117 11299 22151
rect 11241 22111 11299 22117
rect 11790 22108 11796 22160
rect 11848 22108 11854 22160
rect 14642 22148 14648 22160
rect 13832 22120 14648 22148
rect 10643 22052 11008 22080
rect 12989 22083 13047 22089
rect 10643 22049 10655 22052
rect 10597 22043 10655 22049
rect 12989 22049 13001 22083
rect 13035 22080 13047 22083
rect 13832 22080 13860 22120
rect 14642 22108 14648 22120
rect 14700 22108 14706 22160
rect 14918 22080 14924 22092
rect 13035 22052 13860 22080
rect 14476 22052 14924 22080
rect 13035 22049 13047 22052
rect 12989 22043 13047 22049
rect 8110 22012 8116 22024
rect 6512 21984 7604 22012
rect 7668 21984 8116 22012
rect 6512 21972 6518 21984
rect 4154 21836 4160 21888
rect 4212 21836 4218 21888
rect 5994 21836 6000 21888
rect 6052 21836 6058 21888
rect 7098 21836 7104 21888
rect 7156 21876 7162 21888
rect 7668 21876 7696 21984
rect 8110 21972 8116 21984
rect 8168 21972 8174 22024
rect 8202 21972 8208 22024
rect 8260 22012 8266 22024
rect 8297 22015 8355 22021
rect 8297 22012 8309 22015
rect 8260 21984 8309 22012
rect 8260 21972 8266 21984
rect 8297 21981 8309 21984
rect 8343 21981 8355 22015
rect 8297 21975 8355 21981
rect 8478 21972 8484 22024
rect 8536 22012 8542 22024
rect 10060 22012 10088 22043
rect 10226 22012 10232 22024
rect 8536 21984 10232 22012
rect 8536 21972 8542 21984
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 22012 10839 22015
rect 10870 22012 10876 22024
rect 10827 21984 10876 22012
rect 10827 21981 10839 21984
rect 10781 21975 10839 21981
rect 10870 21972 10876 21984
rect 10928 21972 10934 22024
rect 10965 22015 11023 22021
rect 10965 21981 10977 22015
rect 11011 21981 11023 22015
rect 10965 21975 11023 21981
rect 9582 21904 9588 21956
rect 9640 21944 9646 21956
rect 10980 21944 11008 21975
rect 11974 21972 11980 22024
rect 12032 22012 12038 22024
rect 13004 22012 13032 22043
rect 12032 21984 13032 22012
rect 13357 22015 13415 22021
rect 12032 21972 12038 21984
rect 13357 21981 13369 22015
rect 13403 22012 13415 22015
rect 14476 22012 14504 22052
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 15013 22083 15071 22089
rect 15013 22049 15025 22083
rect 15059 22080 15071 22083
rect 15194 22080 15200 22092
rect 15059 22052 15200 22080
rect 15059 22049 15071 22052
rect 15013 22043 15071 22049
rect 15194 22040 15200 22052
rect 15252 22040 15258 22092
rect 15304 22089 15332 22188
rect 15562 22176 15568 22228
rect 15620 22216 15626 22228
rect 16482 22216 16488 22228
rect 15620 22188 16488 22216
rect 15620 22176 15626 22188
rect 16482 22176 16488 22188
rect 16540 22176 16546 22228
rect 17954 22176 17960 22228
rect 18012 22176 18018 22228
rect 20070 22176 20076 22228
rect 20128 22176 20134 22228
rect 21358 22176 21364 22228
rect 21416 22216 21422 22228
rect 21637 22219 21695 22225
rect 21637 22216 21649 22219
rect 21416 22188 21649 22216
rect 21416 22176 21422 22188
rect 21637 22185 21649 22188
rect 21683 22185 21695 22219
rect 21637 22179 21695 22185
rect 23661 22219 23719 22225
rect 23661 22185 23673 22219
rect 23707 22216 23719 22219
rect 24026 22216 24032 22228
rect 23707 22188 24032 22216
rect 23707 22185 23719 22188
rect 23661 22179 23719 22185
rect 24026 22176 24032 22188
rect 24084 22176 24090 22228
rect 24210 22176 24216 22228
rect 24268 22216 24274 22228
rect 24305 22219 24363 22225
rect 24305 22216 24317 22219
rect 24268 22188 24317 22216
rect 24268 22176 24274 22188
rect 24305 22185 24317 22188
rect 24351 22185 24363 22219
rect 24305 22179 24363 22185
rect 25041 22219 25099 22225
rect 25041 22185 25053 22219
rect 25087 22216 25099 22219
rect 25406 22216 25412 22228
rect 25087 22188 25412 22216
rect 25087 22185 25099 22188
rect 25041 22179 25099 22185
rect 25406 22176 25412 22188
rect 25464 22176 25470 22228
rect 27249 22219 27307 22225
rect 25516 22188 26004 22216
rect 18230 22148 18236 22160
rect 17342 22120 18236 22148
rect 18230 22108 18236 22120
rect 18288 22108 18294 22160
rect 19794 22108 19800 22160
rect 19852 22108 19858 22160
rect 20088 22148 20116 22176
rect 20257 22151 20315 22157
rect 20257 22148 20269 22151
rect 20088 22120 20269 22148
rect 20257 22117 20269 22120
rect 20303 22117 20315 22151
rect 20257 22111 20315 22117
rect 21542 22108 21548 22160
rect 21600 22148 21606 22160
rect 21729 22151 21787 22157
rect 21729 22148 21741 22151
rect 21600 22120 21741 22148
rect 21600 22108 21606 22120
rect 21729 22117 21741 22120
rect 21775 22117 21787 22151
rect 21729 22111 21787 22117
rect 22925 22151 22983 22157
rect 22925 22117 22937 22151
rect 22971 22148 22983 22151
rect 23566 22148 23572 22160
rect 22971 22120 23572 22148
rect 22971 22117 22983 22120
rect 22925 22111 22983 22117
rect 23566 22108 23572 22120
rect 23624 22148 23630 22160
rect 24578 22148 24584 22160
rect 23624 22120 24584 22148
rect 23624 22108 23630 22120
rect 24578 22108 24584 22120
rect 24636 22108 24642 22160
rect 24670 22108 24676 22160
rect 24728 22148 24734 22160
rect 25516 22157 25544 22188
rect 25291 22151 25349 22157
rect 25291 22148 25303 22151
rect 24728 22120 25303 22148
rect 24728 22108 24734 22120
rect 25291 22117 25303 22120
rect 25337 22117 25349 22151
rect 25291 22111 25349 22117
rect 25501 22151 25559 22157
rect 25501 22117 25513 22151
rect 25547 22117 25559 22151
rect 25501 22111 25559 22117
rect 15289 22083 15347 22089
rect 15289 22049 15301 22083
rect 15335 22080 15347 22083
rect 15378 22080 15384 22092
rect 15335 22052 15384 22080
rect 15335 22049 15347 22052
rect 15289 22043 15347 22049
rect 15378 22040 15384 22052
rect 15436 22040 15442 22092
rect 15841 22083 15899 22089
rect 15841 22080 15853 22083
rect 15764 22052 15853 22080
rect 13403 21984 14504 22012
rect 14553 22015 14611 22021
rect 13403 21981 13415 21984
rect 13357 21975 13415 21981
rect 14553 21981 14565 22015
rect 14599 21981 14611 22015
rect 14936 22012 14964 22040
rect 15764 22024 15792 22052
rect 15841 22049 15853 22052
rect 15887 22049 15899 22083
rect 15841 22043 15899 22049
rect 18049 22083 18107 22089
rect 18049 22049 18061 22083
rect 18095 22080 18107 22083
rect 23109 22083 23167 22089
rect 18095 22052 19104 22080
rect 18095 22049 18107 22052
rect 18049 22043 18107 22049
rect 15562 22012 15568 22024
rect 14936 21984 15568 22012
rect 14553 21975 14611 21981
rect 9640 21916 11008 21944
rect 13909 21947 13967 21953
rect 9640 21904 9646 21916
rect 13909 21913 13921 21947
rect 13955 21944 13967 21947
rect 14568 21944 14596 21975
rect 15562 21972 15568 21984
rect 15620 21972 15626 22024
rect 15746 21972 15752 22024
rect 15804 21972 15810 22024
rect 16114 21972 16120 22024
rect 16172 21972 16178 22024
rect 18782 21972 18788 22024
rect 18840 22012 18846 22024
rect 18966 22012 18972 22024
rect 18840 21984 18972 22012
rect 18840 21972 18846 21984
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 13955 21916 14596 21944
rect 13955 21913 13967 21916
rect 13909 21907 13967 21913
rect 14642 21904 14648 21956
rect 14700 21944 14706 21956
rect 18046 21944 18052 21956
rect 14700 21916 15976 21944
rect 14700 21904 14706 21916
rect 7156 21848 7696 21876
rect 7156 21836 7162 21848
rect 7926 21836 7932 21888
rect 7984 21876 7990 21888
rect 9674 21876 9680 21888
rect 7984 21848 9680 21876
rect 7984 21836 7990 21848
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 9950 21836 9956 21888
rect 10008 21836 10014 21888
rect 10042 21836 10048 21888
rect 10100 21876 10106 21888
rect 10137 21879 10195 21885
rect 10137 21876 10149 21879
rect 10100 21848 10149 21876
rect 10100 21836 10106 21848
rect 10137 21845 10149 21848
rect 10183 21845 10195 21879
rect 10137 21839 10195 21845
rect 12894 21836 12900 21888
rect 12952 21836 12958 21888
rect 13998 21836 14004 21888
rect 14056 21836 14062 21888
rect 14734 21836 14740 21888
rect 14792 21836 14798 21888
rect 14918 21836 14924 21888
rect 14976 21836 14982 21888
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 15565 21879 15623 21885
rect 15565 21876 15577 21879
rect 15344 21848 15577 21876
rect 15344 21836 15350 21848
rect 15565 21845 15577 21848
rect 15611 21845 15623 21879
rect 15948 21876 15976 21916
rect 17328 21916 18052 21944
rect 17328 21876 17356 21916
rect 18046 21904 18052 21916
rect 18104 21904 18110 21956
rect 18693 21947 18751 21953
rect 18693 21913 18705 21947
rect 18739 21944 18751 21947
rect 18739 21916 19012 21944
rect 18739 21913 18751 21916
rect 18693 21907 18751 21913
rect 18984 21888 19012 21916
rect 15948 21848 17356 21876
rect 17589 21879 17647 21885
rect 15565 21839 15623 21845
rect 17589 21845 17601 21879
rect 17635 21876 17647 21879
rect 17954 21876 17960 21888
rect 17635 21848 17960 21876
rect 17635 21845 17647 21848
rect 17589 21839 17647 21845
rect 17954 21836 17960 21848
rect 18012 21836 18018 21888
rect 18782 21836 18788 21888
rect 18840 21836 18846 21888
rect 18966 21836 18972 21888
rect 19024 21836 19030 21888
rect 19076 21876 19104 22052
rect 20548 22052 21772 22080
rect 19702 21972 19708 22024
rect 19760 22012 19766 22024
rect 20548 22021 20576 22052
rect 20533 22015 20591 22021
rect 19760 21984 20484 22012
rect 19760 21972 19766 21984
rect 20456 21944 20484 21984
rect 20533 21981 20545 22015
rect 20579 21981 20591 22015
rect 20533 21975 20591 21981
rect 20898 21972 20904 22024
rect 20956 22012 20962 22024
rect 21177 22015 21235 22021
rect 21177 22012 21189 22015
rect 20956 21984 21189 22012
rect 20956 21972 20962 21984
rect 21177 21981 21189 21984
rect 21223 21981 21235 22015
rect 21744 22012 21772 22052
rect 23109 22049 23121 22083
rect 23155 22080 23167 22083
rect 23934 22080 23940 22092
rect 23155 22052 23940 22080
rect 23155 22049 23167 22052
rect 23109 22043 23167 22049
rect 23934 22040 23940 22052
rect 23992 22040 23998 22092
rect 25406 22080 25412 22092
rect 24412 22052 25268 22080
rect 25367 22052 25412 22080
rect 22094 22012 22100 22024
rect 21744 21984 22100 22012
rect 21177 21975 21235 21981
rect 22094 21972 22100 21984
rect 22152 22012 22158 22024
rect 22465 22015 22523 22021
rect 22465 22012 22477 22015
rect 22152 21984 22477 22012
rect 22152 21972 22158 21984
rect 22465 21981 22477 21984
rect 22511 21981 22523 22015
rect 22465 21975 22523 21981
rect 23845 22015 23903 22021
rect 23845 21981 23857 22015
rect 23891 22012 23903 22015
rect 24412 22012 24440 22052
rect 25240 22024 25268 22052
rect 25406 22040 25412 22052
rect 25464 22040 25470 22092
rect 25593 22083 25651 22089
rect 25593 22049 25605 22083
rect 25639 22080 25651 22083
rect 25866 22080 25872 22092
rect 25639 22052 25872 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 25866 22040 25872 22052
rect 25924 22040 25930 22092
rect 25976 22080 26004 22188
rect 27249 22185 27261 22219
rect 27295 22216 27307 22219
rect 27798 22216 27804 22228
rect 27295 22188 27804 22216
rect 27295 22185 27307 22188
rect 27249 22179 27307 22185
rect 26694 22108 26700 22160
rect 26752 22148 26758 22160
rect 26789 22151 26847 22157
rect 26789 22148 26801 22151
rect 26752 22120 26801 22148
rect 26752 22108 26758 22120
rect 26789 22117 26801 22120
rect 26835 22117 26847 22151
rect 26789 22111 26847 22117
rect 27264 22080 27292 22179
rect 27798 22176 27804 22188
rect 27856 22176 27862 22228
rect 27338 22108 27344 22160
rect 27396 22108 27402 22160
rect 25976 22052 27292 22080
rect 23891 21984 24440 22012
rect 23891 21981 23903 21984
rect 23845 21975 23903 21981
rect 24486 21972 24492 22024
rect 24544 21972 24550 22024
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 25133 22015 25191 22021
rect 25133 22012 25145 22015
rect 24820 21984 25145 22012
rect 24820 21972 24826 21984
rect 25133 21981 25145 21984
rect 25179 21981 25191 22015
rect 25133 21975 25191 21981
rect 25222 21972 25228 22024
rect 25280 21972 25286 22024
rect 25976 22012 26004 22052
rect 27522 22040 27528 22092
rect 27580 22080 27586 22092
rect 27709 22083 27767 22089
rect 27709 22080 27721 22083
rect 27580 22052 27721 22080
rect 27580 22040 27586 22052
rect 27709 22049 27721 22052
rect 27755 22049 27767 22083
rect 27709 22043 27767 22049
rect 27982 22040 27988 22092
rect 28040 22040 28046 22092
rect 28074 22040 28080 22092
rect 28132 22080 28138 22092
rect 28169 22083 28227 22089
rect 28169 22080 28181 22083
rect 28132 22052 28181 22080
rect 28132 22040 28138 22052
rect 28169 22049 28181 22052
rect 28215 22049 28227 22083
rect 28169 22043 28227 22049
rect 30469 22083 30527 22089
rect 30469 22049 30481 22083
rect 30515 22049 30527 22083
rect 30469 22043 30527 22049
rect 25608 21984 26004 22012
rect 26053 22015 26111 22021
rect 20456 21916 25447 21944
rect 20070 21876 20076 21888
rect 19076 21848 20076 21876
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 20622 21836 20628 21888
rect 20680 21836 20686 21888
rect 23201 21879 23259 21885
rect 23201 21845 23213 21879
rect 23247 21876 23259 21879
rect 24670 21876 24676 21888
rect 23247 21848 24676 21876
rect 23247 21845 23259 21848
rect 23201 21839 23259 21845
rect 24670 21836 24676 21848
rect 24728 21836 24734 21888
rect 25419 21876 25447 21916
rect 25498 21904 25504 21956
rect 25556 21944 25562 21956
rect 25608 21944 25636 21984
rect 26053 21981 26065 22015
rect 26099 22012 26111 22015
rect 26326 22012 26332 22024
rect 26099 21984 26332 22012
rect 26099 21981 26111 21984
rect 26053 21975 26111 21981
rect 26326 21972 26332 21984
rect 26384 21972 26390 22024
rect 27430 21972 27436 22024
rect 27488 21972 27494 22024
rect 30484 21944 30512 22043
rect 31662 22040 31668 22092
rect 31720 22040 31726 22092
rect 25556 21916 25636 21944
rect 25700 21916 30512 21944
rect 25556 21904 25562 21916
rect 25700 21876 25728 21916
rect 25419 21848 25728 21876
rect 25774 21836 25780 21888
rect 25832 21836 25838 21888
rect 26050 21836 26056 21888
rect 26108 21876 26114 21888
rect 26694 21876 26700 21888
rect 26108 21848 26700 21876
rect 26108 21836 26114 21848
rect 26694 21836 26700 21848
rect 26752 21836 26758 21888
rect 26786 21836 26792 21888
rect 26844 21876 26850 21888
rect 26881 21879 26939 21885
rect 26881 21876 26893 21879
rect 26844 21848 26893 21876
rect 26844 21836 26850 21848
rect 26881 21845 26893 21848
rect 26927 21845 26939 21879
rect 26881 21839 26939 21845
rect 26970 21836 26976 21888
rect 27028 21876 27034 21888
rect 27801 21879 27859 21885
rect 27801 21876 27813 21879
rect 27028 21848 27813 21876
rect 27028 21836 27034 21848
rect 27801 21845 27813 21848
rect 27847 21845 27859 21879
rect 27801 21839 27859 21845
rect 2760 21786 32200 21808
rect 2760 21734 6286 21786
rect 6338 21734 6350 21786
rect 6402 21734 6414 21786
rect 6466 21734 6478 21786
rect 6530 21734 6542 21786
rect 6594 21734 13646 21786
rect 13698 21734 13710 21786
rect 13762 21734 13774 21786
rect 13826 21734 13838 21786
rect 13890 21734 13902 21786
rect 13954 21734 21006 21786
rect 21058 21734 21070 21786
rect 21122 21734 21134 21786
rect 21186 21734 21198 21786
rect 21250 21734 21262 21786
rect 21314 21734 28366 21786
rect 28418 21734 28430 21786
rect 28482 21734 28494 21786
rect 28546 21734 28558 21786
rect 28610 21734 28622 21786
rect 28674 21734 32200 21786
rect 2760 21712 32200 21734
rect 3145 21675 3203 21681
rect 3145 21641 3157 21675
rect 3191 21672 3203 21675
rect 3234 21672 3240 21684
rect 3191 21644 3240 21672
rect 3191 21641 3203 21644
rect 3145 21635 3203 21641
rect 3234 21632 3240 21644
rect 3292 21632 3298 21684
rect 6178 21632 6184 21684
rect 6236 21672 6242 21684
rect 6733 21675 6791 21681
rect 6733 21672 6745 21675
rect 6236 21644 6745 21672
rect 6236 21632 6242 21644
rect 6733 21641 6745 21644
rect 6779 21641 6791 21675
rect 6733 21635 6791 21641
rect 7466 21632 7472 21684
rect 7524 21632 7530 21684
rect 7926 21632 7932 21684
rect 7984 21632 7990 21684
rect 8110 21632 8116 21684
rect 8168 21672 8174 21684
rect 8297 21675 8355 21681
rect 8297 21672 8309 21675
rect 8168 21644 8309 21672
rect 8168 21632 8174 21644
rect 8297 21641 8309 21644
rect 8343 21672 8355 21675
rect 11330 21672 11336 21684
rect 8343 21644 11336 21672
rect 8343 21641 8355 21644
rect 8297 21635 8355 21641
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 11790 21632 11796 21684
rect 11848 21632 11854 21684
rect 11977 21675 12035 21681
rect 11977 21641 11989 21675
rect 12023 21672 12035 21675
rect 12802 21672 12808 21684
rect 12023 21644 12808 21672
rect 12023 21641 12035 21644
rect 11977 21635 12035 21641
rect 12802 21632 12808 21644
rect 12860 21632 12866 21684
rect 13467 21675 13525 21681
rect 13467 21641 13479 21675
rect 13513 21672 13525 21675
rect 13998 21672 14004 21684
rect 13513 21644 14004 21672
rect 13513 21641 13525 21644
rect 13467 21635 13525 21641
rect 13998 21632 14004 21644
rect 14056 21632 14062 21684
rect 14384 21644 14780 21672
rect 6822 21604 6828 21616
rect 5736 21576 6828 21604
rect 5077 21539 5135 21545
rect 5077 21536 5089 21539
rect 3528 21508 5089 21536
rect 3528 21454 3556 21508
rect 5077 21505 5089 21508
rect 5123 21505 5135 21539
rect 5077 21499 5135 21505
rect 5736 21477 5764 21576
rect 6822 21564 6828 21576
rect 6880 21604 6886 21616
rect 8478 21604 8484 21616
rect 6880 21576 8484 21604
rect 6880 21564 6886 21576
rect 5994 21496 6000 21548
rect 6052 21496 6058 21548
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21536 6699 21539
rect 6730 21536 6736 21548
rect 6687 21508 6736 21536
rect 6687 21505 6699 21508
rect 6641 21499 6699 21505
rect 6730 21496 6736 21508
rect 6788 21536 6794 21548
rect 6788 21508 7052 21536
rect 6788 21496 6794 21508
rect 7024 21477 7052 21508
rect 4893 21471 4951 21477
rect 4893 21437 4905 21471
rect 4939 21437 4951 21471
rect 4893 21431 4951 21437
rect 5169 21471 5227 21477
rect 5169 21437 5181 21471
rect 5215 21468 5227 21471
rect 5721 21471 5779 21477
rect 5721 21468 5733 21471
rect 5215 21440 5733 21468
rect 5215 21437 5227 21440
rect 5169 21431 5227 21437
rect 5721 21437 5733 21440
rect 5767 21437 5779 21471
rect 5721 21431 5779 21437
rect 6917 21471 6975 21477
rect 6917 21437 6929 21471
rect 6963 21437 6975 21471
rect 6917 21431 6975 21437
rect 7009 21471 7067 21477
rect 7009 21437 7021 21471
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 4614 21360 4620 21412
rect 4672 21360 4678 21412
rect 4908 21400 4936 21431
rect 4724 21372 4936 21400
rect 4724 21344 4752 21372
rect 4706 21292 4712 21344
rect 4764 21292 4770 21344
rect 5718 21292 5724 21344
rect 5776 21332 5782 21344
rect 5813 21335 5871 21341
rect 5813 21332 5825 21335
rect 5776 21304 5825 21332
rect 5776 21292 5782 21304
rect 5813 21301 5825 21304
rect 5859 21301 5871 21335
rect 6932 21332 6960 21431
rect 7098 21428 7104 21480
rect 7156 21428 7162 21480
rect 7282 21428 7288 21480
rect 7340 21468 7346 21480
rect 7576 21477 7604 21576
rect 8478 21564 8484 21576
rect 8536 21564 8542 21616
rect 8386 21496 8392 21548
rect 8444 21536 8450 21548
rect 8665 21539 8723 21545
rect 8665 21536 8677 21539
rect 8444 21508 8677 21536
rect 8444 21496 8450 21508
rect 8665 21505 8677 21508
rect 8711 21536 8723 21539
rect 9582 21536 9588 21548
rect 8711 21508 9588 21536
rect 8711 21505 8723 21508
rect 8665 21499 8723 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 13725 21539 13783 21545
rect 9732 21508 12204 21536
rect 9732 21496 9738 21508
rect 7561 21471 7619 21477
rect 7340 21440 7512 21468
rect 7340 21428 7346 21440
rect 7484 21400 7512 21440
rect 7561 21437 7573 21471
rect 7607 21437 7619 21471
rect 7561 21431 7619 21437
rect 7926 21428 7932 21480
rect 7984 21428 7990 21480
rect 9950 21428 9956 21480
rect 10008 21468 10014 21480
rect 11425 21471 11483 21477
rect 10008 21440 10074 21468
rect 10008 21428 10014 21440
rect 11425 21437 11437 21471
rect 11471 21468 11483 21471
rect 11701 21471 11759 21477
rect 11701 21468 11713 21471
rect 11471 21440 11713 21468
rect 11471 21437 11483 21440
rect 11425 21431 11483 21437
rect 11701 21437 11713 21440
rect 11747 21468 11759 21471
rect 11747 21440 12112 21468
rect 11747 21437 11759 21440
rect 11701 21431 11759 21437
rect 7944 21400 7972 21428
rect 7484 21372 7972 21400
rect 8941 21403 8999 21409
rect 8941 21369 8953 21403
rect 8987 21369 8999 21403
rect 8941 21363 8999 21369
rect 8018 21332 8024 21344
rect 6932 21304 8024 21332
rect 5813 21295 5871 21301
rect 8018 21292 8024 21304
rect 8076 21292 8082 21344
rect 8956 21332 8984 21363
rect 10226 21360 10232 21412
rect 10284 21400 10290 21412
rect 10873 21403 10931 21409
rect 10873 21400 10885 21403
rect 10284 21372 10885 21400
rect 10284 21360 10290 21372
rect 10873 21369 10885 21372
rect 10919 21369 10931 21403
rect 10873 21363 10931 21369
rect 12084 21344 12112 21440
rect 9674 21332 9680 21344
rect 8956 21304 9680 21332
rect 9674 21292 9680 21304
rect 9732 21292 9738 21344
rect 10410 21292 10416 21344
rect 10468 21292 10474 21344
rect 12066 21292 12072 21344
rect 12124 21292 12130 21344
rect 12176 21332 12204 21508
rect 13725 21505 13737 21539
rect 13771 21505 13783 21539
rect 13725 21499 13783 21505
rect 12894 21360 12900 21412
rect 12952 21360 12958 21412
rect 13446 21360 13452 21412
rect 13504 21400 13510 21412
rect 13740 21400 13768 21499
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14277 21539 14335 21545
rect 14277 21536 14289 21539
rect 14240 21508 14289 21536
rect 14240 21496 14246 21508
rect 14277 21505 14289 21508
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 13504 21372 13768 21400
rect 13504 21360 13510 21372
rect 13998 21360 14004 21412
rect 14056 21400 14062 21412
rect 14093 21403 14151 21409
rect 14093 21400 14105 21403
rect 14056 21372 14105 21400
rect 14056 21360 14062 21372
rect 14093 21369 14105 21372
rect 14139 21369 14151 21403
rect 14093 21363 14151 21369
rect 14384 21332 14412 21644
rect 14645 21607 14703 21613
rect 14645 21573 14657 21607
rect 14691 21573 14703 21607
rect 14645 21567 14703 21573
rect 14461 21471 14519 21477
rect 14461 21437 14473 21471
rect 14507 21437 14519 21471
rect 14461 21431 14519 21437
rect 14553 21471 14611 21477
rect 14553 21437 14565 21471
rect 14599 21468 14611 21471
rect 14660 21468 14688 21567
rect 14599 21440 14688 21468
rect 14752 21468 14780 21644
rect 14826 21632 14832 21684
rect 14884 21672 14890 21684
rect 15194 21672 15200 21684
rect 14884 21644 15200 21672
rect 14884 21632 14890 21644
rect 15194 21632 15200 21644
rect 15252 21632 15258 21684
rect 16114 21632 16120 21684
rect 16172 21672 16178 21684
rect 16301 21675 16359 21681
rect 16301 21672 16313 21675
rect 16172 21644 16313 21672
rect 16172 21632 16178 21644
rect 16301 21641 16313 21644
rect 16347 21641 16359 21675
rect 16301 21635 16359 21641
rect 18230 21632 18236 21684
rect 18288 21632 18294 21684
rect 18414 21632 18420 21684
rect 18472 21632 18478 21684
rect 20349 21675 20407 21681
rect 20349 21641 20361 21675
rect 20395 21672 20407 21675
rect 20714 21672 20720 21684
rect 20395 21644 20720 21672
rect 20395 21641 20407 21644
rect 20349 21635 20407 21641
rect 20714 21632 20720 21644
rect 20772 21632 20778 21684
rect 20898 21632 20904 21684
rect 20956 21632 20962 21684
rect 21008 21644 24440 21672
rect 15562 21564 15568 21616
rect 15620 21604 15626 21616
rect 16206 21604 16212 21616
rect 15620 21576 16212 21604
rect 15620 21564 15626 21576
rect 16206 21564 16212 21576
rect 16264 21604 16270 21616
rect 17126 21604 17132 21616
rect 16264 21576 17132 21604
rect 16264 21564 16270 21576
rect 17126 21564 17132 21576
rect 17184 21564 17190 21616
rect 18432 21604 18460 21632
rect 21008 21604 21036 21644
rect 18432 21576 21036 21604
rect 23750 21564 23756 21616
rect 23808 21604 23814 21616
rect 24118 21604 24124 21616
rect 23808 21576 24124 21604
rect 23808 21564 23814 21576
rect 24118 21564 24124 21576
rect 24176 21604 24182 21616
rect 24176 21576 24348 21604
rect 24176 21564 24182 21576
rect 15013 21539 15071 21545
rect 15013 21505 15025 21539
rect 15059 21536 15071 21539
rect 18782 21536 18788 21548
rect 15059 21508 15240 21536
rect 15059 21505 15071 21508
rect 15013 21499 15071 21505
rect 14829 21471 14887 21477
rect 14829 21468 14841 21471
rect 14752 21440 14841 21468
rect 14599 21437 14611 21440
rect 14553 21431 14611 21437
rect 14829 21437 14841 21440
rect 14875 21468 14887 21471
rect 15102 21468 15108 21480
rect 14875 21440 15108 21468
rect 14875 21437 14887 21440
rect 14829 21431 14887 21437
rect 14476 21400 14504 21431
rect 15102 21428 15108 21440
rect 15160 21428 15166 21480
rect 15212 21400 15240 21508
rect 15396 21508 18788 21536
rect 15286 21428 15292 21480
rect 15344 21428 15350 21480
rect 15396 21400 15424 21508
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 19797 21539 19855 21545
rect 19797 21505 19809 21539
rect 19843 21505 19855 21539
rect 20622 21536 20628 21548
rect 19797 21499 19855 21505
rect 19996 21508 20628 21536
rect 15470 21428 15476 21480
rect 15528 21428 15534 21480
rect 15749 21471 15807 21477
rect 15749 21437 15761 21471
rect 15795 21468 15807 21471
rect 15838 21468 15844 21480
rect 15795 21440 15844 21468
rect 15795 21437 15807 21440
rect 15749 21431 15807 21437
rect 15838 21428 15844 21440
rect 15896 21428 15902 21480
rect 16117 21471 16175 21477
rect 16117 21437 16129 21471
rect 16163 21468 16175 21471
rect 16942 21468 16948 21480
rect 16163 21440 16948 21468
rect 16163 21437 16175 21440
rect 16117 21431 16175 21437
rect 16942 21428 16948 21440
rect 17000 21428 17006 21480
rect 17494 21468 17500 21480
rect 17052 21440 17500 21468
rect 14476 21372 15148 21400
rect 15212 21372 15424 21400
rect 15488 21400 15516 21428
rect 15933 21403 15991 21409
rect 15933 21400 15945 21403
rect 15488 21372 15945 21400
rect 12176 21304 14412 21332
rect 14553 21335 14611 21341
rect 14553 21301 14565 21335
rect 14599 21332 14611 21335
rect 15010 21332 15016 21344
rect 14599 21304 15016 21332
rect 14599 21301 14611 21304
rect 14553 21295 14611 21301
rect 15010 21292 15016 21304
rect 15068 21292 15074 21344
rect 15120 21332 15148 21372
rect 15933 21369 15945 21372
rect 15979 21369 15991 21403
rect 15933 21363 15991 21369
rect 16022 21360 16028 21412
rect 16080 21360 16086 21412
rect 16390 21360 16396 21412
rect 16448 21400 16454 21412
rect 16485 21403 16543 21409
rect 16485 21400 16497 21403
rect 16448 21372 16497 21400
rect 16448 21360 16454 21372
rect 16485 21369 16497 21372
rect 16531 21369 16543 21403
rect 16485 21363 16543 21369
rect 16666 21360 16672 21412
rect 16724 21400 16730 21412
rect 17052 21400 17080 21440
rect 17494 21428 17500 21440
rect 17552 21468 17558 21480
rect 17865 21471 17923 21477
rect 17865 21468 17877 21471
rect 17552 21440 17877 21468
rect 17552 21428 17558 21440
rect 17865 21437 17877 21440
rect 17911 21437 17923 21471
rect 17865 21431 17923 21437
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 18141 21471 18199 21477
rect 18141 21468 18153 21471
rect 18104 21440 18153 21468
rect 18104 21428 18110 21440
rect 18141 21437 18153 21440
rect 18187 21437 18199 21471
rect 18141 21431 18199 21437
rect 16724 21372 17080 21400
rect 16724 21360 16730 21372
rect 17126 21360 17132 21412
rect 17184 21360 17190 21412
rect 15654 21332 15660 21344
rect 15120 21304 15660 21332
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 15838 21292 15844 21344
rect 15896 21332 15902 21344
rect 16408 21332 16436 21360
rect 15896 21304 16436 21332
rect 15896 21292 15902 21304
rect 16574 21292 16580 21344
rect 16632 21332 16638 21344
rect 17218 21332 17224 21344
rect 16632 21304 17224 21332
rect 16632 21292 16638 21304
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 18800 21332 18828 21496
rect 19812 21412 19840 21499
rect 19996 21477 20024 21508
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 22373 21539 22431 21545
rect 22373 21505 22385 21539
rect 22419 21536 22431 21539
rect 22741 21539 22799 21545
rect 22741 21536 22753 21539
rect 22419 21508 22753 21536
rect 22419 21505 22431 21508
rect 22373 21499 22431 21505
rect 22741 21505 22753 21508
rect 22787 21505 22799 21539
rect 22741 21499 22799 21505
rect 19981 21471 20039 21477
rect 19981 21437 19993 21471
rect 20027 21437 20039 21471
rect 19981 21431 20039 21437
rect 20070 21428 20076 21480
rect 20128 21468 20134 21480
rect 20530 21468 20536 21480
rect 20128 21440 20536 21468
rect 20128 21428 20134 21440
rect 20530 21428 20536 21440
rect 20588 21428 20594 21480
rect 22649 21471 22707 21477
rect 22649 21437 22661 21471
rect 22695 21437 22707 21471
rect 22649 21431 22707 21437
rect 19794 21360 19800 21412
rect 19852 21400 19858 21412
rect 20625 21403 20683 21409
rect 19852 21372 20024 21400
rect 19852 21360 19858 21372
rect 19889 21335 19947 21341
rect 19889 21332 19901 21335
rect 18800 21304 19901 21332
rect 19889 21301 19901 21304
rect 19935 21301 19947 21335
rect 19996 21332 20024 21372
rect 20625 21369 20637 21403
rect 20671 21400 20683 21403
rect 20671 21372 21206 21400
rect 20671 21369 20683 21372
rect 20625 21363 20683 21369
rect 21450 21332 21456 21344
rect 19996 21304 21456 21332
rect 19889 21295 19947 21301
rect 21450 21292 21456 21304
rect 21508 21292 21514 21344
rect 22094 21292 22100 21344
rect 22152 21332 22158 21344
rect 22664 21332 22692 21431
rect 23290 21428 23296 21480
rect 23348 21428 23354 21480
rect 24121 21471 24179 21477
rect 24121 21437 24133 21471
rect 24167 21468 24179 21471
rect 24213 21471 24271 21477
rect 24213 21468 24225 21471
rect 24167 21440 24225 21468
rect 24167 21437 24179 21440
rect 24121 21431 24179 21437
rect 24213 21437 24225 21440
rect 24259 21437 24271 21471
rect 24320 21468 24348 21576
rect 24412 21536 24440 21644
rect 24486 21632 24492 21684
rect 24544 21672 24550 21684
rect 25501 21675 25559 21681
rect 25501 21672 25513 21675
rect 24544 21644 25513 21672
rect 24544 21632 24550 21644
rect 25501 21641 25513 21644
rect 25547 21641 25559 21675
rect 25501 21635 25559 21641
rect 26050 21632 26056 21684
rect 26108 21672 26114 21684
rect 26237 21675 26295 21681
rect 26237 21672 26249 21675
rect 26108 21644 26249 21672
rect 26108 21632 26114 21644
rect 26237 21641 26249 21644
rect 26283 21641 26295 21675
rect 27982 21672 27988 21684
rect 26237 21635 26295 21641
rect 26344 21644 27988 21672
rect 24581 21607 24639 21613
rect 24581 21573 24593 21607
rect 24627 21604 24639 21607
rect 24670 21604 24676 21616
rect 24627 21576 24676 21604
rect 24627 21573 24639 21576
rect 24581 21567 24639 21573
rect 24670 21564 24676 21576
rect 24728 21564 24734 21616
rect 25222 21564 25228 21616
rect 25280 21604 25286 21616
rect 26344 21604 26372 21644
rect 27982 21632 27988 21644
rect 28040 21632 28046 21684
rect 25280 21576 26372 21604
rect 27724 21576 28764 21604
rect 25280 21564 25286 21576
rect 26142 21536 26148 21548
rect 24412 21508 26148 21536
rect 26142 21496 26148 21508
rect 26200 21496 26206 21548
rect 26418 21496 26424 21548
rect 26476 21496 26482 21548
rect 26697 21539 26755 21545
rect 26697 21505 26709 21539
rect 26743 21536 26755 21539
rect 26786 21536 26792 21548
rect 26743 21508 26792 21536
rect 26743 21505 26755 21508
rect 26697 21499 26755 21505
rect 26786 21496 26792 21508
rect 26844 21496 26850 21548
rect 27062 21496 27068 21548
rect 27120 21536 27126 21548
rect 27724 21536 27752 21576
rect 28629 21539 28687 21545
rect 28629 21536 28641 21539
rect 27120 21508 27752 21536
rect 27816 21508 28641 21536
rect 27120 21496 27126 21508
rect 24397 21471 24455 21477
rect 24397 21468 24409 21471
rect 24320 21440 24409 21468
rect 24213 21431 24271 21437
rect 24397 21437 24409 21440
rect 24443 21437 24455 21471
rect 24397 21431 24455 21437
rect 24673 21471 24731 21477
rect 24673 21437 24685 21471
rect 24719 21468 24731 21471
rect 24946 21468 24952 21480
rect 24719 21440 24952 21468
rect 24719 21437 24731 21440
rect 24673 21431 24731 21437
rect 24946 21428 24952 21440
rect 25004 21428 25010 21480
rect 25038 21428 25044 21480
rect 25096 21468 25102 21480
rect 25317 21471 25375 21477
rect 25317 21468 25329 21471
rect 25096 21440 25329 21468
rect 25096 21428 25102 21440
rect 25317 21437 25329 21440
rect 25363 21437 25375 21471
rect 25317 21431 25375 21437
rect 25424 21440 26004 21468
rect 27816 21454 27844 21508
rect 28629 21505 28641 21508
rect 28675 21505 28687 21539
rect 28629 21499 28687 21505
rect 28736 21477 28764 21576
rect 30190 21496 30196 21548
rect 30248 21496 30254 21548
rect 28445 21471 28503 21477
rect 22830 21360 22836 21412
rect 22888 21400 22894 21412
rect 23382 21400 23388 21412
rect 22888 21372 23388 21400
rect 22888 21360 22894 21372
rect 23382 21360 23388 21372
rect 23440 21400 23446 21412
rect 25424 21400 25452 21440
rect 23440 21372 25452 21400
rect 23440 21360 23446 21372
rect 25682 21360 25688 21412
rect 25740 21360 25746 21412
rect 25866 21360 25872 21412
rect 25924 21360 25930 21412
rect 25976 21400 26004 21440
rect 28445 21437 28457 21471
rect 28491 21437 28503 21471
rect 28445 21431 28503 21437
rect 28721 21471 28779 21477
rect 28721 21437 28733 21471
rect 28767 21468 28779 21471
rect 30208 21468 30236 21496
rect 28767 21440 30236 21468
rect 28767 21437 28779 21440
rect 28721 21431 28779 21437
rect 26970 21400 26976 21412
rect 25976 21372 26976 21400
rect 26970 21360 26976 21372
rect 27028 21360 27034 21412
rect 28353 21403 28411 21409
rect 28353 21400 28365 21403
rect 28000 21372 28365 21400
rect 22152 21304 22692 21332
rect 23477 21335 23535 21341
rect 22152 21292 22158 21304
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 24026 21332 24032 21344
rect 23523 21304 24032 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24210 21292 24216 21344
rect 24268 21332 24274 21344
rect 24765 21335 24823 21341
rect 24765 21332 24777 21335
rect 24268 21304 24777 21332
rect 24268 21292 24274 21304
rect 24765 21301 24777 21304
rect 24811 21301 24823 21335
rect 24765 21295 24823 21301
rect 24946 21292 24952 21344
rect 25004 21332 25010 21344
rect 25406 21332 25412 21344
rect 25004 21304 25412 21332
rect 25004 21292 25010 21304
rect 25406 21292 25412 21304
rect 25464 21292 25470 21344
rect 25884 21332 25912 21360
rect 26510 21332 26516 21344
rect 25884 21304 26516 21332
rect 26510 21292 26516 21304
rect 26568 21332 26574 21344
rect 26786 21332 26792 21344
rect 26568 21304 26792 21332
rect 26568 21292 26574 21304
rect 26786 21292 26792 21304
rect 26844 21292 26850 21344
rect 27706 21292 27712 21344
rect 27764 21332 27770 21344
rect 28000 21332 28028 21372
rect 28353 21369 28365 21372
rect 28399 21369 28411 21403
rect 28460 21400 28488 21431
rect 28460 21372 28764 21400
rect 28353 21363 28411 21369
rect 28736 21344 28764 21372
rect 27764 21304 28028 21332
rect 27764 21292 27770 21304
rect 28166 21292 28172 21344
rect 28224 21292 28230 21344
rect 28718 21292 28724 21344
rect 28776 21292 28782 21344
rect 2760 21242 32200 21264
rect 2760 21190 6946 21242
rect 6998 21190 7010 21242
rect 7062 21190 7074 21242
rect 7126 21190 7138 21242
rect 7190 21190 7202 21242
rect 7254 21190 14306 21242
rect 14358 21190 14370 21242
rect 14422 21190 14434 21242
rect 14486 21190 14498 21242
rect 14550 21190 14562 21242
rect 14614 21190 21666 21242
rect 21718 21190 21730 21242
rect 21782 21190 21794 21242
rect 21846 21190 21858 21242
rect 21910 21190 21922 21242
rect 21974 21190 29026 21242
rect 29078 21190 29090 21242
rect 29142 21190 29154 21242
rect 29206 21190 29218 21242
rect 29270 21190 29282 21242
rect 29334 21190 32200 21242
rect 2760 21168 32200 21190
rect 4154 21088 4160 21140
rect 4212 21128 4218 21140
rect 4525 21131 4583 21137
rect 4525 21128 4537 21131
rect 4212 21100 4537 21128
rect 4212 21088 4218 21100
rect 4525 21097 4537 21100
rect 4571 21097 4583 21131
rect 4525 21091 4583 21097
rect 4614 21088 4620 21140
rect 4672 21128 4678 21140
rect 4893 21131 4951 21137
rect 4893 21128 4905 21131
rect 4672 21100 4905 21128
rect 4672 21088 4678 21100
rect 4893 21097 4905 21100
rect 4939 21097 4951 21131
rect 4893 21091 4951 21097
rect 11054 21088 11060 21140
rect 11112 21128 11118 21140
rect 11517 21131 11575 21137
rect 11112 21100 11468 21128
rect 11112 21088 11118 21100
rect 10042 21020 10048 21072
rect 10100 21020 10106 21072
rect 10778 21020 10784 21072
rect 10836 21020 10842 21072
rect 11440 21060 11468 21100
rect 11517 21097 11529 21131
rect 11563 21128 11575 21131
rect 11606 21128 11612 21140
rect 11563 21100 11612 21128
rect 11563 21097 11575 21100
rect 11517 21091 11575 21097
rect 11606 21088 11612 21100
rect 11664 21088 11670 21140
rect 14090 21088 14096 21140
rect 14148 21128 14154 21140
rect 14277 21131 14335 21137
rect 14277 21128 14289 21131
rect 14148 21100 14289 21128
rect 14148 21088 14154 21100
rect 14277 21097 14289 21100
rect 14323 21097 14335 21131
rect 14277 21091 14335 21097
rect 15102 21088 15108 21140
rect 15160 21128 15166 21140
rect 15841 21131 15899 21137
rect 15841 21128 15853 21131
rect 15160 21100 15853 21128
rect 15160 21088 15166 21100
rect 15841 21097 15853 21100
rect 15887 21128 15899 21131
rect 15887 21100 20576 21128
rect 15887 21097 15899 21100
rect 15841 21091 15899 21097
rect 11974 21060 11980 21072
rect 11440 21032 11980 21060
rect 11974 21020 11980 21032
rect 12032 21060 12038 21072
rect 12161 21063 12219 21069
rect 12161 21060 12173 21063
rect 12032 21032 12173 21060
rect 12032 21020 12038 21032
rect 12161 21029 12173 21032
rect 12207 21029 12219 21063
rect 12161 21023 12219 21029
rect 12434 21020 12440 21072
rect 12492 21060 12498 21072
rect 12713 21063 12771 21069
rect 12713 21060 12725 21063
rect 12492 21032 12725 21060
rect 12492 21020 12498 21032
rect 12713 21029 12725 21032
rect 12759 21060 12771 21063
rect 13354 21060 13360 21072
rect 12759 21032 13360 21060
rect 12759 21029 12771 21032
rect 12713 21023 12771 21029
rect 13354 21020 13360 21032
rect 13412 21020 13418 21072
rect 13538 21020 13544 21072
rect 13596 21060 13602 21072
rect 13909 21063 13967 21069
rect 13909 21060 13921 21063
rect 13596 21032 13921 21060
rect 13596 21020 13602 21032
rect 13909 21029 13921 21032
rect 13955 21029 13967 21063
rect 13909 21023 13967 21029
rect 14200 21032 15608 21060
rect 14200 21004 14228 21032
rect 3326 20952 3332 21004
rect 3384 20952 3390 21004
rect 4433 20995 4491 21001
rect 4433 20961 4445 20995
rect 4479 20992 4491 20995
rect 5902 20992 5908 21004
rect 4479 20964 5908 20992
rect 4479 20961 4491 20964
rect 4433 20955 4491 20961
rect 5902 20952 5908 20964
rect 5960 20992 5966 21004
rect 6181 20995 6239 21001
rect 6181 20992 6193 20995
rect 5960 20964 6193 20992
rect 5960 20952 5966 20964
rect 6181 20961 6193 20964
rect 6227 20961 6239 20995
rect 6181 20955 6239 20961
rect 9582 20952 9588 21004
rect 9640 20992 9646 21004
rect 9769 20995 9827 21001
rect 9769 20992 9781 20995
rect 9640 20964 9781 20992
rect 9640 20952 9646 20964
rect 9769 20961 9781 20964
rect 9815 20961 9827 20995
rect 9769 20955 9827 20961
rect 12176 20964 13032 20992
rect 3050 20884 3056 20936
rect 3108 20884 3114 20936
rect 4246 20884 4252 20936
rect 4304 20884 4310 20936
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 6730 20884 6736 20936
rect 6788 20884 6794 20936
rect 8202 20884 8208 20936
rect 8260 20924 8266 20936
rect 12176 20924 12204 20964
rect 13004 20936 13032 20964
rect 13262 20952 13268 21004
rect 13320 20992 13326 21004
rect 13449 20995 13507 21001
rect 13449 20992 13461 20995
rect 13320 20964 13461 20992
rect 13320 20952 13326 20964
rect 13449 20961 13461 20964
rect 13495 20992 13507 20995
rect 13495 20964 13860 20992
rect 13495 20961 13507 20964
rect 13449 20955 13507 20961
rect 13832 20936 13860 20964
rect 13998 20952 14004 21004
rect 14056 21001 14062 21004
rect 14056 20995 14084 21001
rect 14072 20961 14084 20995
rect 14056 20955 14084 20961
rect 14056 20952 14062 20955
rect 14182 20952 14188 21004
rect 14240 20952 14246 21004
rect 14458 20952 14464 21004
rect 14516 20992 14522 21004
rect 14829 20995 14887 21001
rect 14829 20992 14841 20995
rect 14516 20964 14841 20992
rect 14516 20952 14522 20964
rect 14829 20961 14841 20964
rect 14875 20961 14887 20995
rect 14829 20955 14887 20961
rect 15010 20952 15016 21004
rect 15068 20992 15074 21004
rect 15473 20995 15531 21001
rect 15473 20992 15485 20995
rect 15068 20964 15485 20992
rect 15068 20952 15074 20964
rect 15473 20961 15485 20964
rect 15519 20961 15531 20995
rect 15473 20955 15531 20961
rect 8260 20896 12204 20924
rect 8260 20884 8266 20896
rect 12250 20884 12256 20936
rect 12308 20884 12314 20936
rect 12986 20884 12992 20936
rect 13044 20884 13050 20936
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 12618 20816 12624 20868
rect 12676 20856 12682 20868
rect 12713 20859 12771 20865
rect 12713 20856 12725 20859
rect 12676 20828 12725 20856
rect 12676 20816 12682 20828
rect 12713 20825 12725 20828
rect 12759 20825 12771 20859
rect 12713 20819 12771 20825
rect 5258 20748 5264 20800
rect 5316 20748 5322 20800
rect 11977 20791 12035 20797
rect 11977 20757 11989 20791
rect 12023 20788 12035 20791
rect 12802 20788 12808 20800
rect 12023 20760 12808 20788
rect 12023 20757 12035 20760
rect 11977 20751 12035 20757
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 13556 20788 13584 20887
rect 13814 20884 13820 20936
rect 13872 20884 13878 20936
rect 15197 20927 15255 20933
rect 15197 20924 15209 20927
rect 14200 20896 15209 20924
rect 14200 20865 14228 20896
rect 15197 20893 15209 20896
rect 15243 20893 15255 20927
rect 15197 20887 15255 20893
rect 15289 20927 15347 20933
rect 15289 20893 15301 20927
rect 15335 20893 15347 20927
rect 15289 20887 15347 20893
rect 15381 20927 15439 20933
rect 15381 20893 15393 20927
rect 15427 20924 15439 20927
rect 15580 20924 15608 21032
rect 15930 21020 15936 21072
rect 15988 21060 15994 21072
rect 16485 21063 16543 21069
rect 16485 21060 16497 21063
rect 15988 21032 16497 21060
rect 15988 21020 15994 21032
rect 16485 21029 16497 21032
rect 16531 21060 16543 21063
rect 16850 21060 16856 21072
rect 16531 21032 16856 21060
rect 16531 21029 16543 21032
rect 16485 21023 16543 21029
rect 16850 21020 16856 21032
rect 16908 21020 16914 21072
rect 19058 21020 19064 21072
rect 19116 21020 19122 21072
rect 20073 21063 20131 21069
rect 20073 21029 20085 21063
rect 20119 21060 20131 21063
rect 20441 21063 20499 21069
rect 20441 21060 20453 21063
rect 20119 21032 20453 21060
rect 20119 21029 20131 21032
rect 20073 21023 20131 21029
rect 20441 21029 20453 21032
rect 20487 21029 20499 21063
rect 20548 21060 20576 21100
rect 20622 21088 20628 21140
rect 20680 21128 20686 21140
rect 22005 21131 22063 21137
rect 22005 21128 22017 21131
rect 20680 21100 22017 21128
rect 20680 21088 20686 21100
rect 22005 21097 22017 21100
rect 22051 21097 22063 21131
rect 22005 21091 22063 21097
rect 22465 21131 22523 21137
rect 22465 21097 22477 21131
rect 22511 21128 22523 21131
rect 23290 21128 23296 21140
rect 22511 21100 23296 21128
rect 22511 21097 22523 21100
rect 22465 21091 22523 21097
rect 23290 21088 23296 21100
rect 23348 21088 23354 21140
rect 23753 21131 23811 21137
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 23799 21100 24164 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 20898 21060 20904 21072
rect 20548 21032 20904 21060
rect 20441 21023 20499 21029
rect 20898 21020 20904 21032
rect 20956 21020 20962 21072
rect 21542 21020 21548 21072
rect 21600 21020 21606 21072
rect 22097 21063 22155 21069
rect 22097 21029 22109 21063
rect 22143 21060 22155 21063
rect 24136 21060 24164 21100
rect 24670 21088 24676 21140
rect 24728 21128 24734 21140
rect 25317 21131 25375 21137
rect 25317 21128 25329 21131
rect 24728 21100 25329 21128
rect 24728 21088 24734 21100
rect 25317 21097 25329 21100
rect 25363 21128 25375 21131
rect 27798 21128 27804 21140
rect 25363 21100 27804 21128
rect 25363 21097 25375 21100
rect 25317 21091 25375 21097
rect 27798 21088 27804 21100
rect 27856 21088 27862 21140
rect 28166 21088 28172 21140
rect 28224 21088 28230 21140
rect 25133 21063 25191 21069
rect 22143 21032 24072 21060
rect 22143 21029 22155 21032
rect 22097 21023 22155 21029
rect 15654 20952 15660 21004
rect 15712 20952 15718 21004
rect 20806 20952 20812 21004
rect 20864 20992 20870 21004
rect 21560 20992 21588 21020
rect 24044 21004 24072 21032
rect 24136 21032 24532 21060
rect 20864 20964 21588 20992
rect 20864 20952 20870 20964
rect 23566 20952 23572 21004
rect 23624 20992 23630 21004
rect 23661 20995 23719 21001
rect 23661 20992 23673 20995
rect 23624 20964 23673 20992
rect 23624 20952 23630 20964
rect 23661 20961 23673 20964
rect 23707 20961 23719 20995
rect 23661 20955 23719 20961
rect 24026 20952 24032 21004
rect 24084 20952 24090 21004
rect 24136 21001 24164 21032
rect 24121 20995 24179 21001
rect 24121 20961 24133 20995
rect 24167 20961 24179 20995
rect 24121 20955 24179 20961
rect 24210 20952 24216 21004
rect 24268 20992 24274 21004
rect 24305 20995 24363 21001
rect 24305 20992 24317 20995
rect 24268 20964 24317 20992
rect 24268 20952 24274 20964
rect 24305 20961 24317 20964
rect 24351 20961 24363 20995
rect 24305 20955 24363 20961
rect 24394 20952 24400 21004
rect 24452 20952 24458 21004
rect 15427 20896 15608 20924
rect 15427 20893 15439 20896
rect 15381 20887 15439 20893
rect 14185 20859 14243 20865
rect 14185 20825 14197 20859
rect 14231 20825 14243 20859
rect 15304 20856 15332 20887
rect 15672 20856 15700 20952
rect 18322 20884 18328 20936
rect 18380 20884 18386 20936
rect 20349 20927 20407 20933
rect 20349 20893 20361 20927
rect 20395 20893 20407 20927
rect 20349 20887 20407 20893
rect 15304 20828 15700 20856
rect 14185 20819 14243 20825
rect 14550 20788 14556 20800
rect 13556 20760 14556 20788
rect 14550 20748 14556 20760
rect 14608 20748 14614 20800
rect 14918 20748 14924 20800
rect 14976 20788 14982 20800
rect 15013 20791 15071 20797
rect 15013 20788 15025 20791
rect 14976 20760 15025 20788
rect 14976 20748 14982 20760
rect 15013 20757 15025 20760
rect 15059 20757 15071 20791
rect 15013 20751 15071 20757
rect 16666 20748 16672 20800
rect 16724 20788 16730 20800
rect 16853 20791 16911 20797
rect 16853 20788 16865 20791
rect 16724 20760 16865 20788
rect 16724 20748 16730 20760
rect 16853 20757 16865 20760
rect 16899 20788 16911 20791
rect 17034 20788 17040 20800
rect 16899 20760 17040 20788
rect 16899 20757 16911 20760
rect 16853 20751 16911 20757
rect 17034 20748 17040 20760
rect 17092 20788 17098 20800
rect 18340 20788 18368 20884
rect 20364 20856 20392 20887
rect 20714 20884 20720 20936
rect 20772 20924 20778 20936
rect 20993 20927 21051 20933
rect 20993 20924 21005 20927
rect 20772 20896 21005 20924
rect 20772 20884 20778 20896
rect 20993 20893 21005 20896
rect 21039 20893 21051 20927
rect 20993 20887 21051 20893
rect 21913 20927 21971 20933
rect 21913 20893 21925 20927
rect 21959 20924 21971 20927
rect 21959 20896 24164 20924
rect 21959 20893 21971 20896
rect 21913 20887 21971 20893
rect 24136 20868 24164 20896
rect 22094 20856 22100 20868
rect 20364 20828 22100 20856
rect 22094 20816 22100 20828
rect 22152 20816 22158 20868
rect 23014 20816 23020 20868
rect 23072 20856 23078 20868
rect 23072 20828 24072 20856
rect 23072 20816 23078 20828
rect 18690 20788 18696 20800
rect 17092 20760 18696 20788
rect 17092 20748 17098 20760
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 23934 20748 23940 20800
rect 23992 20748 23998 20800
rect 24044 20788 24072 20828
rect 24118 20816 24124 20868
rect 24176 20816 24182 20868
rect 24213 20859 24271 20865
rect 24213 20825 24225 20859
rect 24259 20825 24271 20859
rect 24504 20856 24532 21032
rect 25133 21029 25145 21063
rect 25179 21060 25191 21063
rect 25498 21060 25504 21072
rect 25179 21032 25504 21060
rect 25179 21029 25191 21032
rect 25133 21023 25191 21029
rect 25498 21020 25504 21032
rect 25556 21020 25562 21072
rect 27706 21060 27712 21072
rect 27278 21032 27712 21060
rect 27706 21020 27712 21032
rect 27764 21020 27770 21072
rect 24578 20952 24584 21004
rect 24636 20952 24642 21004
rect 24762 20952 24768 21004
rect 24820 20952 24826 21004
rect 24854 20952 24860 21004
rect 24912 20992 24918 21004
rect 25041 20995 25099 21001
rect 25041 20992 25053 20995
rect 24912 20964 25053 20992
rect 24912 20952 24918 20964
rect 25041 20961 25053 20964
rect 25087 20961 25099 20995
rect 25041 20955 25099 20961
rect 25409 20995 25467 21001
rect 25409 20961 25421 20995
rect 25455 20961 25467 20995
rect 25409 20955 25467 20961
rect 25314 20884 25320 20936
rect 25372 20924 25378 20936
rect 25424 20924 25452 20955
rect 25682 20952 25688 21004
rect 25740 20952 25746 21004
rect 28184 21001 28212 21088
rect 28169 20995 28227 21001
rect 28169 20961 28181 20995
rect 28215 20961 28227 20995
rect 28169 20955 28227 20961
rect 31849 20995 31907 21001
rect 31849 20961 31861 20995
rect 31895 20961 31907 20995
rect 31849 20955 31907 20961
rect 25372 20896 25452 20924
rect 25372 20884 25378 20896
rect 25498 20884 25504 20936
rect 25556 20884 25562 20936
rect 25700 20856 25728 20952
rect 25777 20927 25835 20933
rect 25777 20893 25789 20927
rect 25823 20893 25835 20927
rect 25777 20887 25835 20893
rect 24504 20828 25728 20856
rect 24213 20819 24271 20825
rect 24228 20788 24256 20819
rect 24857 20791 24915 20797
rect 24857 20788 24869 20791
rect 24044 20760 24869 20788
rect 24857 20757 24869 20760
rect 24903 20788 24915 20791
rect 24946 20788 24952 20800
rect 24903 20760 24952 20788
rect 24903 20757 24915 20760
rect 24857 20751 24915 20757
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 25682 20748 25688 20800
rect 25740 20748 25746 20800
rect 25792 20788 25820 20887
rect 26050 20884 26056 20936
rect 26108 20884 26114 20936
rect 26142 20884 26148 20936
rect 26200 20924 26206 20936
rect 27525 20927 27583 20933
rect 26200 20896 27108 20924
rect 26200 20884 26206 20896
rect 27080 20856 27108 20896
rect 27525 20893 27537 20927
rect 27571 20924 27583 20927
rect 29181 20927 29239 20933
rect 29181 20924 29193 20927
rect 27571 20896 29193 20924
rect 27571 20893 27583 20896
rect 27525 20887 27583 20893
rect 29181 20893 29193 20896
rect 29227 20893 29239 20927
rect 29181 20887 29239 20893
rect 29457 20927 29515 20933
rect 29457 20893 29469 20927
rect 29503 20924 29515 20927
rect 29546 20924 29552 20936
rect 29503 20896 29552 20924
rect 29503 20893 29515 20896
rect 29457 20887 29515 20893
rect 29546 20884 29552 20896
rect 29604 20884 29610 20936
rect 29638 20884 29644 20936
rect 29696 20924 29702 20936
rect 30653 20927 30711 20933
rect 30653 20924 30665 20927
rect 29696 20896 30665 20924
rect 29696 20884 29702 20896
rect 30653 20893 30665 20896
rect 30699 20893 30711 20927
rect 31864 20924 31892 20955
rect 33042 20924 33048 20936
rect 31864 20896 33048 20924
rect 30653 20887 30711 20893
rect 33042 20884 33048 20896
rect 33100 20884 33106 20936
rect 31665 20859 31723 20865
rect 31665 20856 31677 20859
rect 27080 20828 31677 20856
rect 31665 20825 31677 20828
rect 31711 20825 31723 20859
rect 31665 20819 31723 20825
rect 26418 20788 26424 20800
rect 25792 20760 26424 20788
rect 26418 20748 26424 20760
rect 26476 20748 26482 20800
rect 27614 20748 27620 20800
rect 27672 20748 27678 20800
rect 27706 20748 27712 20800
rect 27764 20788 27770 20800
rect 28629 20791 28687 20797
rect 28629 20788 28641 20791
rect 27764 20760 28641 20788
rect 27764 20748 27770 20760
rect 28629 20757 28641 20760
rect 28675 20757 28687 20791
rect 28629 20751 28687 20757
rect 30006 20748 30012 20800
rect 30064 20748 30070 20800
rect 30098 20748 30104 20800
rect 30156 20748 30162 20800
rect 2760 20698 32200 20720
rect 2760 20646 6286 20698
rect 6338 20646 6350 20698
rect 6402 20646 6414 20698
rect 6466 20646 6478 20698
rect 6530 20646 6542 20698
rect 6594 20646 13646 20698
rect 13698 20646 13710 20698
rect 13762 20646 13774 20698
rect 13826 20646 13838 20698
rect 13890 20646 13902 20698
rect 13954 20646 21006 20698
rect 21058 20646 21070 20698
rect 21122 20646 21134 20698
rect 21186 20646 21198 20698
rect 21250 20646 21262 20698
rect 21314 20646 28366 20698
rect 28418 20646 28430 20698
rect 28482 20646 28494 20698
rect 28546 20646 28558 20698
rect 28610 20646 28622 20698
rect 28674 20646 32200 20698
rect 2760 20624 32200 20646
rect 4246 20544 4252 20596
rect 4304 20584 4310 20596
rect 4801 20587 4859 20593
rect 4801 20584 4813 20587
rect 4304 20556 4813 20584
rect 4304 20544 4310 20556
rect 4801 20553 4813 20556
rect 4847 20553 4859 20587
rect 4801 20547 4859 20553
rect 5445 20587 5503 20593
rect 5445 20553 5457 20587
rect 5491 20584 5503 20587
rect 5810 20584 5816 20596
rect 5491 20556 5816 20584
rect 5491 20553 5503 20556
rect 5445 20547 5503 20553
rect 5810 20544 5816 20556
rect 5868 20544 5874 20596
rect 5920 20556 8064 20584
rect 5920 20516 5948 20556
rect 8036 20528 8064 20556
rect 9674 20544 9680 20596
rect 9732 20584 9738 20596
rect 10413 20587 10471 20593
rect 9732 20556 9996 20584
rect 9732 20544 9738 20556
rect 5644 20488 5948 20516
rect 5644 20389 5672 20488
rect 8018 20476 8024 20528
rect 8076 20476 8082 20528
rect 9968 20516 9996 20556
rect 10413 20553 10425 20587
rect 10459 20584 10471 20587
rect 10502 20584 10508 20596
rect 10459 20556 10508 20584
rect 10459 20553 10471 20556
rect 10413 20547 10471 20553
rect 10502 20544 10508 20556
rect 10560 20544 10566 20596
rect 11146 20544 11152 20596
rect 11204 20584 11210 20596
rect 11606 20584 11612 20596
rect 11204 20556 11612 20584
rect 11204 20544 11210 20556
rect 10597 20519 10655 20525
rect 10597 20516 10609 20519
rect 9968 20488 10609 20516
rect 10597 20485 10609 20488
rect 10643 20485 10655 20519
rect 10597 20479 10655 20485
rect 5810 20408 5816 20460
rect 5868 20448 5874 20460
rect 6086 20448 6092 20460
rect 5868 20420 6092 20448
rect 5868 20408 5874 20420
rect 6086 20408 6092 20420
rect 6144 20408 6150 20460
rect 7837 20451 7895 20457
rect 7837 20417 7849 20451
rect 7883 20448 7895 20451
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7883 20420 7941 20448
rect 7883 20417 7895 20420
rect 7837 20411 7895 20417
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 8386 20408 8392 20460
rect 8444 20448 8450 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 8444 20420 8677 20448
rect 8444 20408 8450 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 9582 20408 9588 20460
rect 9640 20448 9646 20460
rect 10870 20448 10876 20460
rect 9640 20420 10876 20448
rect 9640 20408 9646 20420
rect 10870 20408 10876 20420
rect 10928 20448 10934 20460
rect 11149 20451 11207 20457
rect 11149 20448 11161 20451
rect 10928 20420 11161 20448
rect 10928 20408 10934 20420
rect 11149 20417 11161 20420
rect 11195 20417 11207 20451
rect 11149 20411 11207 20417
rect 5629 20383 5687 20389
rect 5629 20349 5641 20383
rect 5675 20349 5687 20383
rect 5629 20343 5687 20349
rect 5721 20383 5779 20389
rect 5721 20349 5733 20383
rect 5767 20380 5779 20383
rect 5902 20380 5908 20392
rect 5767 20352 5908 20380
rect 5767 20349 5779 20352
rect 5721 20343 5779 20349
rect 5902 20340 5908 20352
rect 5960 20340 5966 20392
rect 5997 20383 6055 20389
rect 5997 20349 6009 20383
rect 6043 20380 6055 20383
rect 6043 20352 6132 20380
rect 6043 20349 6055 20352
rect 5997 20343 6055 20349
rect 5813 20315 5871 20321
rect 5813 20281 5825 20315
rect 5859 20281 5871 20315
rect 5813 20275 5871 20281
rect 5261 20247 5319 20253
rect 5261 20213 5273 20247
rect 5307 20244 5319 20247
rect 5828 20244 5856 20275
rect 5994 20244 6000 20256
rect 5307 20216 6000 20244
rect 5307 20213 5319 20216
rect 5261 20207 5319 20213
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6104 20244 6132 20352
rect 10042 20340 10048 20392
rect 10100 20340 10106 20392
rect 10965 20383 11023 20389
rect 10965 20349 10977 20383
rect 11011 20380 11023 20383
rect 11256 20380 11284 20556
rect 11606 20544 11612 20556
rect 11664 20544 11670 20596
rect 14182 20544 14188 20596
rect 14240 20544 14246 20596
rect 14550 20544 14556 20596
rect 14608 20584 14614 20596
rect 15286 20584 15292 20596
rect 14608 20556 15292 20584
rect 14608 20544 14614 20556
rect 15286 20544 15292 20556
rect 15344 20544 15350 20596
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15436 20556 15945 20584
rect 15436 20544 15442 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 18690 20544 18696 20596
rect 18748 20584 18754 20596
rect 18877 20587 18935 20593
rect 18877 20584 18889 20587
rect 18748 20556 18889 20584
rect 18748 20544 18754 20556
rect 18877 20553 18889 20556
rect 18923 20553 18935 20587
rect 18877 20547 18935 20553
rect 19058 20544 19064 20596
rect 19116 20584 19122 20596
rect 19153 20587 19211 20593
rect 19153 20584 19165 20587
rect 19116 20556 19165 20584
rect 19116 20544 19122 20556
rect 19153 20553 19165 20556
rect 19199 20553 19211 20587
rect 19153 20547 19211 20553
rect 20073 20587 20131 20593
rect 20073 20553 20085 20587
rect 20119 20584 20131 20587
rect 20714 20584 20720 20596
rect 20119 20556 20720 20584
rect 20119 20553 20131 20556
rect 20073 20547 20131 20553
rect 20714 20544 20720 20556
rect 20772 20544 20778 20596
rect 23934 20544 23940 20596
rect 23992 20544 23998 20596
rect 24118 20544 24124 20596
rect 24176 20584 24182 20596
rect 24397 20587 24455 20593
rect 24397 20584 24409 20587
rect 24176 20556 24409 20584
rect 24176 20544 24182 20556
rect 24397 20553 24409 20556
rect 24443 20553 24455 20587
rect 24397 20547 24455 20553
rect 24765 20587 24823 20593
rect 24765 20553 24777 20587
rect 24811 20584 24823 20587
rect 25038 20584 25044 20596
rect 24811 20556 25044 20584
rect 24811 20553 24823 20556
rect 24765 20547 24823 20553
rect 16574 20516 16580 20528
rect 12176 20488 16580 20516
rect 11974 20408 11980 20460
rect 12032 20408 12038 20460
rect 11011 20352 11284 20380
rect 11011 20349 11023 20352
rect 10965 20343 11023 20349
rect 6362 20272 6368 20324
rect 6420 20272 6426 20324
rect 7374 20272 7380 20324
rect 7432 20272 7438 20324
rect 8938 20272 8944 20324
rect 8996 20272 9002 20324
rect 11054 20272 11060 20324
rect 11112 20272 11118 20324
rect 7282 20244 7288 20256
rect 6104 20216 7288 20244
rect 7282 20204 7288 20216
rect 7340 20204 7346 20256
rect 8110 20204 8116 20256
rect 8168 20244 8174 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8168 20216 8585 20244
rect 8168 20204 8174 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9306 20204 9312 20256
rect 9364 20244 9370 20256
rect 12176 20244 12204 20488
rect 16574 20476 16580 20488
rect 16632 20476 16638 20528
rect 16684 20488 21404 20516
rect 12250 20408 12256 20460
rect 12308 20408 12314 20460
rect 12434 20408 12440 20460
rect 12492 20457 12498 20460
rect 12492 20451 12520 20457
rect 12508 20417 12520 20451
rect 14642 20448 14648 20460
rect 12492 20411 12520 20417
rect 14016 20420 14648 20448
rect 12492 20408 12498 20411
rect 12268 20380 12296 20408
rect 12345 20383 12403 20389
rect 12345 20380 12357 20383
rect 12268 20352 12357 20380
rect 12345 20349 12357 20352
rect 12391 20349 12403 20383
rect 12345 20343 12403 20349
rect 12618 20340 12624 20392
rect 12676 20340 12682 20392
rect 14016 20389 14044 20420
rect 14642 20408 14648 20420
rect 14700 20408 14706 20460
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 15252 20420 15485 20448
rect 15252 20408 15258 20420
rect 15473 20417 15485 20420
rect 15519 20448 15531 20451
rect 16684 20448 16712 20488
rect 21376 20460 21404 20488
rect 15519 20420 16712 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 18690 20408 18696 20460
rect 18748 20448 18754 20460
rect 19521 20451 19579 20457
rect 18748 20420 19472 20448
rect 18748 20408 18754 20420
rect 14001 20383 14059 20389
rect 14001 20349 14013 20383
rect 14047 20349 14059 20383
rect 14001 20343 14059 20349
rect 14093 20383 14151 20389
rect 14093 20349 14105 20383
rect 14139 20380 14151 20383
rect 14139 20352 14688 20380
rect 14139 20349 14151 20352
rect 14093 20343 14151 20349
rect 12636 20312 12664 20340
rect 12268 20284 12434 20312
rect 12268 20253 12296 20284
rect 9364 20216 12204 20244
rect 12253 20247 12311 20253
rect 9364 20204 9370 20216
rect 12253 20213 12265 20247
rect 12299 20213 12311 20247
rect 12406 20244 12434 20284
rect 12544 20284 12664 20312
rect 12544 20244 12572 20284
rect 14660 20256 14688 20352
rect 14734 20340 14740 20392
rect 14792 20380 14798 20392
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 14792 20352 15025 20380
rect 14792 20340 14798 20352
rect 15013 20349 15025 20352
rect 15059 20380 15071 20383
rect 15378 20380 15384 20392
rect 15059 20352 15384 20380
rect 15059 20349 15071 20352
rect 15013 20343 15071 20349
rect 15378 20340 15384 20352
rect 15436 20380 15442 20392
rect 15930 20380 15936 20392
rect 15436 20352 15936 20380
rect 15436 20340 15442 20352
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 19058 20340 19064 20392
rect 19116 20380 19122 20392
rect 19444 20380 19472 20420
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19794 20448 19800 20460
rect 19567 20420 19800 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 21358 20408 21364 20460
rect 21416 20408 21422 20460
rect 22094 20408 22100 20460
rect 22152 20448 22158 20460
rect 22833 20451 22891 20457
rect 22833 20448 22845 20451
rect 22152 20420 22845 20448
rect 22152 20408 22158 20420
rect 22833 20417 22845 20420
rect 22879 20417 22891 20451
rect 22833 20411 22891 20417
rect 23569 20451 23627 20457
rect 23569 20417 23581 20451
rect 23615 20448 23627 20451
rect 23952 20448 23980 20544
rect 23615 20420 23980 20448
rect 23615 20417 23627 20420
rect 23569 20411 23627 20417
rect 24026 20408 24032 20460
rect 24084 20408 24090 20460
rect 24670 20408 24676 20460
rect 24728 20408 24734 20460
rect 19613 20383 19671 20389
rect 19613 20380 19625 20383
rect 19116 20352 19288 20380
rect 19444 20352 19625 20380
rect 19116 20340 19122 20352
rect 19260 20312 19288 20352
rect 19613 20349 19625 20352
rect 19659 20349 19671 20383
rect 19613 20343 19671 20349
rect 22922 20340 22928 20392
rect 22980 20380 22986 20392
rect 23293 20383 23351 20389
rect 23293 20380 23305 20383
rect 22980 20352 23305 20380
rect 22980 20340 22986 20352
rect 23293 20349 23305 20352
rect 23339 20349 23351 20383
rect 23293 20343 23351 20349
rect 19978 20312 19984 20324
rect 19260 20284 19984 20312
rect 19978 20272 19984 20284
rect 20036 20272 20042 20324
rect 22002 20272 22008 20324
rect 22060 20272 22066 20324
rect 22557 20315 22615 20321
rect 22557 20281 22569 20315
rect 22603 20312 22615 20315
rect 22603 20284 23152 20312
rect 22603 20281 22615 20284
rect 22557 20275 22615 20281
rect 12406 20216 12572 20244
rect 12621 20247 12679 20253
rect 12253 20207 12311 20213
rect 12621 20213 12633 20247
rect 12667 20244 12679 20247
rect 12710 20244 12716 20256
rect 12667 20216 12716 20244
rect 12667 20213 12679 20216
rect 12621 20207 12679 20213
rect 12710 20204 12716 20216
rect 12768 20204 12774 20256
rect 13078 20204 13084 20256
rect 13136 20244 13142 20256
rect 13538 20244 13544 20256
rect 13136 20216 13544 20244
rect 13136 20204 13142 20216
rect 13538 20204 13544 20216
rect 13596 20244 13602 20256
rect 13633 20247 13691 20253
rect 13633 20244 13645 20247
rect 13596 20216 13645 20244
rect 13596 20204 13602 20216
rect 13633 20213 13645 20216
rect 13679 20213 13691 20247
rect 13633 20207 13691 20213
rect 13909 20247 13967 20253
rect 13909 20213 13921 20247
rect 13955 20244 13967 20247
rect 14090 20244 14096 20256
rect 13955 20216 14096 20244
rect 13955 20213 13967 20216
rect 13909 20207 13967 20213
rect 14090 20204 14096 20216
rect 14148 20204 14154 20256
rect 14642 20204 14648 20256
rect 14700 20204 14706 20256
rect 14734 20204 14740 20256
rect 14792 20244 14798 20256
rect 15654 20244 15660 20256
rect 14792 20216 15660 20244
rect 14792 20204 14798 20216
rect 15654 20204 15660 20216
rect 15712 20204 15718 20256
rect 19705 20247 19763 20253
rect 19705 20213 19717 20247
rect 19751 20244 19763 20247
rect 20438 20244 20444 20256
rect 19751 20216 20444 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 21082 20204 21088 20256
rect 21140 20204 21146 20256
rect 23124 20253 23152 20284
rect 23109 20247 23167 20253
rect 23109 20213 23121 20247
rect 23155 20213 23167 20247
rect 23308 20244 23336 20343
rect 23382 20340 23388 20392
rect 23440 20340 23446 20392
rect 23477 20383 23535 20389
rect 23477 20349 23489 20383
rect 23523 20380 23535 20383
rect 23750 20380 23756 20392
rect 23523 20352 23756 20380
rect 23523 20349 23535 20352
rect 23477 20343 23535 20349
rect 23750 20340 23756 20352
rect 23808 20340 23814 20392
rect 23842 20340 23848 20392
rect 23900 20340 23906 20392
rect 23937 20383 23995 20389
rect 23937 20349 23949 20383
rect 23983 20349 23995 20383
rect 23937 20343 23995 20349
rect 23400 20312 23428 20340
rect 23952 20312 23980 20343
rect 24118 20340 24124 20392
rect 24176 20340 24182 20392
rect 23400 20284 23980 20312
rect 23934 20244 23940 20256
rect 23308 20216 23940 20244
rect 23109 20207 23167 20213
rect 23934 20204 23940 20216
rect 23992 20204 23998 20256
rect 24302 20204 24308 20256
rect 24360 20204 24366 20256
rect 24670 20204 24676 20256
rect 24728 20244 24734 20256
rect 24780 20244 24808 20547
rect 25038 20544 25044 20556
rect 25096 20544 25102 20596
rect 25133 20587 25191 20593
rect 25133 20553 25145 20587
rect 25179 20584 25191 20587
rect 25498 20584 25504 20596
rect 25179 20556 25504 20584
rect 25179 20553 25191 20556
rect 25133 20547 25191 20553
rect 25498 20544 25504 20556
rect 25556 20544 25562 20596
rect 25590 20544 25596 20596
rect 25648 20544 25654 20596
rect 25682 20544 25688 20596
rect 25740 20584 25746 20596
rect 26678 20587 26736 20593
rect 26678 20584 26690 20587
rect 25740 20556 26690 20584
rect 25740 20544 25746 20556
rect 26678 20553 26690 20556
rect 26724 20553 26736 20587
rect 26678 20547 26736 20553
rect 26786 20544 26792 20596
rect 26844 20584 26850 20596
rect 27982 20584 27988 20596
rect 26844 20556 27988 20584
rect 26844 20544 26850 20556
rect 27982 20544 27988 20556
rect 28040 20544 28046 20596
rect 28169 20587 28227 20593
rect 28169 20553 28181 20587
rect 28215 20584 28227 20587
rect 29638 20584 29644 20596
rect 28215 20556 29644 20584
rect 28215 20553 28227 20556
rect 28169 20547 28227 20553
rect 29638 20544 29644 20556
rect 29696 20544 29702 20596
rect 29822 20544 29828 20596
rect 29880 20584 29886 20596
rect 30561 20587 30619 20593
rect 30561 20584 30573 20587
rect 29880 20556 30573 20584
rect 29880 20544 29886 20556
rect 30561 20553 30573 20556
rect 30607 20553 30619 20587
rect 30561 20547 30619 20553
rect 25608 20516 25636 20544
rect 26142 20516 26148 20528
rect 25608 20488 26148 20516
rect 26142 20476 26148 20488
rect 26200 20476 26206 20528
rect 25130 20408 25136 20460
rect 25188 20448 25194 20460
rect 25498 20448 25504 20460
rect 25188 20420 25504 20448
rect 25188 20408 25194 20420
rect 25498 20408 25504 20420
rect 25556 20408 25562 20460
rect 26418 20408 26424 20460
rect 26476 20448 26482 20460
rect 29362 20448 29368 20460
rect 26476 20420 29368 20448
rect 26476 20408 26482 20420
rect 29362 20408 29368 20420
rect 29420 20448 29426 20460
rect 30285 20451 30343 20457
rect 30285 20448 30297 20451
rect 29420 20420 30297 20448
rect 29420 20408 29426 20420
rect 30285 20417 30297 20420
rect 30331 20417 30343 20451
rect 30285 20411 30343 20417
rect 24854 20340 24860 20392
rect 24912 20380 24918 20392
rect 24949 20383 25007 20389
rect 24949 20380 24961 20383
rect 24912 20352 24961 20380
rect 24912 20340 24918 20352
rect 24949 20349 24961 20352
rect 24995 20349 25007 20383
rect 24949 20343 25007 20349
rect 25409 20383 25467 20389
rect 25409 20349 25421 20383
rect 25455 20349 25467 20383
rect 25409 20343 25467 20349
rect 25424 20312 25452 20343
rect 25682 20340 25688 20392
rect 25740 20340 25746 20392
rect 25774 20340 25780 20392
rect 25832 20380 25838 20392
rect 25869 20383 25927 20389
rect 25869 20380 25881 20383
rect 25832 20352 25881 20380
rect 25832 20340 25838 20352
rect 25869 20349 25881 20352
rect 25915 20349 25927 20383
rect 25869 20343 25927 20349
rect 26053 20383 26111 20389
rect 26053 20349 26065 20383
rect 26099 20380 26111 20383
rect 26326 20380 26332 20392
rect 26099 20352 26332 20380
rect 26099 20349 26111 20352
rect 26053 20343 26111 20349
rect 26326 20340 26332 20352
rect 26384 20340 26390 20392
rect 28166 20340 28172 20392
rect 28224 20380 28230 20392
rect 28261 20383 28319 20389
rect 28261 20380 28273 20383
rect 28224 20352 28273 20380
rect 28224 20340 28230 20352
rect 28261 20349 28273 20352
rect 28307 20349 28319 20383
rect 28261 20343 28319 20349
rect 28074 20312 28080 20324
rect 25424 20284 27108 20312
rect 27922 20284 28080 20312
rect 26694 20244 26700 20256
rect 24728 20216 26700 20244
rect 24728 20204 24734 20216
rect 26694 20204 26700 20216
rect 26752 20204 26758 20256
rect 27080 20244 27108 20284
rect 28074 20272 28080 20284
rect 28132 20272 28138 20324
rect 29454 20272 29460 20324
rect 29512 20272 29518 20324
rect 30006 20272 30012 20324
rect 30064 20272 30070 20324
rect 28166 20244 28172 20256
rect 27080 20216 28172 20244
rect 28166 20204 28172 20216
rect 28224 20244 28230 20256
rect 30098 20244 30104 20256
rect 28224 20216 30104 20244
rect 28224 20204 28230 20216
rect 30098 20204 30104 20216
rect 30156 20204 30162 20256
rect 30650 20204 30656 20256
rect 30708 20244 30714 20256
rect 30929 20247 30987 20253
rect 30929 20244 30941 20247
rect 30708 20216 30941 20244
rect 30708 20204 30714 20216
rect 30929 20213 30941 20216
rect 30975 20213 30987 20247
rect 30929 20207 30987 20213
rect 31202 20204 31208 20256
rect 31260 20244 31266 20256
rect 31389 20247 31447 20253
rect 31389 20244 31401 20247
rect 31260 20216 31401 20244
rect 31260 20204 31266 20216
rect 31389 20213 31401 20216
rect 31435 20213 31447 20247
rect 31389 20207 31447 20213
rect 2760 20154 32200 20176
rect 2760 20102 6946 20154
rect 6998 20102 7010 20154
rect 7062 20102 7074 20154
rect 7126 20102 7138 20154
rect 7190 20102 7202 20154
rect 7254 20102 14306 20154
rect 14358 20102 14370 20154
rect 14422 20102 14434 20154
rect 14486 20102 14498 20154
rect 14550 20102 14562 20154
rect 14614 20102 21666 20154
rect 21718 20102 21730 20154
rect 21782 20102 21794 20154
rect 21846 20102 21858 20154
rect 21910 20102 21922 20154
rect 21974 20102 29026 20154
rect 29078 20102 29090 20154
rect 29142 20102 29154 20154
rect 29206 20102 29218 20154
rect 29270 20102 29282 20154
rect 29334 20102 32200 20154
rect 2760 20080 32200 20102
rect 6362 20000 6368 20052
rect 6420 20000 6426 20052
rect 6457 20043 6515 20049
rect 6457 20009 6469 20043
rect 6503 20040 6515 20043
rect 6730 20040 6736 20052
rect 6503 20012 6736 20040
rect 6503 20009 6515 20012
rect 6457 20003 6515 20009
rect 6730 20000 6736 20012
rect 6788 20000 6794 20052
rect 7101 20043 7159 20049
rect 7101 20009 7113 20043
rect 7147 20040 7159 20043
rect 7374 20040 7380 20052
rect 7147 20012 7380 20040
rect 7147 20009 7159 20012
rect 7101 20003 7159 20009
rect 7374 20000 7380 20012
rect 7432 20000 7438 20052
rect 8021 20043 8079 20049
rect 8021 20009 8033 20043
rect 8067 20009 8079 20043
rect 8021 20003 8079 20009
rect 4985 19975 5043 19981
rect 4985 19941 4997 19975
rect 5031 19972 5043 19975
rect 5258 19972 5264 19984
rect 5031 19944 5264 19972
rect 5031 19941 5043 19944
rect 4985 19935 5043 19941
rect 5258 19932 5264 19944
rect 5316 19932 5322 19984
rect 5718 19932 5724 19984
rect 5776 19932 5782 19984
rect 6380 19972 6408 20000
rect 8036 19972 8064 20003
rect 8938 20000 8944 20052
rect 8996 20040 9002 20052
rect 9401 20043 9459 20049
rect 9401 20040 9413 20043
rect 8996 20012 9413 20040
rect 8996 20000 9002 20012
rect 9401 20009 9413 20012
rect 9447 20009 9459 20043
rect 9401 20003 9459 20009
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 10137 20043 10195 20049
rect 10137 20040 10149 20043
rect 10100 20012 10149 20040
rect 10100 20000 10106 20012
rect 10137 20009 10149 20012
rect 10183 20009 10195 20043
rect 10137 20003 10195 20009
rect 11606 20000 11612 20052
rect 11664 20040 11670 20052
rect 14369 20043 14427 20049
rect 14369 20040 14381 20043
rect 11664 20012 14381 20040
rect 11664 20000 11670 20012
rect 14369 20009 14381 20012
rect 14415 20040 14427 20043
rect 14734 20040 14740 20052
rect 14415 20012 14740 20040
rect 14415 20009 14427 20012
rect 14369 20003 14427 20009
rect 14734 20000 14740 20012
rect 14792 20000 14798 20052
rect 14829 20043 14887 20049
rect 14829 20009 14841 20043
rect 14875 20040 14887 20043
rect 15102 20040 15108 20052
rect 14875 20012 15108 20040
rect 14875 20009 14887 20012
rect 14829 20003 14887 20009
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15197 20043 15255 20049
rect 15197 20009 15209 20043
rect 15243 20040 15255 20043
rect 16482 20040 16488 20052
rect 15243 20012 16488 20040
rect 15243 20009 15255 20012
rect 15197 20003 15255 20009
rect 16482 20000 16488 20012
rect 16540 20000 16546 20052
rect 19058 20000 19064 20052
rect 19116 20000 19122 20052
rect 19242 20000 19248 20052
rect 19300 20000 19306 20052
rect 20438 20000 20444 20052
rect 20496 20000 20502 20052
rect 21082 20000 21088 20052
rect 21140 20000 21146 20052
rect 22002 20000 22008 20052
rect 22060 20040 22066 20052
rect 22097 20043 22155 20049
rect 22097 20040 22109 20043
rect 22060 20012 22109 20040
rect 22060 20000 22066 20012
rect 22097 20009 22109 20012
rect 22143 20009 22155 20043
rect 23658 20040 23664 20052
rect 22097 20003 22155 20009
rect 22664 20012 23664 20040
rect 6380 19944 8064 19972
rect 8110 19932 8116 19984
rect 8168 19972 8174 19984
rect 8297 19975 8355 19981
rect 8297 19972 8309 19975
rect 8168 19944 8309 19972
rect 8168 19932 8174 19944
rect 8297 19941 8309 19944
rect 8343 19941 8355 19975
rect 8297 19935 8355 19941
rect 8389 19975 8447 19981
rect 8389 19941 8401 19975
rect 8435 19972 8447 19975
rect 9858 19972 9864 19984
rect 8435 19944 9864 19972
rect 8435 19941 8447 19944
rect 8389 19935 8447 19941
rect 9858 19932 9864 19944
rect 9916 19932 9922 19984
rect 14274 19932 14280 19984
rect 14332 19972 14338 19984
rect 14553 19975 14611 19981
rect 14553 19972 14565 19975
rect 14332 19944 14565 19972
rect 14332 19932 14338 19944
rect 14553 19941 14565 19944
rect 14599 19941 14611 19975
rect 14553 19935 14611 19941
rect 15013 19975 15071 19981
rect 15013 19941 15025 19975
rect 15059 19972 15071 19975
rect 15470 19972 15476 19984
rect 15059 19944 15476 19972
rect 15059 19941 15071 19944
rect 15013 19935 15071 19941
rect 15470 19932 15476 19944
rect 15528 19932 15534 19984
rect 15654 19932 15660 19984
rect 15712 19972 15718 19984
rect 16209 19975 16267 19981
rect 16209 19972 16221 19975
rect 15712 19944 16221 19972
rect 15712 19932 15718 19944
rect 16209 19941 16221 19944
rect 16255 19972 16267 19975
rect 16758 19972 16764 19984
rect 16255 19944 16764 19972
rect 16255 19941 16267 19944
rect 16209 19935 16267 19941
rect 16758 19932 16764 19944
rect 16816 19932 16822 19984
rect 6914 19864 6920 19916
rect 6972 19904 6978 19916
rect 7009 19907 7067 19913
rect 7009 19904 7021 19907
rect 6972 19876 7021 19904
rect 6972 19864 6978 19876
rect 7009 19873 7021 19876
rect 7055 19873 7067 19907
rect 7009 19867 7067 19873
rect 7282 19864 7288 19916
rect 7340 19864 7346 19916
rect 7374 19864 7380 19916
rect 7432 19904 7438 19916
rect 8128 19904 8156 19932
rect 7432 19876 8156 19904
rect 8205 19907 8263 19913
rect 7432 19864 7438 19876
rect 8205 19873 8217 19907
rect 8251 19873 8263 19907
rect 8205 19867 8263 19873
rect 8573 19907 8631 19913
rect 8573 19873 8585 19907
rect 8619 19904 8631 19907
rect 9306 19904 9312 19916
rect 8619 19876 9312 19904
rect 8619 19873 8631 19876
rect 8573 19867 8631 19873
rect 4706 19796 4712 19848
rect 4764 19836 4770 19848
rect 5718 19836 5724 19848
rect 4764 19808 5724 19836
rect 4764 19796 4770 19808
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 6825 19839 6883 19845
rect 6825 19805 6837 19839
rect 6871 19836 6883 19839
rect 7300 19836 7328 19864
rect 6871 19808 7328 19836
rect 6871 19805 6883 19808
rect 6825 19799 6883 19805
rect 8018 19796 8024 19848
rect 8076 19836 8082 19848
rect 8220 19836 8248 19867
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 9582 19864 9588 19916
rect 9640 19864 9646 19916
rect 9674 19864 9680 19916
rect 9732 19864 9738 19916
rect 9766 19864 9772 19916
rect 9824 19864 9830 19916
rect 9953 19907 10011 19913
rect 9953 19873 9965 19907
rect 9999 19873 10011 19907
rect 9953 19867 10011 19873
rect 9600 19836 9628 19864
rect 8076 19808 9628 19836
rect 9968 19836 9996 19867
rect 10226 19864 10232 19916
rect 10284 19864 10290 19916
rect 10410 19864 10416 19916
rect 10468 19904 10474 19916
rect 10781 19907 10839 19913
rect 10781 19904 10793 19907
rect 10468 19876 10793 19904
rect 10468 19864 10474 19876
rect 10781 19873 10793 19876
rect 10827 19873 10839 19907
rect 10781 19867 10839 19873
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11425 19907 11483 19913
rect 11425 19904 11437 19907
rect 11112 19876 11437 19904
rect 11112 19864 11118 19876
rect 11425 19873 11437 19876
rect 11471 19904 11483 19907
rect 12250 19904 12256 19916
rect 11471 19876 12256 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 12250 19864 12256 19876
rect 12308 19864 12314 19916
rect 12802 19864 12808 19916
rect 12860 19864 12866 19916
rect 12894 19864 12900 19916
rect 12952 19904 12958 19916
rect 13541 19907 13599 19913
rect 13541 19904 13553 19907
rect 12952 19876 13553 19904
rect 12952 19864 12958 19876
rect 13541 19873 13553 19876
rect 13587 19873 13599 19907
rect 14185 19907 14243 19913
rect 14185 19904 14197 19907
rect 13541 19867 13599 19873
rect 13740 19876 14197 19904
rect 9968 19808 10272 19836
rect 8076 19796 8082 19808
rect 5994 19728 6000 19780
rect 6052 19768 6058 19780
rect 9766 19768 9772 19780
rect 6052 19740 9772 19768
rect 6052 19728 6058 19740
rect 9766 19728 9772 19740
rect 9824 19728 9830 19780
rect 10244 19712 10272 19808
rect 11330 19728 11336 19780
rect 11388 19768 11394 19780
rect 11606 19768 11612 19780
rect 11388 19740 11612 19768
rect 11388 19728 11394 19740
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 12618 19728 12624 19780
rect 12676 19768 12682 19780
rect 12820 19768 12848 19864
rect 13262 19796 13268 19848
rect 13320 19796 13326 19848
rect 13354 19796 13360 19848
rect 13412 19796 13418 19848
rect 13740 19845 13768 19876
rect 14185 19873 14197 19876
rect 14231 19873 14243 19907
rect 14185 19867 14243 19873
rect 14734 19864 14740 19916
rect 14792 19864 14798 19916
rect 15105 19907 15163 19913
rect 15105 19873 15117 19907
rect 15151 19873 15163 19907
rect 15105 19867 15163 19873
rect 13449 19839 13507 19845
rect 13449 19805 13461 19839
rect 13495 19805 13507 19839
rect 13449 19799 13507 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 14645 19839 14703 19845
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14918 19836 14924 19848
rect 14691 19808 14924 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 13464 19768 13492 19799
rect 14292 19768 14320 19799
rect 14918 19796 14924 19808
rect 14976 19796 14982 19848
rect 15120 19836 15148 19867
rect 15562 19864 15568 19916
rect 15620 19864 15626 19916
rect 17957 19907 18015 19913
rect 17957 19873 17969 19907
rect 18003 19904 18015 19907
rect 18414 19904 18420 19916
rect 18003 19876 18420 19904
rect 18003 19873 18015 19876
rect 17957 19867 18015 19873
rect 18414 19864 18420 19876
rect 18472 19864 18478 19916
rect 18509 19907 18567 19913
rect 18509 19873 18521 19907
rect 18555 19904 18567 19907
rect 19076 19904 19104 20000
rect 21100 19913 21128 20000
rect 22204 19944 22600 19972
rect 22204 19913 22232 19944
rect 18555 19876 19104 19904
rect 21085 19907 21143 19913
rect 18555 19873 18567 19876
rect 18509 19867 18567 19873
rect 21085 19873 21097 19907
rect 21131 19873 21143 19907
rect 21085 19867 21143 19873
rect 22189 19907 22247 19913
rect 22189 19873 22201 19907
rect 22235 19873 22247 19907
rect 22189 19867 22247 19873
rect 22465 19907 22523 19913
rect 22465 19873 22477 19907
rect 22511 19873 22523 19907
rect 22465 19867 22523 19873
rect 15194 19836 15200 19848
rect 15120 19808 15200 19836
rect 15194 19796 15200 19808
rect 15252 19836 15258 19848
rect 15933 19839 15991 19845
rect 15933 19836 15945 19839
rect 15252 19808 15945 19836
rect 15252 19796 15258 19808
rect 15933 19805 15945 19808
rect 15979 19836 15991 19839
rect 18138 19836 18144 19848
rect 15979 19808 18144 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 18138 19796 18144 19808
rect 18196 19836 18202 19848
rect 18196 19808 20300 19836
rect 18196 19796 18202 19808
rect 12676 19740 13492 19768
rect 13556 19740 14688 19768
rect 12676 19728 12682 19740
rect 9214 19660 9220 19712
rect 9272 19660 9278 19712
rect 10226 19660 10232 19712
rect 10284 19700 10290 19712
rect 10597 19703 10655 19709
rect 10597 19700 10609 19703
rect 10284 19672 10609 19700
rect 10284 19660 10290 19672
rect 10597 19669 10609 19672
rect 10643 19700 10655 19703
rect 13556 19700 13584 19740
rect 10643 19672 13584 19700
rect 10643 19669 10655 19672
rect 10597 19663 10655 19669
rect 13998 19660 14004 19712
rect 14056 19660 14062 19712
rect 14660 19700 14688 19740
rect 14734 19728 14740 19780
rect 14792 19768 14798 19780
rect 15013 19771 15071 19777
rect 15013 19768 15025 19771
rect 14792 19740 15025 19768
rect 14792 19728 14798 19740
rect 15013 19737 15025 19740
rect 15059 19737 15071 19771
rect 15013 19731 15071 19737
rect 15381 19771 15439 19777
rect 15381 19737 15393 19771
rect 15427 19768 15439 19771
rect 16666 19768 16672 19780
rect 15427 19740 16672 19768
rect 15427 19737 15439 19740
rect 15381 19731 15439 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 16758 19728 16764 19780
rect 16816 19768 16822 19780
rect 20162 19768 20168 19780
rect 16816 19740 20168 19768
rect 16816 19728 16822 19740
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 20272 19712 20300 19808
rect 21726 19796 21732 19848
rect 21784 19796 21790 19848
rect 15286 19700 15292 19712
rect 14660 19672 15292 19700
rect 15286 19660 15292 19672
rect 15344 19660 15350 19712
rect 15470 19660 15476 19712
rect 15528 19700 15534 19712
rect 16206 19700 16212 19712
rect 15528 19672 16212 19700
rect 15528 19660 15534 19672
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 17678 19660 17684 19712
rect 17736 19700 17742 19712
rect 17865 19703 17923 19709
rect 17865 19700 17877 19703
rect 17736 19672 17877 19700
rect 17736 19660 17742 19672
rect 17865 19669 17877 19672
rect 17911 19669 17923 19703
rect 17865 19663 17923 19669
rect 18414 19660 18420 19712
rect 18472 19660 18478 19712
rect 20254 19660 20260 19712
rect 20312 19660 20318 19712
rect 21177 19703 21235 19709
rect 21177 19669 21189 19703
rect 21223 19700 21235 19703
rect 21542 19700 21548 19712
rect 21223 19672 21548 19700
rect 21223 19669 21235 19672
rect 21177 19663 21235 19669
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 22480 19700 22508 19867
rect 22572 19836 22600 19944
rect 22664 19913 22692 20012
rect 23658 20000 23664 20012
rect 23716 20000 23722 20052
rect 23842 20000 23848 20052
rect 23900 20000 23906 20052
rect 24578 20000 24584 20052
rect 24636 20040 24642 20052
rect 26326 20040 26332 20052
rect 24636 20012 26332 20040
rect 24636 20000 24642 20012
rect 26326 20000 26332 20012
rect 26384 20040 26390 20052
rect 27430 20040 27436 20052
rect 26384 20012 27436 20040
rect 26384 20000 26390 20012
rect 27430 20000 27436 20012
rect 27488 20000 27494 20052
rect 27522 20000 27528 20052
rect 27580 20040 27586 20052
rect 27580 20012 27844 20040
rect 27580 20000 27586 20012
rect 22741 19975 22799 19981
rect 22741 19941 22753 19975
rect 22787 19972 22799 19975
rect 23860 19972 23888 20000
rect 22787 19944 23888 19972
rect 22787 19941 22799 19944
rect 22741 19935 22799 19941
rect 23934 19932 23940 19984
rect 23992 19972 23998 19984
rect 23992 19944 26372 19972
rect 23992 19932 23998 19944
rect 26344 19916 26372 19944
rect 26528 19944 27660 19972
rect 22649 19907 22707 19913
rect 22649 19873 22661 19907
rect 22695 19873 22707 19907
rect 22649 19867 22707 19873
rect 22830 19864 22836 19916
rect 22888 19864 22894 19916
rect 22925 19907 22983 19913
rect 22925 19873 22937 19907
rect 22971 19873 22983 19907
rect 22925 19867 22983 19873
rect 22848 19836 22876 19864
rect 22572 19808 22876 19836
rect 22940 19836 22968 19867
rect 23014 19864 23020 19916
rect 23072 19864 23078 19916
rect 23198 19864 23204 19916
rect 23256 19864 23262 19916
rect 23566 19864 23572 19916
rect 23624 19904 23630 19916
rect 24029 19907 24087 19913
rect 24029 19904 24041 19907
rect 23624 19876 24041 19904
rect 23624 19864 23630 19876
rect 24029 19873 24041 19876
rect 24075 19904 24087 19907
rect 24489 19907 24547 19913
rect 24489 19904 24501 19907
rect 24075 19876 24501 19904
rect 24075 19873 24087 19876
rect 24029 19867 24087 19873
rect 24489 19873 24501 19876
rect 24535 19873 24547 19907
rect 24489 19867 24547 19873
rect 25682 19864 25688 19916
rect 25740 19904 25746 19916
rect 26053 19907 26111 19913
rect 26053 19904 26065 19907
rect 25740 19876 26065 19904
rect 25740 19864 25746 19876
rect 26053 19873 26065 19876
rect 26099 19904 26111 19907
rect 26099 19876 26188 19904
rect 26099 19873 26111 19876
rect 26053 19867 26111 19873
rect 23584 19836 23612 19864
rect 22940 19808 23612 19836
rect 23842 19796 23848 19848
rect 23900 19836 23906 19848
rect 24121 19839 24179 19845
rect 24121 19836 24133 19839
rect 23900 19808 24133 19836
rect 23900 19796 23906 19808
rect 24121 19805 24133 19808
rect 24167 19836 24179 19839
rect 24581 19839 24639 19845
rect 24581 19836 24593 19839
rect 24167 19808 24593 19836
rect 24167 19805 24179 19808
rect 24121 19799 24179 19805
rect 24581 19805 24593 19808
rect 24627 19836 24639 19839
rect 24762 19836 24768 19848
rect 24627 19808 24768 19836
rect 24627 19805 24639 19808
rect 24581 19799 24639 19805
rect 24762 19796 24768 19808
rect 24820 19836 24826 19848
rect 25700 19836 25728 19864
rect 24820 19808 25728 19836
rect 25777 19839 25835 19845
rect 24820 19796 24826 19808
rect 25777 19805 25789 19839
rect 25823 19805 25835 19839
rect 25777 19799 25835 19805
rect 22649 19771 22707 19777
rect 22649 19737 22661 19771
rect 22695 19768 22707 19771
rect 22922 19768 22928 19780
rect 22695 19740 22928 19768
rect 22695 19737 22707 19740
rect 22649 19731 22707 19737
rect 22922 19728 22928 19740
rect 22980 19728 22986 19780
rect 23109 19771 23167 19777
rect 23109 19737 23121 19771
rect 23155 19768 23167 19771
rect 24210 19768 24216 19780
rect 23155 19740 24216 19768
rect 23155 19737 23167 19740
rect 23109 19731 23167 19737
rect 24210 19728 24216 19740
rect 24268 19728 24274 19780
rect 25682 19768 25688 19780
rect 24688 19740 25688 19768
rect 22738 19700 22744 19712
rect 22480 19672 22744 19700
rect 22738 19660 22744 19672
rect 22796 19660 22802 19712
rect 23198 19660 23204 19712
rect 23256 19700 23262 19712
rect 24688 19700 24716 19740
rect 25682 19728 25688 19740
rect 25740 19728 25746 19780
rect 25792 19768 25820 19799
rect 26160 19768 26188 19876
rect 26326 19864 26332 19916
rect 26384 19864 26390 19916
rect 26528 19913 26556 19944
rect 27632 19916 27660 19944
rect 27706 19932 27712 19984
rect 27764 19932 27770 19984
rect 26513 19907 26571 19913
rect 26513 19873 26525 19907
rect 26559 19873 26571 19907
rect 26513 19867 26571 19873
rect 27525 19907 27583 19913
rect 27525 19873 27537 19907
rect 27571 19873 27583 19907
rect 27525 19867 27583 19873
rect 26694 19796 26700 19848
rect 26752 19836 26758 19848
rect 27540 19836 27568 19867
rect 27614 19864 27620 19916
rect 27672 19864 27678 19916
rect 27724 19836 27752 19932
rect 27816 19913 27844 20012
rect 28166 20000 28172 20052
rect 28224 20040 28230 20052
rect 28997 20043 29055 20049
rect 28997 20040 29009 20043
rect 28224 20012 29009 20040
rect 28224 20000 28230 20012
rect 28997 20009 29009 20012
rect 29043 20009 29055 20043
rect 28997 20003 29055 20009
rect 29365 20043 29423 20049
rect 29365 20009 29377 20043
rect 29411 20040 29423 20043
rect 29546 20040 29552 20052
rect 29411 20012 29552 20040
rect 29411 20009 29423 20012
rect 29365 20003 29423 20009
rect 29546 20000 29552 20012
rect 29604 20000 29610 20052
rect 29822 20000 29828 20052
rect 29880 20040 29886 20052
rect 29880 20012 31754 20040
rect 29880 20000 29886 20012
rect 28258 19932 28264 19984
rect 28316 19972 28322 19984
rect 28902 19972 28908 19984
rect 28316 19944 28908 19972
rect 28316 19932 28322 19944
rect 28902 19932 28908 19944
rect 28960 19932 28966 19984
rect 29914 19972 29920 19984
rect 29564 19944 29920 19972
rect 27801 19907 27859 19913
rect 27801 19873 27813 19907
rect 27847 19873 27859 19907
rect 27801 19867 27859 19873
rect 27893 19907 27951 19913
rect 27893 19873 27905 19907
rect 27939 19904 27951 19907
rect 27982 19904 27988 19916
rect 27939 19876 27988 19904
rect 27939 19873 27951 19876
rect 27893 19867 27951 19873
rect 27982 19864 27988 19876
rect 28040 19864 28046 19916
rect 28077 19907 28135 19913
rect 28077 19873 28089 19907
rect 28123 19873 28135 19907
rect 28077 19867 28135 19873
rect 26752 19808 27384 19836
rect 27540 19808 27752 19836
rect 26752 19796 26758 19808
rect 27356 19768 27384 19808
rect 27985 19771 28043 19777
rect 27985 19768 27997 19771
rect 25792 19740 26096 19768
rect 26160 19740 27292 19768
rect 27356 19740 27997 19768
rect 23256 19672 24716 19700
rect 23256 19660 23262 19672
rect 24762 19660 24768 19712
rect 24820 19700 24826 19712
rect 24857 19703 24915 19709
rect 24857 19700 24869 19703
rect 24820 19672 24869 19700
rect 24820 19660 24826 19672
rect 24857 19669 24869 19672
rect 24903 19669 24915 19703
rect 24857 19663 24915 19669
rect 25130 19660 25136 19712
rect 25188 19660 25194 19712
rect 25958 19660 25964 19712
rect 26016 19660 26022 19712
rect 26068 19700 26096 19740
rect 27264 19712 27292 19740
rect 27985 19737 27997 19740
rect 28031 19737 28043 19771
rect 27985 19731 28043 19737
rect 26602 19700 26608 19712
rect 26068 19672 26608 19700
rect 26602 19660 26608 19672
rect 26660 19660 26666 19712
rect 27246 19660 27252 19712
rect 27304 19660 27310 19712
rect 27798 19660 27804 19712
rect 27856 19700 27862 19712
rect 28092 19700 28120 19867
rect 28813 19839 28871 19845
rect 28813 19805 28825 19839
rect 28859 19836 28871 19839
rect 28994 19836 29000 19848
rect 28859 19808 29000 19836
rect 28859 19805 28871 19808
rect 28813 19799 28871 19805
rect 28994 19796 29000 19808
rect 29052 19836 29058 19848
rect 29564 19836 29592 19944
rect 29914 19932 29920 19944
rect 29972 19932 29978 19984
rect 29641 19907 29699 19913
rect 29641 19873 29653 19907
rect 29687 19873 29699 19907
rect 29641 19867 29699 19873
rect 29052 19808 29592 19836
rect 29052 19796 29058 19808
rect 28718 19728 28724 19780
rect 28776 19768 28782 19780
rect 29656 19768 29684 19867
rect 30650 19864 30656 19916
rect 30708 19864 30714 19916
rect 30834 19913 30840 19916
rect 30812 19907 30840 19913
rect 30812 19873 30824 19907
rect 30812 19867 30840 19873
rect 30834 19864 30840 19867
rect 30892 19864 30898 19916
rect 30929 19907 30987 19913
rect 30929 19873 30941 19907
rect 30975 19873 30987 19907
rect 31726 19904 31754 20012
rect 31849 19907 31907 19913
rect 31849 19904 31861 19907
rect 31726 19876 31861 19904
rect 30929 19867 30987 19873
rect 31849 19873 31861 19876
rect 31895 19873 31907 19907
rect 31849 19867 31907 19873
rect 30944 19836 30972 19867
rect 31478 19836 31484 19848
rect 30944 19808 31484 19836
rect 31478 19796 31484 19808
rect 31536 19796 31542 19848
rect 31665 19839 31723 19845
rect 31665 19805 31677 19839
rect 31711 19805 31723 19839
rect 31665 19799 31723 19805
rect 28776 19740 29684 19768
rect 28776 19728 28782 19740
rect 31202 19728 31208 19780
rect 31260 19728 31266 19780
rect 31386 19728 31392 19780
rect 31444 19768 31450 19780
rect 31680 19768 31708 19799
rect 31444 19740 31708 19768
rect 31444 19728 31450 19740
rect 27856 19672 28120 19700
rect 27856 19660 27862 19672
rect 28258 19660 28264 19712
rect 28316 19660 28322 19712
rect 29454 19660 29460 19712
rect 29512 19700 29518 19712
rect 29549 19703 29607 19709
rect 29549 19700 29561 19703
rect 29512 19672 29561 19700
rect 29512 19660 29518 19672
rect 29549 19669 29561 19672
rect 29595 19669 29607 19703
rect 29549 19663 29607 19669
rect 30006 19660 30012 19712
rect 30064 19660 30070 19712
rect 30650 19660 30656 19712
rect 30708 19700 30714 19712
rect 31220 19700 31248 19728
rect 30708 19672 31248 19700
rect 30708 19660 30714 19672
rect 2760 19610 32200 19632
rect 2760 19558 6286 19610
rect 6338 19558 6350 19610
rect 6402 19558 6414 19610
rect 6466 19558 6478 19610
rect 6530 19558 6542 19610
rect 6594 19558 13646 19610
rect 13698 19558 13710 19610
rect 13762 19558 13774 19610
rect 13826 19558 13838 19610
rect 13890 19558 13902 19610
rect 13954 19558 21006 19610
rect 21058 19558 21070 19610
rect 21122 19558 21134 19610
rect 21186 19558 21198 19610
rect 21250 19558 21262 19610
rect 21314 19558 28366 19610
rect 28418 19558 28430 19610
rect 28482 19558 28494 19610
rect 28546 19558 28558 19610
rect 28610 19558 28622 19610
rect 28674 19558 32200 19610
rect 2760 19536 32200 19558
rect 14182 19496 14188 19508
rect 12477 19468 14188 19496
rect 12477 19428 12505 19468
rect 14182 19456 14188 19468
rect 14240 19496 14246 19508
rect 14240 19468 18644 19496
rect 14240 19456 14246 19468
rect 12452 19400 12505 19428
rect 14277 19431 14335 19437
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19329 8539 19363
rect 8481 19323 8539 19329
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19360 9459 19363
rect 9582 19360 9588 19372
rect 9447 19332 9588 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 1302 19252 1308 19304
rect 1360 19292 1366 19304
rect 3053 19295 3111 19301
rect 3053 19292 3065 19295
rect 1360 19264 3065 19292
rect 1360 19252 1366 19264
rect 3053 19261 3065 19264
rect 3099 19261 3111 19295
rect 3053 19255 3111 19261
rect 7834 19252 7840 19304
rect 7892 19252 7898 19304
rect 8496 19292 8524 19323
rect 9582 19320 9588 19332
rect 9640 19360 9646 19372
rect 10042 19360 10048 19372
rect 9640 19332 10048 19360
rect 9640 19320 9646 19332
rect 10042 19320 10048 19332
rect 10100 19320 10106 19372
rect 9125 19295 9183 19301
rect 8496 19264 8892 19292
rect 8864 19168 8892 19264
rect 9125 19261 9137 19295
rect 9171 19292 9183 19295
rect 9214 19292 9220 19304
rect 9171 19264 9220 19292
rect 9171 19261 9183 19264
rect 9125 19255 9183 19261
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 10502 19292 10508 19304
rect 9324 19264 10508 19292
rect 3234 19116 3240 19168
rect 3292 19116 3298 19168
rect 8754 19116 8760 19168
rect 8812 19116 8818 19168
rect 8846 19116 8852 19168
rect 8904 19116 8910 19168
rect 8938 19116 8944 19168
rect 8996 19156 9002 19168
rect 9217 19159 9275 19165
rect 9217 19156 9229 19159
rect 8996 19128 9229 19156
rect 8996 19116 9002 19128
rect 9217 19125 9229 19128
rect 9263 19156 9275 19159
rect 9324 19156 9352 19264
rect 10502 19252 10508 19264
rect 10560 19252 10566 19304
rect 10686 19252 10692 19304
rect 10744 19252 10750 19304
rect 11790 19252 11796 19304
rect 11848 19292 11854 19304
rect 12158 19292 12164 19304
rect 11848 19264 12164 19292
rect 11848 19252 11854 19264
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 11882 19224 11888 19236
rect 9416 19196 11888 19224
rect 9416 19168 9444 19196
rect 11882 19184 11888 19196
rect 11940 19224 11946 19236
rect 11940 19196 12112 19224
rect 11940 19184 11946 19196
rect 9263 19128 9352 19156
rect 9263 19125 9275 19128
rect 9217 19119 9275 19125
rect 9398 19116 9404 19168
rect 9456 19116 9462 19168
rect 9766 19116 9772 19168
rect 9824 19156 9830 19168
rect 9950 19156 9956 19168
rect 9824 19128 9956 19156
rect 9824 19116 9830 19128
rect 9950 19116 9956 19128
rect 10008 19156 10014 19168
rect 10045 19159 10103 19165
rect 10045 19156 10057 19159
rect 10008 19128 10057 19156
rect 10008 19116 10014 19128
rect 10045 19125 10057 19128
rect 10091 19125 10103 19159
rect 10045 19119 10103 19125
rect 11330 19116 11336 19168
rect 11388 19116 11394 19168
rect 11422 19116 11428 19168
rect 11480 19156 11486 19168
rect 11974 19156 11980 19168
rect 11480 19128 11980 19156
rect 11480 19116 11486 19128
rect 11974 19116 11980 19128
rect 12032 19116 12038 19168
rect 12084 19156 12112 19196
rect 12452 19156 12480 19400
rect 14277 19397 14289 19431
rect 14323 19428 14335 19431
rect 14323 19400 14412 19428
rect 14323 19397 14335 19400
rect 14277 19391 14335 19397
rect 14384 19360 14412 19400
rect 14458 19360 14464 19372
rect 14384 19332 14464 19360
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 15120 19332 15332 19360
rect 12526 19252 12532 19304
rect 12584 19252 12590 19304
rect 14645 19295 14703 19301
rect 14645 19261 14657 19295
rect 14691 19292 14703 19295
rect 14734 19292 14740 19304
rect 14691 19264 14740 19292
rect 14691 19261 14703 19264
rect 14645 19255 14703 19261
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 15120 19292 15148 19332
rect 15028 19264 15148 19292
rect 15304 19292 15332 19332
rect 16684 19332 16896 19360
rect 15381 19295 15439 19301
rect 15381 19292 15393 19295
rect 15304 19264 15393 19292
rect 12802 19184 12808 19236
rect 12860 19184 12866 19236
rect 14090 19224 14096 19236
rect 14030 19196 14096 19224
rect 14090 19184 14096 19196
rect 14148 19184 14154 19236
rect 15028 19168 15056 19264
rect 15381 19261 15393 19264
rect 15427 19261 15439 19295
rect 15381 19255 15439 19261
rect 15565 19295 15623 19301
rect 15565 19261 15577 19295
rect 15611 19292 15623 19295
rect 16684 19292 16712 19332
rect 16868 19304 16896 19332
rect 16960 19332 17172 19360
rect 15611 19264 16712 19292
rect 15611 19261 15623 19264
rect 15565 19255 15623 19261
rect 16758 19252 16764 19304
rect 16816 19252 16822 19304
rect 16850 19252 16856 19304
rect 16908 19252 16914 19304
rect 15194 19184 15200 19236
rect 15252 19224 15258 19236
rect 15746 19224 15752 19236
rect 15252 19196 15752 19224
rect 15252 19184 15258 19196
rect 15746 19184 15752 19196
rect 15804 19224 15810 19236
rect 16960 19224 16988 19332
rect 17029 19297 17087 19303
rect 17144 19301 17172 19332
rect 17029 19263 17041 19297
rect 17075 19263 17087 19297
rect 17029 19257 17087 19263
rect 17118 19295 17176 19301
rect 17118 19261 17130 19295
rect 17164 19261 17176 19295
rect 15804 19196 16988 19224
rect 15804 19184 15810 19196
rect 12084 19128 12480 19156
rect 14722 19116 14728 19168
rect 14780 19156 14786 19168
rect 14829 19159 14887 19165
rect 14829 19156 14841 19159
rect 14780 19128 14841 19156
rect 14780 19116 14786 19128
rect 14829 19125 14841 19128
rect 14875 19125 14887 19159
rect 14829 19119 14887 19125
rect 15010 19116 15016 19168
rect 15068 19116 15074 19168
rect 15286 19116 15292 19168
rect 15344 19116 15350 19168
rect 15565 19159 15623 19165
rect 15565 19125 15577 19159
rect 15611 19156 15623 19159
rect 16022 19156 16028 19168
rect 15611 19128 16028 19156
rect 15611 19125 15623 19128
rect 15565 19119 15623 19125
rect 16022 19116 16028 19128
rect 16080 19116 16086 19168
rect 16114 19116 16120 19168
rect 16172 19116 16178 19168
rect 16942 19116 16948 19168
rect 17000 19116 17006 19168
rect 17052 19156 17080 19257
rect 17118 19255 17176 19261
rect 18414 19252 18420 19304
rect 18472 19292 18478 19304
rect 18616 19292 18644 19468
rect 19794 19456 19800 19508
rect 19852 19496 19858 19508
rect 21637 19499 21695 19505
rect 19852 19468 20576 19496
rect 19852 19456 19858 19468
rect 19981 19431 20039 19437
rect 19981 19397 19993 19431
rect 20027 19397 20039 19431
rect 19981 19391 20039 19397
rect 19889 19295 19947 19301
rect 18472 19264 18538 19292
rect 18616 19264 19288 19292
rect 18472 19252 18478 19264
rect 17402 19184 17408 19236
rect 17460 19184 17466 19236
rect 19150 19184 19156 19236
rect 19208 19184 19214 19236
rect 19260 19224 19288 19264
rect 19889 19261 19901 19295
rect 19935 19292 19947 19295
rect 19996 19292 20024 19391
rect 20548 19369 20576 19468
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 21726 19496 21732 19508
rect 21683 19468 21732 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 21726 19456 21732 19468
rect 21784 19456 21790 19508
rect 22738 19456 22744 19508
rect 22796 19496 22802 19508
rect 22796 19468 23336 19496
rect 22796 19456 22802 19468
rect 23308 19428 23336 19468
rect 23658 19456 23664 19508
rect 23716 19496 23722 19508
rect 23937 19499 23995 19505
rect 23937 19496 23949 19499
rect 23716 19468 23949 19496
rect 23716 19456 23722 19468
rect 23937 19465 23949 19468
rect 23983 19465 23995 19499
rect 23937 19459 23995 19465
rect 24026 19456 24032 19508
rect 24084 19496 24090 19508
rect 24121 19499 24179 19505
rect 24121 19496 24133 19499
rect 24084 19468 24133 19496
rect 24084 19456 24090 19468
rect 24121 19465 24133 19468
rect 24167 19496 24179 19499
rect 24578 19496 24584 19508
rect 24167 19468 24584 19496
rect 24167 19465 24179 19468
rect 24121 19459 24179 19465
rect 24578 19456 24584 19468
rect 24636 19456 24642 19508
rect 24670 19456 24676 19508
rect 24728 19456 24734 19508
rect 24762 19456 24768 19508
rect 24820 19496 24826 19508
rect 26237 19499 26295 19505
rect 26237 19496 26249 19499
rect 24820 19468 26249 19496
rect 24820 19456 24826 19468
rect 26237 19465 26249 19468
rect 26283 19465 26295 19499
rect 26237 19459 26295 19465
rect 26326 19456 26332 19508
rect 26384 19496 26390 19508
rect 26384 19468 26464 19496
rect 26384 19456 26390 19468
rect 23308 19400 24072 19428
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 20622 19360 20628 19372
rect 20579 19332 20628 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 23109 19363 23167 19369
rect 23109 19329 23121 19363
rect 23155 19360 23167 19363
rect 23474 19360 23480 19372
rect 23155 19332 23480 19360
rect 23155 19329 23167 19332
rect 23109 19323 23167 19329
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 24044 19369 24072 19400
rect 24029 19363 24087 19369
rect 24029 19329 24041 19363
rect 24075 19360 24087 19363
rect 24688 19360 24716 19456
rect 25498 19388 25504 19440
rect 25556 19428 25562 19440
rect 26436 19428 26464 19468
rect 26602 19456 26608 19508
rect 26660 19496 26666 19508
rect 27525 19499 27583 19505
rect 27525 19496 27537 19499
rect 26660 19468 27537 19496
rect 26660 19456 26666 19468
rect 27525 19465 27537 19468
rect 27571 19465 27583 19499
rect 27525 19459 27583 19465
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 28537 19499 28595 19505
rect 28537 19496 28549 19499
rect 28132 19468 28549 19496
rect 28132 19456 28138 19468
rect 28537 19465 28549 19468
rect 28583 19465 28595 19499
rect 28537 19459 28595 19465
rect 28902 19456 28908 19508
rect 28960 19456 28966 19508
rect 25556 19400 26372 19428
rect 26436 19400 27752 19428
rect 25556 19388 25562 19400
rect 25958 19360 25964 19372
rect 24075 19332 24716 19360
rect 24872 19332 25964 19360
rect 24075 19329 24087 19332
rect 24029 19323 24087 19329
rect 19935 19264 20024 19292
rect 20349 19295 20407 19301
rect 19935 19261 19947 19264
rect 19889 19255 19947 19261
rect 20349 19261 20361 19295
rect 20395 19292 20407 19295
rect 23385 19295 23443 19301
rect 20395 19264 21588 19292
rect 20395 19261 20407 19264
rect 20349 19255 20407 19261
rect 19260 19196 20576 19224
rect 18046 19156 18052 19168
rect 17052 19128 18052 19156
rect 18046 19116 18052 19128
rect 18104 19116 18110 19168
rect 19242 19116 19248 19168
rect 19300 19116 19306 19168
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 20441 19159 20499 19165
rect 20441 19156 20453 19159
rect 20404 19128 20453 19156
rect 20404 19116 20410 19128
rect 20441 19125 20453 19128
rect 20487 19125 20499 19159
rect 20548 19156 20576 19196
rect 20898 19184 20904 19236
rect 20956 19224 20962 19236
rect 21085 19227 21143 19233
rect 21085 19224 21097 19227
rect 20956 19196 21097 19224
rect 20956 19184 20962 19196
rect 21085 19193 21097 19196
rect 21131 19224 21143 19227
rect 21453 19227 21511 19233
rect 21453 19224 21465 19227
rect 21131 19196 21465 19224
rect 21131 19193 21143 19196
rect 21085 19187 21143 19193
rect 21453 19193 21465 19196
rect 21499 19193 21511 19227
rect 21453 19187 21511 19193
rect 21560 19168 21588 19264
rect 23385 19261 23397 19295
rect 23431 19292 23443 19295
rect 23750 19292 23756 19304
rect 23431 19264 23756 19292
rect 23431 19261 23443 19264
rect 23385 19255 23443 19261
rect 23750 19252 23756 19264
rect 23808 19252 23814 19304
rect 23845 19295 23903 19301
rect 23845 19261 23857 19295
rect 23891 19261 23903 19295
rect 23845 19255 23903 19261
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 24872 19292 24900 19332
rect 25958 19320 25964 19332
rect 26016 19320 26022 19372
rect 26344 19369 26372 19400
rect 26329 19363 26387 19369
rect 26329 19329 26341 19363
rect 26375 19329 26387 19363
rect 26329 19323 26387 19329
rect 26528 19332 26740 19360
rect 24351 19264 24900 19292
rect 24949 19295 25007 19301
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 24949 19261 24961 19295
rect 24995 19261 25007 19295
rect 24949 19255 25007 19261
rect 25133 19295 25191 19301
rect 25133 19261 25145 19295
rect 25179 19261 25191 19295
rect 25133 19255 25191 19261
rect 22646 19184 22652 19236
rect 22704 19184 22710 19236
rect 23860 19224 23888 19255
rect 24964 19224 24992 19255
rect 23492 19196 23888 19224
rect 24320 19196 24992 19224
rect 21266 19156 21272 19168
rect 20548 19128 21272 19156
rect 20441 19119 20499 19125
rect 21266 19116 21272 19128
rect 21324 19156 21330 19168
rect 21361 19159 21419 19165
rect 21361 19156 21373 19159
rect 21324 19128 21373 19156
rect 21324 19116 21330 19128
rect 21361 19125 21373 19128
rect 21407 19125 21419 19159
rect 21361 19119 21419 19125
rect 21542 19116 21548 19168
rect 21600 19156 21606 19168
rect 23492 19156 23520 19196
rect 21600 19128 23520 19156
rect 23569 19159 23627 19165
rect 21600 19116 21606 19128
rect 23569 19125 23581 19159
rect 23615 19156 23627 19159
rect 24320 19156 24348 19196
rect 23615 19128 24348 19156
rect 23615 19125 23627 19128
rect 23569 19119 23627 19125
rect 24394 19116 24400 19168
rect 24452 19116 24458 19168
rect 24578 19116 24584 19168
rect 24636 19156 24642 19168
rect 25148 19156 25176 19255
rect 25406 19252 25412 19304
rect 25464 19292 25470 19304
rect 26528 19292 26556 19332
rect 25464 19264 26556 19292
rect 26605 19295 26663 19301
rect 25464 19252 25470 19264
rect 26605 19261 26617 19295
rect 26651 19261 26663 19295
rect 26712 19292 26740 19332
rect 27246 19320 27252 19372
rect 27304 19360 27310 19372
rect 27724 19369 27752 19400
rect 27709 19363 27767 19369
rect 27304 19332 27568 19360
rect 27304 19320 27310 19332
rect 26712 19264 27292 19292
rect 26605 19255 26663 19261
rect 26620 19224 26648 19255
rect 25792 19196 26648 19224
rect 27264 19224 27292 19264
rect 27430 19252 27436 19304
rect 27488 19252 27494 19304
rect 27540 19292 27568 19332
rect 27709 19329 27721 19363
rect 27755 19329 27767 19363
rect 27709 19323 27767 19329
rect 27798 19320 27804 19372
rect 27856 19320 27862 19372
rect 27890 19320 27896 19372
rect 27948 19320 27954 19372
rect 27985 19363 28043 19369
rect 27985 19329 27997 19363
rect 28031 19360 28043 19363
rect 28258 19360 28264 19372
rect 28031 19332 28264 19360
rect 28031 19329 28043 19332
rect 27985 19323 28043 19329
rect 28258 19320 28264 19332
rect 28316 19320 28322 19372
rect 28169 19295 28227 19301
rect 28169 19292 28181 19295
rect 27540 19286 27844 19292
rect 27908 19286 28181 19292
rect 27540 19264 28181 19286
rect 27816 19258 27936 19264
rect 28169 19261 28181 19264
rect 28215 19261 28227 19295
rect 28169 19255 28227 19261
rect 28353 19295 28411 19301
rect 28353 19261 28365 19295
rect 28399 19261 28411 19295
rect 28353 19255 28411 19261
rect 28629 19295 28687 19301
rect 28629 19261 28641 19295
rect 28675 19292 28687 19295
rect 28718 19292 28724 19304
rect 28675 19264 28724 19292
rect 28675 19261 28687 19264
rect 28629 19255 28687 19261
rect 27706 19224 27712 19236
rect 27264 19196 27712 19224
rect 25792 19168 25820 19196
rect 24636 19128 25176 19156
rect 24636 19116 24642 19128
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 25866 19116 25872 19168
rect 25924 19156 25930 19168
rect 27264 19165 27292 19196
rect 27706 19184 27712 19196
rect 27764 19184 27770 19236
rect 28368 19224 28396 19255
rect 27908 19196 28396 19224
rect 26053 19159 26111 19165
rect 26053 19156 26065 19159
rect 25924 19128 26065 19156
rect 25924 19116 25930 19128
rect 26053 19125 26065 19128
rect 26099 19125 26111 19159
rect 26053 19119 26111 19125
rect 27249 19159 27307 19165
rect 27249 19125 27261 19159
rect 27295 19125 27307 19159
rect 27249 19119 27307 19125
rect 27338 19116 27344 19168
rect 27396 19156 27402 19168
rect 27908 19156 27936 19196
rect 27396 19128 27936 19156
rect 27396 19116 27402 19128
rect 27982 19116 27988 19168
rect 28040 19156 28046 19168
rect 28169 19159 28227 19165
rect 28169 19156 28181 19159
rect 28040 19128 28181 19156
rect 28040 19116 28046 19128
rect 28169 19125 28181 19128
rect 28215 19125 28227 19159
rect 28169 19119 28227 19125
rect 28350 19116 28356 19168
rect 28408 19156 28414 19168
rect 28644 19156 28672 19255
rect 28718 19252 28724 19264
rect 28776 19252 28782 19304
rect 29273 19295 29331 19301
rect 29273 19261 29285 19295
rect 29319 19261 29331 19295
rect 29273 19255 29331 19261
rect 31757 19295 31815 19301
rect 31757 19261 31769 19295
rect 31803 19261 31815 19295
rect 31757 19255 31815 19261
rect 29288 19224 29316 19255
rect 29288 19196 29408 19224
rect 29380 19168 29408 19196
rect 29546 19184 29552 19236
rect 29604 19184 29610 19236
rect 30282 19184 30288 19236
rect 30340 19184 30346 19236
rect 31772 19224 31800 19255
rect 31036 19196 31800 19224
rect 31036 19168 31064 19196
rect 28408 19128 28672 19156
rect 28408 19116 28414 19128
rect 29362 19116 29368 19168
rect 29420 19116 29426 19168
rect 31018 19116 31024 19168
rect 31076 19116 31082 19168
rect 31202 19116 31208 19168
rect 31260 19116 31266 19168
rect 2760 19066 32200 19088
rect 2760 19014 6946 19066
rect 6998 19014 7010 19066
rect 7062 19014 7074 19066
rect 7126 19014 7138 19066
rect 7190 19014 7202 19066
rect 7254 19014 14306 19066
rect 14358 19014 14370 19066
rect 14422 19014 14434 19066
rect 14486 19014 14498 19066
rect 14550 19014 14562 19066
rect 14614 19014 21666 19066
rect 21718 19014 21730 19066
rect 21782 19014 21794 19066
rect 21846 19014 21858 19066
rect 21910 19014 21922 19066
rect 21974 19014 29026 19066
rect 29078 19014 29090 19066
rect 29142 19014 29154 19066
rect 29206 19014 29218 19066
rect 29270 19014 29282 19066
rect 29334 19014 32200 19066
rect 2760 18992 32200 19014
rect 7837 18955 7895 18961
rect 7837 18921 7849 18955
rect 7883 18952 7895 18955
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 7883 18924 8493 18952
rect 7883 18921 7895 18924
rect 7837 18915 7895 18921
rect 8481 18921 8493 18924
rect 8527 18952 8539 18955
rect 9769 18955 9827 18961
rect 8527 18924 9168 18952
rect 8527 18921 8539 18924
rect 8481 18915 8539 18921
rect 8938 18844 8944 18896
rect 8996 18884 9002 18896
rect 9033 18887 9091 18893
rect 9033 18884 9045 18887
rect 8996 18856 9045 18884
rect 8996 18844 9002 18856
rect 9033 18853 9045 18856
rect 9079 18853 9091 18887
rect 9140 18884 9168 18924
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 9815 18924 10088 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 9858 18884 9864 18896
rect 9140 18856 9864 18884
rect 9033 18847 9091 18853
rect 9858 18844 9864 18856
rect 9916 18844 9922 18896
rect 10060 18884 10088 18924
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13173 18955 13231 18961
rect 13173 18952 13185 18955
rect 12860 18924 13185 18952
rect 12860 18912 12866 18924
rect 13173 18921 13185 18924
rect 13219 18921 13231 18955
rect 13173 18915 13231 18921
rect 13633 18955 13691 18961
rect 13633 18921 13645 18955
rect 13679 18952 13691 18955
rect 13814 18952 13820 18964
rect 13679 18924 13820 18952
rect 13679 18921 13691 18924
rect 13633 18915 13691 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 14090 18912 14096 18964
rect 14148 18952 14154 18964
rect 14461 18955 14519 18961
rect 14461 18952 14473 18955
rect 14148 18924 14473 18952
rect 14148 18912 14154 18924
rect 14461 18921 14473 18924
rect 14507 18921 14519 18955
rect 14461 18915 14519 18921
rect 14550 18912 14556 18964
rect 14608 18952 14614 18964
rect 14734 18952 14740 18964
rect 14608 18924 14740 18952
rect 14608 18912 14614 18924
rect 14734 18912 14740 18924
rect 14792 18912 14798 18964
rect 15286 18912 15292 18964
rect 15344 18912 15350 18964
rect 17313 18955 17371 18961
rect 17313 18921 17325 18955
rect 17359 18952 17371 18955
rect 17402 18952 17408 18964
rect 17359 18924 17408 18952
rect 17359 18921 17371 18924
rect 17313 18915 17371 18921
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 17586 18912 17592 18964
rect 17644 18952 17650 18964
rect 17644 18924 21404 18952
rect 17644 18912 17650 18924
rect 10060 18856 11744 18884
rect 6086 18776 6092 18828
rect 6144 18776 6150 18828
rect 8573 18819 8631 18825
rect 8573 18785 8585 18819
rect 8619 18816 8631 18819
rect 9585 18819 9643 18825
rect 9585 18816 9597 18819
rect 8619 18788 9597 18816
rect 8619 18785 8631 18788
rect 8573 18779 8631 18785
rect 9585 18785 9597 18788
rect 9631 18816 9643 18819
rect 9674 18816 9680 18828
rect 9631 18788 9680 18816
rect 9631 18785 9643 18788
rect 9585 18779 9643 18785
rect 9674 18776 9680 18788
rect 9732 18776 9738 18828
rect 10873 18819 10931 18825
rect 10873 18785 10885 18819
rect 10919 18816 10931 18819
rect 10962 18816 10968 18828
rect 10919 18788 10968 18816
rect 10919 18785 10931 18788
rect 10873 18779 10931 18785
rect 10962 18776 10968 18788
rect 11020 18776 11026 18828
rect 4706 18708 4712 18760
rect 4764 18708 4770 18760
rect 4982 18708 4988 18760
rect 5040 18708 5046 18760
rect 7101 18751 7159 18757
rect 7101 18748 7113 18751
rect 6656 18720 7113 18748
rect 4724 18612 4752 18708
rect 6178 18640 6184 18692
rect 6236 18680 6242 18692
rect 6549 18683 6607 18689
rect 6549 18680 6561 18683
rect 6236 18652 6561 18680
rect 6236 18640 6242 18652
rect 6549 18649 6561 18652
rect 6595 18649 6607 18683
rect 6549 18643 6607 18649
rect 5166 18612 5172 18624
rect 4724 18584 5172 18612
rect 5166 18572 5172 18584
rect 5224 18572 5230 18624
rect 5994 18572 6000 18624
rect 6052 18612 6058 18624
rect 6457 18615 6515 18621
rect 6457 18612 6469 18615
rect 6052 18584 6469 18612
rect 6052 18572 6058 18584
rect 6457 18581 6469 18584
rect 6503 18612 6515 18615
rect 6656 18612 6684 18720
rect 7101 18717 7113 18720
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 7926 18708 7932 18760
rect 7984 18748 7990 18760
rect 8757 18751 8815 18757
rect 8757 18748 8769 18751
rect 7984 18720 8769 18748
rect 7984 18708 7990 18720
rect 8757 18717 8769 18720
rect 8803 18748 8815 18751
rect 9493 18751 9551 18757
rect 8803 18720 9168 18748
rect 8803 18717 8815 18720
rect 8757 18711 8815 18717
rect 8846 18640 8852 18692
rect 8904 18680 8910 18692
rect 9033 18683 9091 18689
rect 9033 18680 9045 18683
rect 8904 18652 9045 18680
rect 8904 18640 8910 18652
rect 9033 18649 9045 18652
rect 9079 18649 9091 18683
rect 9140 18680 9168 18720
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 9766 18748 9772 18760
rect 9539 18720 9772 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 9858 18708 9864 18760
rect 9916 18708 9922 18760
rect 10042 18708 10048 18760
rect 10100 18708 10106 18760
rect 11716 18748 11744 18856
rect 12526 18844 12532 18896
rect 12584 18884 12590 18896
rect 13446 18884 13452 18896
rect 12584 18856 13452 18884
rect 12584 18844 12590 18856
rect 13446 18844 13452 18856
rect 13504 18884 13510 18896
rect 15304 18884 15332 18912
rect 15746 18884 15752 18896
rect 13504 18856 15231 18884
rect 15304 18856 15752 18884
rect 13504 18844 13510 18856
rect 15203 18828 15231 18856
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 16942 18884 16948 18896
rect 16698 18856 16948 18884
rect 16942 18844 16948 18856
rect 17000 18844 17006 18896
rect 19242 18844 19248 18896
rect 19300 18884 19306 18896
rect 19613 18887 19671 18893
rect 19613 18884 19625 18887
rect 19300 18856 19625 18884
rect 19300 18844 19306 18856
rect 19613 18853 19625 18856
rect 19659 18853 19671 18887
rect 21082 18884 21088 18896
rect 20838 18856 21088 18884
rect 19613 18847 19671 18853
rect 21082 18844 21088 18856
rect 21140 18844 21146 18896
rect 12066 18776 12072 18828
rect 12124 18776 12130 18828
rect 12894 18816 12900 18828
rect 12544 18788 12900 18816
rect 12544 18757 12572 18788
rect 12894 18776 12900 18788
rect 12952 18776 12958 18828
rect 13354 18776 13360 18828
rect 13412 18816 13418 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 13412 18788 13553 18816
rect 13412 18776 13418 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 14093 18819 14151 18825
rect 14093 18785 14105 18819
rect 14139 18816 14151 18819
rect 14182 18816 14188 18828
rect 14139 18788 14188 18816
rect 14139 18785 14151 18788
rect 14093 18779 14151 18785
rect 14182 18776 14188 18788
rect 14240 18776 14246 18828
rect 15010 18816 15016 18828
rect 14292 18788 15016 18816
rect 12529 18751 12587 18757
rect 12529 18748 12541 18751
rect 11716 18720 12541 18748
rect 12529 18717 12541 18720
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 12618 18708 12624 18760
rect 12676 18708 12682 18760
rect 12986 18708 12992 18760
rect 13044 18708 13050 18760
rect 13446 18708 13452 18760
rect 13504 18748 13510 18760
rect 13725 18751 13783 18757
rect 13725 18748 13737 18751
rect 13504 18720 13737 18748
rect 13504 18708 13510 18720
rect 13725 18717 13737 18720
rect 13771 18717 13783 18751
rect 14292 18748 14320 18788
rect 15010 18776 15016 18788
rect 15068 18776 15074 18828
rect 15194 18776 15200 18828
rect 15252 18776 15258 18828
rect 17681 18819 17739 18825
rect 17681 18785 17693 18819
rect 17727 18816 17739 18819
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 17727 18788 18429 18816
rect 17727 18785 17739 18788
rect 17681 18779 17739 18785
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 13725 18711 13783 18717
rect 14108 18720 14320 18748
rect 14369 18751 14427 18757
rect 10060 18680 10088 18708
rect 9140 18652 10088 18680
rect 9033 18643 9091 18649
rect 6503 18584 6684 18612
rect 6503 18581 6515 18584
rect 6457 18575 6515 18581
rect 8110 18572 8116 18624
rect 8168 18572 8174 18624
rect 9048 18612 9076 18643
rect 10134 18640 10140 18692
rect 10192 18640 10198 18692
rect 12161 18683 12219 18689
rect 12161 18649 12173 18683
rect 12207 18680 12219 18683
rect 12207 18652 13124 18680
rect 12207 18649 12219 18652
rect 12161 18643 12219 18649
rect 10152 18612 10180 18640
rect 13096 18624 13124 18652
rect 14108 18624 14136 18720
rect 14369 18717 14381 18751
rect 14415 18748 14427 18751
rect 14415 18720 15341 18748
rect 14415 18717 14427 18720
rect 14369 18711 14427 18717
rect 14185 18683 14243 18689
rect 14185 18649 14197 18683
rect 14231 18680 14243 18683
rect 14274 18680 14280 18692
rect 14231 18652 14280 18680
rect 14231 18649 14243 18652
rect 14185 18643 14243 18649
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 9048 18584 10180 18612
rect 10502 18572 10508 18624
rect 10560 18572 10566 18624
rect 12345 18615 12403 18621
rect 12345 18581 12357 18615
rect 12391 18612 12403 18615
rect 12434 18612 12440 18624
rect 12391 18584 12440 18612
rect 12391 18581 12403 18584
rect 12345 18575 12403 18581
rect 12434 18572 12440 18584
rect 12492 18572 12498 18624
rect 13078 18572 13084 18624
rect 13136 18572 13142 18624
rect 14090 18572 14096 18624
rect 14148 18572 14154 18624
rect 15313 18612 15341 18720
rect 15470 18708 15476 18760
rect 15528 18708 15534 18760
rect 16942 18708 16948 18760
rect 17000 18748 17006 18760
rect 17770 18748 17776 18760
rect 17000 18720 17776 18748
rect 17000 18708 17006 18720
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 17862 18708 17868 18760
rect 17920 18708 17926 18760
rect 19061 18751 19119 18757
rect 19061 18717 19073 18751
rect 19107 18748 19119 18751
rect 19150 18748 19156 18760
rect 19107 18720 19156 18748
rect 19107 18717 19119 18720
rect 19061 18711 19119 18717
rect 19150 18708 19156 18720
rect 19208 18708 19214 18760
rect 19334 18708 19340 18760
rect 19392 18708 19398 18760
rect 20346 18748 20352 18760
rect 19444 18720 20352 18748
rect 16482 18640 16488 18692
rect 16540 18680 16546 18692
rect 16540 18652 17080 18680
rect 16540 18640 16546 18652
rect 16114 18612 16120 18624
rect 15313 18584 16120 18612
rect 16114 18572 16120 18584
rect 16172 18572 16178 18624
rect 16758 18572 16764 18624
rect 16816 18612 16822 18624
rect 16945 18615 17003 18621
rect 16945 18612 16957 18615
rect 16816 18584 16957 18612
rect 16816 18572 16822 18584
rect 16945 18581 16957 18584
rect 16991 18581 17003 18615
rect 17052 18612 17080 18652
rect 18506 18640 18512 18692
rect 18564 18680 18570 18692
rect 19444 18680 19472 18720
rect 20346 18708 20352 18720
rect 20404 18748 20410 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20404 18720 21097 18748
rect 20404 18708 20410 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 18564 18652 19472 18680
rect 21376 18680 21404 18924
rect 22646 18912 22652 18964
rect 22704 18912 22710 18964
rect 23201 18955 23259 18961
rect 23201 18921 23213 18955
rect 23247 18952 23259 18955
rect 23382 18952 23388 18964
rect 23247 18924 23388 18952
rect 23247 18921 23259 18924
rect 23201 18915 23259 18921
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 23842 18952 23848 18964
rect 23492 18924 23848 18952
rect 23492 18884 23520 18924
rect 23842 18912 23848 18924
rect 23900 18912 23906 18964
rect 24118 18912 24124 18964
rect 24176 18952 24182 18964
rect 24673 18955 24731 18961
rect 24673 18952 24685 18955
rect 24176 18924 24685 18952
rect 24176 18912 24182 18924
rect 24673 18921 24685 18924
rect 24719 18921 24731 18955
rect 26418 18952 26424 18964
rect 24673 18915 24731 18921
rect 24872 18924 26424 18952
rect 23124 18856 23520 18884
rect 21637 18819 21695 18825
rect 21637 18785 21649 18819
rect 21683 18816 21695 18819
rect 22738 18816 22744 18828
rect 21683 18788 22744 18816
rect 21683 18785 21695 18788
rect 21637 18779 21695 18785
rect 21450 18708 21456 18760
rect 21508 18748 21514 18760
rect 21652 18748 21680 18779
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 23124 18825 23152 18856
rect 23750 18844 23756 18896
rect 23808 18884 23814 18896
rect 24872 18884 24900 18924
rect 26418 18912 26424 18924
rect 26476 18912 26482 18964
rect 26510 18912 26516 18964
rect 26568 18952 26574 18964
rect 27798 18952 27804 18964
rect 26568 18924 27804 18952
rect 26568 18912 26574 18924
rect 27798 18912 27804 18924
rect 27856 18912 27862 18964
rect 29365 18955 29423 18961
rect 29365 18921 29377 18955
rect 29411 18952 29423 18955
rect 29546 18952 29552 18964
rect 29411 18924 29552 18952
rect 29411 18921 29423 18924
rect 29365 18915 29423 18921
rect 29546 18912 29552 18924
rect 29604 18912 29610 18964
rect 30282 18912 30288 18964
rect 30340 18912 30346 18964
rect 31202 18912 31208 18964
rect 31260 18912 31266 18964
rect 23808 18856 24900 18884
rect 23808 18844 23814 18856
rect 23109 18819 23167 18825
rect 23109 18785 23121 18819
rect 23155 18785 23167 18819
rect 23109 18779 23167 18785
rect 23293 18819 23351 18825
rect 23293 18785 23305 18819
rect 23339 18816 23351 18819
rect 24026 18816 24032 18828
rect 23339 18788 24032 18816
rect 23339 18785 23351 18788
rect 23293 18779 23351 18785
rect 24026 18776 24032 18788
rect 24084 18776 24090 18828
rect 24581 18819 24639 18825
rect 24581 18785 24593 18819
rect 24627 18816 24639 18819
rect 24670 18816 24676 18828
rect 24627 18788 24676 18816
rect 24627 18785 24639 18788
rect 24581 18779 24639 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 24762 18776 24768 18828
rect 24820 18776 24826 18828
rect 24872 18825 24900 18856
rect 25130 18844 25136 18896
rect 25188 18844 25194 18896
rect 25590 18844 25596 18896
rect 25648 18844 25654 18896
rect 26786 18844 26792 18896
rect 26844 18884 26850 18896
rect 29733 18887 29791 18893
rect 26844 18856 28948 18884
rect 26844 18844 26850 18856
rect 28920 18828 28948 18856
rect 29733 18853 29745 18887
rect 29779 18884 29791 18887
rect 31220 18884 31248 18912
rect 29779 18856 31248 18884
rect 31665 18887 31723 18893
rect 29779 18853 29791 18856
rect 29733 18847 29791 18853
rect 31665 18853 31677 18887
rect 31711 18884 31723 18887
rect 33134 18884 33140 18896
rect 31711 18856 33140 18884
rect 31711 18853 31723 18856
rect 31665 18847 31723 18853
rect 33134 18844 33140 18856
rect 33192 18844 33198 18896
rect 24857 18819 24915 18825
rect 24857 18785 24869 18819
rect 24903 18785 24915 18819
rect 28350 18816 28356 18828
rect 24857 18779 24915 18785
rect 26528 18788 28356 18816
rect 21508 18720 21680 18748
rect 24489 18751 24547 18757
rect 21508 18708 21514 18720
rect 24489 18717 24501 18751
rect 24535 18748 24547 18751
rect 25866 18748 25872 18760
rect 24535 18720 25872 18748
rect 24535 18717 24547 18720
rect 24489 18711 24547 18717
rect 25866 18708 25872 18720
rect 25924 18708 25930 18760
rect 26528 18748 26556 18788
rect 28350 18776 28356 18788
rect 28408 18776 28414 18828
rect 28902 18776 28908 18828
rect 28960 18776 28966 18828
rect 30190 18776 30196 18828
rect 30248 18776 30254 18828
rect 30653 18819 30711 18825
rect 30653 18785 30665 18819
rect 30699 18816 30711 18819
rect 31018 18816 31024 18828
rect 30699 18788 31024 18816
rect 30699 18785 30711 18788
rect 30653 18779 30711 18785
rect 31018 18776 31024 18788
rect 31076 18776 31082 18828
rect 26252 18720 26556 18748
rect 26605 18751 26663 18757
rect 26252 18692 26280 18720
rect 26605 18717 26617 18751
rect 26651 18748 26663 18751
rect 26881 18751 26939 18757
rect 26881 18748 26893 18751
rect 26651 18720 26893 18748
rect 26651 18717 26663 18720
rect 26605 18711 26663 18717
rect 26881 18717 26893 18720
rect 26927 18717 26939 18751
rect 27801 18751 27859 18757
rect 27801 18748 27813 18751
rect 26881 18711 26939 18717
rect 26988 18720 27813 18748
rect 26988 18692 27016 18720
rect 27801 18717 27813 18720
rect 27847 18717 27859 18751
rect 27801 18711 27859 18717
rect 29822 18708 29828 18760
rect 29880 18708 29886 18760
rect 29917 18751 29975 18757
rect 29917 18717 29929 18751
rect 29963 18717 29975 18751
rect 29917 18711 29975 18717
rect 21376 18652 24256 18680
rect 18564 18640 18570 18652
rect 20070 18612 20076 18624
rect 17052 18584 20076 18612
rect 16945 18575 17003 18581
rect 20070 18572 20076 18584
rect 20128 18572 20134 18624
rect 21082 18572 21088 18624
rect 21140 18612 21146 18624
rect 21545 18615 21603 18621
rect 21545 18612 21557 18615
rect 21140 18584 21557 18612
rect 21140 18572 21146 18584
rect 21545 18581 21557 18584
rect 21591 18581 21603 18615
rect 21545 18575 21603 18581
rect 23566 18572 23572 18624
rect 23624 18612 23630 18624
rect 23845 18615 23903 18621
rect 23845 18612 23857 18615
rect 23624 18584 23857 18612
rect 23624 18572 23630 18584
rect 23845 18581 23857 18584
rect 23891 18581 23903 18615
rect 24228 18612 24256 18652
rect 26234 18640 26240 18692
rect 26292 18640 26298 18692
rect 26970 18640 26976 18692
rect 27028 18640 27034 18692
rect 27522 18640 27528 18692
rect 27580 18640 27586 18692
rect 28902 18680 28908 18692
rect 27632 18652 28908 18680
rect 27632 18612 27660 18652
rect 28902 18640 28908 18652
rect 28960 18680 28966 18692
rect 29932 18680 29960 18711
rect 28960 18652 29960 18680
rect 28960 18640 28966 18652
rect 24228 18584 27660 18612
rect 23845 18575 23903 18581
rect 27890 18572 27896 18624
rect 27948 18612 27954 18624
rect 28261 18615 28319 18621
rect 28261 18612 28273 18615
rect 27948 18584 28273 18612
rect 27948 18572 27954 18584
rect 28261 18581 28273 18584
rect 28307 18581 28319 18615
rect 28261 18575 28319 18581
rect 28718 18572 28724 18624
rect 28776 18612 28782 18624
rect 28997 18615 29055 18621
rect 28997 18612 29009 18615
rect 28776 18584 29009 18612
rect 28776 18572 28782 18584
rect 28997 18581 29009 18584
rect 29043 18612 29055 18615
rect 29822 18612 29828 18624
rect 29043 18584 29828 18612
rect 29043 18581 29055 18584
rect 28997 18575 29055 18581
rect 29822 18572 29828 18584
rect 29880 18572 29886 18624
rect 2760 18522 32200 18544
rect 2760 18470 6286 18522
rect 6338 18470 6350 18522
rect 6402 18470 6414 18522
rect 6466 18470 6478 18522
rect 6530 18470 6542 18522
rect 6594 18470 13646 18522
rect 13698 18470 13710 18522
rect 13762 18470 13774 18522
rect 13826 18470 13838 18522
rect 13890 18470 13902 18522
rect 13954 18470 21006 18522
rect 21058 18470 21070 18522
rect 21122 18470 21134 18522
rect 21186 18470 21198 18522
rect 21250 18470 21262 18522
rect 21314 18470 28366 18522
rect 28418 18470 28430 18522
rect 28482 18470 28494 18522
rect 28546 18470 28558 18522
rect 28610 18470 28622 18522
rect 28674 18470 32200 18522
rect 2760 18448 32200 18470
rect 4982 18368 4988 18420
rect 5040 18408 5046 18420
rect 5445 18411 5503 18417
rect 5445 18408 5457 18411
rect 5040 18380 5457 18408
rect 5040 18368 5046 18380
rect 5445 18377 5457 18380
rect 5491 18377 5503 18411
rect 5445 18371 5503 18377
rect 6086 18368 6092 18420
rect 6144 18408 6150 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 6144 18380 6377 18408
rect 6144 18368 6150 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 6454 18368 6460 18420
rect 6512 18408 6518 18420
rect 6733 18411 6791 18417
rect 6733 18408 6745 18411
rect 6512 18380 6745 18408
rect 6512 18368 6518 18380
rect 6733 18377 6745 18380
rect 6779 18377 6791 18411
rect 6733 18371 6791 18377
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 8202 18408 8208 18420
rect 6972 18380 8208 18408
rect 6972 18368 6978 18380
rect 8202 18368 8208 18380
rect 8260 18368 8266 18420
rect 8376 18411 8434 18417
rect 8376 18377 8388 18411
rect 8422 18408 8434 18411
rect 8754 18408 8760 18420
rect 8422 18380 8760 18408
rect 8422 18377 8434 18380
rect 8376 18371 8434 18377
rect 8754 18368 8760 18380
rect 8812 18368 8818 18420
rect 9858 18368 9864 18420
rect 9916 18368 9922 18420
rect 11882 18368 11888 18420
rect 11940 18368 11946 18420
rect 12161 18411 12219 18417
rect 12161 18377 12173 18411
rect 12207 18408 12219 18411
rect 12986 18408 12992 18420
rect 12207 18380 12992 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 12986 18368 12992 18380
rect 13044 18408 13050 18420
rect 14093 18411 14151 18417
rect 13044 18380 13676 18408
rect 13044 18368 13050 18380
rect 5166 18300 5172 18352
rect 5224 18340 5230 18352
rect 5224 18312 7052 18340
rect 5224 18300 5230 18312
rect 5626 18232 5632 18284
rect 5684 18272 5690 18284
rect 5997 18275 6055 18281
rect 5997 18272 6009 18275
rect 5684 18244 6009 18272
rect 5684 18232 5690 18244
rect 5997 18241 6009 18244
rect 6043 18272 6055 18275
rect 6086 18272 6092 18284
rect 6043 18244 6092 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 6086 18232 6092 18244
rect 6144 18272 6150 18284
rect 6362 18272 6368 18284
rect 6144 18244 6368 18272
rect 6144 18232 6150 18244
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 6914 18272 6920 18284
rect 6472 18244 6920 18272
rect 5813 18207 5871 18213
rect 5813 18173 5825 18207
rect 5859 18204 5871 18207
rect 6178 18204 6184 18216
rect 5859 18176 6184 18204
rect 5859 18173 5871 18176
rect 5813 18167 5871 18173
rect 6178 18164 6184 18176
rect 6236 18164 6242 18216
rect 6472 18213 6500 18244
rect 6914 18232 6920 18244
rect 6972 18232 6978 18284
rect 6457 18207 6515 18213
rect 6457 18173 6469 18207
rect 6503 18173 6515 18207
rect 7024 18204 7052 18312
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 10597 18343 10655 18349
rect 10597 18340 10609 18343
rect 9732 18312 10609 18340
rect 9732 18300 9738 18312
rect 10597 18309 10609 18312
rect 10643 18309 10655 18343
rect 13648 18340 13676 18380
rect 14093 18377 14105 18411
rect 14139 18408 14151 18411
rect 14366 18408 14372 18420
rect 14139 18380 14372 18408
rect 14139 18377 14151 18380
rect 14093 18371 14151 18377
rect 14366 18368 14372 18380
rect 14424 18408 14430 18420
rect 14734 18408 14740 18420
rect 14424 18380 14740 18408
rect 14424 18368 14430 18380
rect 14734 18368 14740 18380
rect 14792 18368 14798 18420
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 15749 18411 15807 18417
rect 15749 18408 15761 18411
rect 15528 18380 15761 18408
rect 15528 18368 15534 18380
rect 15749 18377 15761 18380
rect 15795 18377 15807 18411
rect 15749 18371 15807 18377
rect 15838 18368 15844 18420
rect 15896 18408 15902 18420
rect 15896 18380 17264 18408
rect 15896 18368 15902 18380
rect 16482 18340 16488 18352
rect 13648 18312 16488 18340
rect 10597 18303 10655 18309
rect 16482 18300 16488 18312
rect 16540 18300 16546 18352
rect 16592 18312 17060 18340
rect 7926 18232 7932 18284
rect 7984 18232 7990 18284
rect 8386 18232 8392 18284
rect 8444 18272 8450 18284
rect 16592 18272 16620 18312
rect 8444 18244 16620 18272
rect 8444 18232 8450 18244
rect 8113 18207 8171 18213
rect 8113 18204 8125 18207
rect 7024 18176 8125 18204
rect 6457 18167 6515 18173
rect 8113 18173 8125 18176
rect 8159 18173 8171 18207
rect 8113 18167 8171 18173
rect 10042 18164 10048 18216
rect 10100 18204 10106 18216
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 10100 18176 10149 18204
rect 10100 18164 10106 18176
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18173 10471 18207
rect 10413 18167 10471 18173
rect 4062 18096 4068 18148
rect 4120 18136 4126 18148
rect 8386 18136 8392 18148
rect 4120 18108 8392 18136
rect 4120 18096 4126 18108
rect 8386 18096 8392 18108
rect 8444 18096 8450 18148
rect 9122 18096 9128 18148
rect 9180 18096 9186 18148
rect 10428 18136 10456 18167
rect 10594 18164 10600 18216
rect 10652 18204 10658 18216
rect 11149 18207 11207 18213
rect 11149 18204 11161 18207
rect 10652 18176 11161 18204
rect 10652 18164 10658 18176
rect 11149 18173 11161 18176
rect 11195 18173 11207 18207
rect 11149 18167 11207 18173
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 12253 18207 12311 18213
rect 12253 18173 12265 18207
rect 12299 18173 12311 18207
rect 12253 18167 12311 18173
rect 12345 18207 12403 18213
rect 12345 18173 12357 18207
rect 12391 18173 12403 18207
rect 12345 18167 12403 18173
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 14642 18204 14648 18216
rect 14323 18176 14648 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 10962 18136 10968 18148
rect 10428 18108 10968 18136
rect 10962 18096 10968 18108
rect 11020 18096 11026 18148
rect 12084 18080 12112 18167
rect 5905 18071 5963 18077
rect 5905 18037 5917 18071
rect 5951 18068 5963 18071
rect 7190 18068 7196 18080
rect 5951 18040 7196 18068
rect 5951 18037 5963 18040
rect 5905 18031 5963 18037
rect 7190 18028 7196 18040
rect 7248 18028 7254 18080
rect 7285 18071 7343 18077
rect 7285 18037 7297 18071
rect 7331 18068 7343 18071
rect 7374 18068 7380 18080
rect 7331 18040 7380 18068
rect 7331 18037 7343 18040
rect 7285 18031 7343 18037
rect 7374 18028 7380 18040
rect 7432 18028 7438 18080
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 7650 18068 7656 18080
rect 7524 18040 7656 18068
rect 7524 18028 7530 18040
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 7745 18071 7803 18077
rect 7745 18037 7757 18071
rect 7791 18068 7803 18071
rect 10134 18068 10140 18080
rect 7791 18040 10140 18068
rect 7791 18037 7803 18040
rect 7745 18031 7803 18037
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 11514 18028 11520 18080
rect 11572 18028 11578 18080
rect 12066 18028 12072 18080
rect 12124 18028 12130 18080
rect 12268 18068 12296 18167
rect 12360 18136 12388 18167
rect 14642 18164 14648 18176
rect 14700 18204 14706 18216
rect 14921 18207 14979 18213
rect 14921 18204 14933 18207
rect 14700 18176 14933 18204
rect 14700 18164 14706 18176
rect 14921 18173 14933 18176
rect 14967 18173 14979 18207
rect 15933 18207 15991 18213
rect 15933 18206 15945 18207
rect 14921 18167 14979 18173
rect 15672 18178 15945 18206
rect 12526 18136 12532 18148
rect 12360 18108 12532 18136
rect 12526 18096 12532 18108
rect 12584 18096 12590 18148
rect 12618 18096 12624 18148
rect 12676 18096 12682 18148
rect 13078 18096 13084 18148
rect 13136 18096 13142 18148
rect 15672 18136 15700 18178
rect 15933 18173 15945 18178
rect 15979 18173 15991 18207
rect 15933 18167 15991 18173
rect 16022 18164 16028 18216
rect 16080 18164 16086 18216
rect 16206 18164 16212 18216
rect 16264 18164 16270 18216
rect 16482 18164 16488 18216
rect 16540 18164 16546 18216
rect 16577 18207 16635 18213
rect 16577 18173 16589 18207
rect 16623 18173 16635 18207
rect 16577 18167 16635 18173
rect 16761 18207 16819 18213
rect 16761 18173 16773 18207
rect 16807 18173 16819 18207
rect 16761 18167 16819 18173
rect 13924 18108 15700 18136
rect 12710 18068 12716 18080
rect 12268 18040 12716 18068
rect 12710 18028 12716 18040
rect 12768 18028 12774 18080
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 13924 18068 13952 18108
rect 15838 18096 15844 18148
rect 15896 18096 15902 18148
rect 16224 18136 16252 18164
rect 16592 18136 16620 18167
rect 16224 18108 16620 18136
rect 13044 18040 13952 18068
rect 14829 18071 14887 18077
rect 13044 18028 13050 18040
rect 14829 18037 14841 18071
rect 14875 18068 14887 18071
rect 14918 18068 14924 18080
rect 14875 18040 14924 18068
rect 14875 18037 14887 18040
rect 14829 18031 14887 18037
rect 14918 18028 14924 18040
rect 14976 18028 14982 18080
rect 15565 18071 15623 18077
rect 15565 18037 15577 18071
rect 15611 18068 15623 18071
rect 15746 18068 15752 18080
rect 15611 18040 15752 18068
rect 15611 18037 15623 18040
rect 15565 18031 15623 18037
rect 15746 18028 15752 18040
rect 15804 18028 15810 18080
rect 15856 18068 15884 18096
rect 16390 18068 16396 18080
rect 15856 18040 16396 18068
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 16776 18068 16804 18167
rect 16850 18164 16856 18216
rect 16908 18164 16914 18216
rect 17032 18204 17060 18312
rect 17129 18207 17187 18213
rect 17129 18204 17141 18207
rect 17032 18176 17141 18204
rect 17129 18173 17141 18176
rect 17175 18173 17187 18207
rect 17236 18204 17264 18380
rect 17770 18368 17776 18420
rect 17828 18368 17834 18420
rect 18322 18368 18328 18420
rect 18380 18408 18386 18420
rect 20165 18411 20223 18417
rect 20165 18408 20177 18411
rect 18380 18380 20177 18408
rect 18380 18368 18386 18380
rect 20165 18377 20177 18380
rect 20211 18377 20223 18411
rect 20165 18371 20223 18377
rect 23474 18368 23480 18420
rect 23532 18368 23538 18420
rect 23658 18368 23664 18420
rect 23716 18408 23722 18420
rect 23842 18408 23848 18420
rect 23716 18380 23848 18408
rect 23716 18368 23722 18380
rect 23842 18368 23848 18380
rect 23900 18368 23906 18420
rect 23934 18368 23940 18420
rect 23992 18368 23998 18420
rect 24394 18368 24400 18420
rect 24452 18368 24458 18420
rect 24578 18368 24584 18420
rect 24636 18368 24642 18420
rect 25041 18411 25099 18417
rect 25041 18377 25053 18411
rect 25087 18408 25099 18411
rect 25590 18408 25596 18420
rect 25087 18380 25596 18408
rect 25087 18377 25099 18380
rect 25041 18371 25099 18377
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 25682 18368 25688 18420
rect 25740 18408 25746 18420
rect 25869 18411 25927 18417
rect 25869 18408 25881 18411
rect 25740 18380 25881 18408
rect 25740 18368 25746 18380
rect 25869 18377 25881 18380
rect 25915 18377 25927 18411
rect 25869 18371 25927 18377
rect 26421 18411 26479 18417
rect 26421 18377 26433 18411
rect 26467 18408 26479 18411
rect 26510 18408 26516 18420
rect 26467 18380 26516 18408
rect 26467 18377 26479 18380
rect 26421 18371 26479 18377
rect 26510 18368 26516 18380
rect 26568 18368 26574 18420
rect 27430 18368 27436 18420
rect 27488 18408 27494 18420
rect 28261 18411 28319 18417
rect 28261 18408 28273 18411
rect 27488 18380 28273 18408
rect 27488 18368 27494 18380
rect 28261 18377 28273 18380
rect 28307 18377 28319 18411
rect 28261 18371 28319 18377
rect 17788 18340 17816 18368
rect 18969 18343 19027 18349
rect 18969 18340 18981 18343
rect 17788 18312 18981 18340
rect 18969 18309 18981 18312
rect 19015 18309 19027 18343
rect 18969 18303 19027 18309
rect 19058 18300 19064 18352
rect 19116 18300 19122 18352
rect 19150 18300 19156 18352
rect 19208 18340 19214 18352
rect 19426 18340 19432 18352
rect 19208 18312 19432 18340
rect 19208 18300 19214 18312
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 21729 18343 21787 18349
rect 21729 18309 21741 18343
rect 21775 18340 21787 18343
rect 23952 18340 23980 18368
rect 21775 18312 22094 18340
rect 21775 18309 21787 18312
rect 21729 18303 21787 18309
rect 18877 18275 18935 18281
rect 18877 18241 18889 18275
rect 18923 18272 18935 18275
rect 19610 18272 19616 18284
rect 18923 18244 19616 18272
rect 18923 18241 18935 18244
rect 18877 18235 18935 18241
rect 19610 18232 19616 18244
rect 19668 18232 19674 18284
rect 20622 18232 20628 18284
rect 20680 18272 20686 18284
rect 21085 18275 21143 18281
rect 21085 18272 21097 18275
rect 20680 18244 21097 18272
rect 20680 18232 20686 18244
rect 21085 18241 21097 18244
rect 21131 18241 21143 18275
rect 22066 18272 22094 18312
rect 23676 18312 23980 18340
rect 23676 18281 23704 18312
rect 22373 18275 22431 18281
rect 22373 18272 22385 18275
rect 22066 18244 22385 18272
rect 21085 18235 21143 18241
rect 22373 18241 22385 18244
rect 22419 18241 22431 18275
rect 22373 18235 22431 18241
rect 23661 18275 23719 18281
rect 23661 18241 23673 18275
rect 23707 18241 23719 18275
rect 23661 18235 23719 18241
rect 23937 18275 23995 18281
rect 23937 18241 23949 18275
rect 23983 18272 23995 18275
rect 24412 18272 24440 18368
rect 27341 18343 27399 18349
rect 27341 18309 27353 18343
rect 27387 18340 27399 18343
rect 27387 18312 27476 18340
rect 27387 18309 27399 18312
rect 27341 18303 27399 18309
rect 26050 18272 26056 18284
rect 23983 18244 24440 18272
rect 24964 18244 26056 18272
rect 23983 18241 23995 18244
rect 23937 18235 23995 18241
rect 24964 18216 24992 18244
rect 26050 18232 26056 18244
rect 26108 18232 26114 18284
rect 26786 18232 26792 18284
rect 26844 18232 26850 18284
rect 26878 18232 26884 18284
rect 26936 18232 26942 18284
rect 27448 18281 27476 18312
rect 27433 18275 27491 18281
rect 27433 18241 27445 18275
rect 27479 18241 27491 18275
rect 27433 18235 27491 18241
rect 29181 18275 29239 18281
rect 29181 18241 29193 18275
rect 29227 18272 29239 18275
rect 30282 18272 30288 18284
rect 29227 18244 30288 18272
rect 29227 18241 29239 18244
rect 29181 18235 29239 18241
rect 30282 18232 30288 18244
rect 30340 18272 30346 18284
rect 30340 18244 30880 18272
rect 30340 18232 30346 18244
rect 19518 18204 19524 18216
rect 17236 18176 19524 18204
rect 17129 18167 17187 18173
rect 19518 18164 19524 18176
rect 19576 18164 19582 18216
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 19794 18204 19800 18216
rect 19751 18176 19800 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 19794 18164 19800 18176
rect 19852 18164 19858 18216
rect 19978 18164 19984 18216
rect 20036 18164 20042 18216
rect 20070 18164 20076 18216
rect 20128 18164 20134 18216
rect 20254 18164 20260 18216
rect 20312 18204 20318 18216
rect 20533 18207 20591 18213
rect 20533 18204 20545 18207
rect 20312 18176 20545 18204
rect 20312 18164 20318 18176
rect 20533 18173 20545 18176
rect 20579 18173 20591 18207
rect 20533 18167 20591 18173
rect 22554 18164 22560 18216
rect 22612 18164 22618 18216
rect 23753 18207 23811 18213
rect 23753 18173 23765 18207
rect 23799 18173 23811 18207
rect 23753 18167 23811 18173
rect 16868 18136 16896 18164
rect 16868 18108 17356 18136
rect 17328 18080 17356 18108
rect 19426 18096 19432 18148
rect 19484 18096 19490 18148
rect 19613 18139 19671 18145
rect 19613 18105 19625 18139
rect 19659 18136 19671 18139
rect 20346 18136 20352 18148
rect 19659 18108 20352 18136
rect 19659 18105 19671 18108
rect 19613 18099 19671 18105
rect 20346 18096 20352 18108
rect 20404 18096 20410 18148
rect 21361 18139 21419 18145
rect 21361 18105 21373 18139
rect 21407 18136 21419 18139
rect 22830 18136 22836 18148
rect 21407 18108 22836 18136
rect 21407 18105 21419 18108
rect 21361 18099 21419 18105
rect 22830 18096 22836 18108
rect 22888 18096 22894 18148
rect 16850 18068 16856 18080
rect 16776 18040 16856 18068
rect 16850 18028 16856 18040
rect 16908 18028 16914 18080
rect 17034 18028 17040 18080
rect 17092 18028 17098 18080
rect 17310 18028 17316 18080
rect 17368 18028 17374 18080
rect 19242 18028 19248 18080
rect 19300 18068 19306 18080
rect 19889 18071 19947 18077
rect 19889 18068 19901 18071
rect 19300 18040 19901 18068
rect 19300 18028 19306 18040
rect 19889 18037 19901 18040
rect 19935 18037 19947 18071
rect 19889 18031 19947 18037
rect 21266 18028 21272 18080
rect 21324 18028 21330 18080
rect 21821 18071 21879 18077
rect 21821 18037 21833 18071
rect 21867 18068 21879 18071
rect 22002 18068 22008 18080
rect 21867 18040 22008 18068
rect 21867 18037 21879 18040
rect 21821 18031 21879 18037
rect 22002 18028 22008 18040
rect 22060 18028 22066 18080
rect 23106 18028 23112 18080
rect 23164 18068 23170 18080
rect 23201 18071 23259 18077
rect 23201 18068 23213 18071
rect 23164 18040 23213 18068
rect 23164 18028 23170 18040
rect 23201 18037 23213 18040
rect 23247 18037 23259 18071
rect 23768 18068 23796 18167
rect 23842 18164 23848 18216
rect 23900 18164 23906 18216
rect 24397 18207 24455 18213
rect 24397 18173 24409 18207
rect 24443 18173 24455 18207
rect 24397 18167 24455 18173
rect 24412 18136 24440 18167
rect 24486 18164 24492 18216
rect 24544 18204 24550 18216
rect 24581 18207 24639 18213
rect 24581 18204 24593 18207
rect 24544 18176 24593 18204
rect 24544 18164 24550 18176
rect 24581 18173 24593 18176
rect 24627 18173 24639 18207
rect 24581 18167 24639 18173
rect 24946 18164 24952 18216
rect 25004 18164 25010 18216
rect 25314 18164 25320 18216
rect 25372 18164 25378 18216
rect 25958 18164 25964 18216
rect 26016 18204 26022 18216
rect 26237 18207 26295 18213
rect 26237 18204 26249 18207
rect 26016 18176 26249 18204
rect 26016 18164 26022 18176
rect 26237 18173 26249 18176
rect 26283 18173 26295 18207
rect 26237 18167 26295 18173
rect 26418 18164 26424 18216
rect 26476 18164 26482 18216
rect 26973 18207 27031 18213
rect 26973 18173 26985 18207
rect 27019 18204 27031 18207
rect 27522 18204 27528 18216
rect 27019 18176 27528 18204
rect 27019 18173 27031 18176
rect 26973 18167 27031 18173
rect 27522 18164 27528 18176
rect 27580 18164 27586 18216
rect 28905 18207 28963 18213
rect 28905 18173 28917 18207
rect 28951 18204 28963 18207
rect 29454 18204 29460 18216
rect 28951 18176 29460 18204
rect 28951 18173 28963 18176
rect 28905 18167 28963 18173
rect 29454 18164 29460 18176
rect 29512 18164 29518 18216
rect 30852 18213 30880 18244
rect 29917 18207 29975 18213
rect 29917 18173 29929 18207
rect 29963 18204 29975 18207
rect 30837 18207 30895 18213
rect 29963 18176 30788 18204
rect 29963 18173 29975 18176
rect 29917 18167 29975 18173
rect 25976 18136 26004 18164
rect 30760 18148 30788 18176
rect 30837 18173 30849 18207
rect 30883 18204 30895 18207
rect 31389 18207 31447 18213
rect 31389 18204 31401 18207
rect 30883 18176 31401 18204
rect 30883 18173 30895 18176
rect 30837 18167 30895 18173
rect 31389 18173 31401 18176
rect 31435 18173 31447 18207
rect 31389 18167 31447 18173
rect 24412 18108 26004 18136
rect 30193 18139 30251 18145
rect 30193 18105 30205 18139
rect 30239 18136 30251 18139
rect 30374 18136 30380 18148
rect 30239 18108 30380 18136
rect 30239 18105 30251 18108
rect 30193 18099 30251 18105
rect 30374 18096 30380 18108
rect 30432 18096 30438 18148
rect 30742 18096 30748 18148
rect 30800 18136 30806 18148
rect 31757 18139 31815 18145
rect 31757 18136 31769 18139
rect 30800 18108 31769 18136
rect 30800 18096 30806 18108
rect 31757 18105 31769 18108
rect 31803 18105 31815 18139
rect 31757 18099 31815 18105
rect 25774 18068 25780 18080
rect 23768 18040 25780 18068
rect 23201 18031 23259 18037
rect 25774 18028 25780 18040
rect 25832 18028 25838 18080
rect 28074 18028 28080 18080
rect 28132 18028 28138 18080
rect 2760 17978 32200 18000
rect 2760 17926 6946 17978
rect 6998 17926 7010 17978
rect 7062 17926 7074 17978
rect 7126 17926 7138 17978
rect 7190 17926 7202 17978
rect 7254 17926 14306 17978
rect 14358 17926 14370 17978
rect 14422 17926 14434 17978
rect 14486 17926 14498 17978
rect 14550 17926 14562 17978
rect 14614 17926 21666 17978
rect 21718 17926 21730 17978
rect 21782 17926 21794 17978
rect 21846 17926 21858 17978
rect 21910 17926 21922 17978
rect 21974 17926 29026 17978
rect 29078 17926 29090 17978
rect 29142 17926 29154 17978
rect 29206 17926 29218 17978
rect 29270 17926 29282 17978
rect 29334 17926 32200 17978
rect 2760 17904 32200 17926
rect 7282 17864 7288 17876
rect 6104 17836 7288 17864
rect 6104 17737 6132 17836
rect 7282 17824 7288 17836
rect 7340 17864 7346 17876
rect 7340 17836 8064 17864
rect 7340 17824 7346 17836
rect 7926 17796 7932 17808
rect 7590 17768 7932 17796
rect 7926 17756 7932 17768
rect 7984 17756 7990 17808
rect 6089 17731 6147 17737
rect 6089 17697 6101 17731
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 7374 17688 7380 17740
rect 7432 17688 7438 17740
rect 8036 17737 8064 17836
rect 9766 17824 9772 17876
rect 9824 17864 9830 17876
rect 10229 17867 10287 17873
rect 10229 17864 10241 17867
rect 9824 17836 10241 17864
rect 9824 17824 9830 17836
rect 10229 17833 10241 17836
rect 10275 17864 10287 17867
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 10275 17836 10609 17864
rect 10275 17833 10287 17836
rect 10229 17827 10287 17833
rect 10597 17833 10609 17836
rect 10643 17833 10655 17867
rect 10597 17827 10655 17833
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17833 11391 17867
rect 11333 17827 11391 17833
rect 8846 17756 8852 17808
rect 8904 17756 8910 17808
rect 10134 17756 10140 17808
rect 10192 17756 10198 17808
rect 10346 17799 10404 17805
rect 10346 17765 10358 17799
rect 10392 17796 10404 17799
rect 10502 17796 10508 17808
rect 10392 17768 10508 17796
rect 10392 17765 10404 17768
rect 10346 17759 10404 17765
rect 10502 17756 10508 17768
rect 10560 17756 10566 17808
rect 11348 17796 11376 17827
rect 11882 17824 11888 17876
rect 11940 17824 11946 17876
rect 12437 17867 12495 17873
rect 12437 17833 12449 17867
rect 12483 17864 12495 17867
rect 12618 17864 12624 17876
rect 12483 17836 12624 17864
rect 12483 17833 12495 17836
rect 12437 17827 12495 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 12710 17824 12716 17876
rect 12768 17864 12774 17876
rect 13373 17867 13431 17873
rect 13373 17864 13385 17867
rect 12768 17836 13385 17864
rect 12768 17824 12774 17836
rect 13373 17833 13385 17836
rect 13419 17833 13431 17867
rect 13373 17827 13431 17833
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 13771 17836 14504 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 10612 17768 11376 17796
rect 8021 17731 8079 17737
rect 8021 17697 8033 17731
rect 8067 17697 8079 17731
rect 8021 17691 8079 17697
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 9861 17731 9919 17737
rect 9861 17728 9873 17731
rect 9732 17700 9873 17728
rect 9732 17688 9738 17700
rect 9861 17697 9873 17700
rect 9907 17697 9919 17731
rect 10612 17728 10640 17768
rect 11900 17737 11928 17824
rect 13170 17796 13176 17808
rect 12820 17768 13176 17796
rect 9861 17691 9919 17697
rect 10152 17700 10640 17728
rect 11885 17731 11943 17737
rect 6365 17663 6423 17669
rect 6365 17629 6377 17663
rect 6411 17660 6423 17663
rect 7392 17660 7420 17688
rect 10152 17672 10180 17700
rect 11885 17697 11897 17731
rect 11931 17697 11943 17731
rect 11885 17691 11943 17697
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 12820 17737 12848 17768
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 13262 17756 13268 17808
rect 13320 17796 13326 17808
rect 14001 17799 14059 17805
rect 14001 17796 14013 17799
rect 13320 17768 14013 17796
rect 13320 17756 13326 17768
rect 14001 17765 14013 17768
rect 14047 17765 14059 17799
rect 14476 17796 14504 17836
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 16298 17864 16304 17876
rect 14884 17836 16304 17864
rect 14884 17824 14890 17836
rect 16298 17824 16304 17836
rect 16356 17864 16362 17876
rect 16853 17867 16911 17873
rect 16853 17864 16865 17867
rect 16356 17836 16865 17864
rect 16356 17824 16362 17836
rect 16853 17833 16865 17836
rect 16899 17833 16911 17867
rect 16853 17827 16911 17833
rect 22373 17867 22431 17873
rect 22373 17833 22385 17867
rect 22419 17864 22431 17867
rect 22554 17864 22560 17876
rect 22419 17836 22560 17864
rect 22419 17833 22431 17836
rect 22373 17827 22431 17833
rect 22554 17824 22560 17836
rect 22612 17824 22618 17876
rect 22830 17824 22836 17876
rect 22888 17824 22894 17876
rect 23842 17824 23848 17876
rect 23900 17824 23906 17876
rect 25314 17824 25320 17876
rect 25372 17864 25378 17876
rect 25501 17867 25559 17873
rect 25501 17864 25513 17867
rect 25372 17836 25513 17864
rect 25372 17824 25378 17836
rect 25501 17833 25513 17836
rect 25547 17833 25559 17867
rect 25501 17827 25559 17833
rect 25682 17824 25688 17876
rect 25740 17864 25746 17876
rect 25961 17867 26019 17873
rect 25961 17864 25973 17867
rect 25740 17836 25973 17864
rect 25740 17824 25746 17836
rect 25961 17833 25973 17836
rect 26007 17833 26019 17867
rect 28718 17864 28724 17876
rect 25961 17827 26019 17833
rect 26896 17836 28724 17864
rect 14642 17796 14648 17808
rect 14476 17768 14648 17796
rect 14001 17759 14059 17765
rect 14642 17756 14648 17768
rect 14700 17796 14706 17808
rect 15010 17796 15016 17808
rect 14700 17768 15016 17796
rect 14700 17756 14706 17768
rect 15010 17756 15016 17768
rect 15068 17756 15074 17808
rect 16390 17756 16396 17808
rect 16448 17796 16454 17808
rect 16448 17768 16528 17796
rect 16448 17756 16454 17768
rect 12621 17731 12679 17737
rect 12621 17728 12633 17731
rect 12492 17700 12633 17728
rect 12492 17688 12498 17700
rect 12621 17697 12633 17700
rect 12667 17697 12679 17731
rect 12621 17691 12679 17697
rect 12805 17731 12863 17737
rect 12805 17697 12817 17731
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 12897 17731 12955 17737
rect 12897 17697 12909 17731
rect 12943 17728 12955 17731
rect 13538 17728 13544 17740
rect 12943 17700 13544 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 13538 17688 13544 17700
rect 13596 17688 13602 17740
rect 13817 17731 13875 17737
rect 13817 17697 13829 17731
rect 13863 17728 13875 17731
rect 14277 17731 14335 17737
rect 13863 17700 14044 17728
rect 13863 17697 13875 17700
rect 13817 17691 13875 17697
rect 14016 17672 14044 17700
rect 14277 17697 14289 17731
rect 14323 17728 14335 17731
rect 14553 17731 14611 17737
rect 14323 17700 14504 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 6411 17632 7420 17660
rect 6411 17629 6423 17632
rect 6365 17623 6423 17629
rect 8294 17620 8300 17672
rect 8352 17620 8358 17672
rect 10134 17620 10140 17672
rect 10192 17620 10198 17672
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 11609 17663 11667 17669
rect 11609 17629 11621 17663
rect 11655 17660 11667 17663
rect 11974 17660 11980 17672
rect 11655 17632 11980 17660
rect 11655 17629 11667 17632
rect 11609 17623 11667 17629
rect 7834 17552 7840 17604
rect 7892 17552 7898 17604
rect 9769 17595 9827 17601
rect 9769 17561 9781 17595
rect 9815 17592 9827 17595
rect 11164 17592 11192 17623
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17660 12771 17663
rect 12759 17632 13492 17660
rect 12759 17629 12771 17632
rect 12713 17623 12771 17629
rect 13464 17604 13492 17632
rect 13998 17620 14004 17672
rect 14056 17620 14062 17672
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14369 17663 14427 17669
rect 14369 17660 14381 17663
rect 14240 17632 14381 17660
rect 14240 17620 14246 17632
rect 14369 17629 14381 17632
rect 14415 17629 14427 17663
rect 14476 17660 14504 17700
rect 14553 17697 14565 17731
rect 14599 17728 14611 17731
rect 14734 17728 14740 17740
rect 14599 17700 14740 17728
rect 14599 17697 14611 17700
rect 14553 17691 14611 17697
rect 14734 17688 14740 17700
rect 14792 17688 14798 17740
rect 15746 17688 15752 17740
rect 15804 17688 15810 17740
rect 15841 17731 15899 17737
rect 15841 17697 15853 17731
rect 15887 17697 15899 17731
rect 15841 17691 15899 17697
rect 15105 17663 15163 17669
rect 14476 17632 15056 17660
rect 14369 17623 14427 17629
rect 12066 17592 12072 17604
rect 9815 17564 11192 17592
rect 11256 17564 12072 17592
rect 9815 17561 9827 17564
rect 9769 17555 9827 17561
rect 10505 17527 10563 17533
rect 10505 17493 10517 17527
rect 10551 17524 10563 17527
rect 11256 17524 11284 17564
rect 12066 17552 12072 17564
rect 12124 17592 12130 17604
rect 12124 17564 13400 17592
rect 12124 17552 12130 17564
rect 10551 17496 11284 17524
rect 10551 17493 10563 17496
rect 10505 17487 10563 17493
rect 11514 17484 11520 17536
rect 11572 17524 11578 17536
rect 11793 17527 11851 17533
rect 11793 17524 11805 17527
rect 11572 17496 11805 17524
rect 11572 17484 11578 17496
rect 11793 17493 11805 17496
rect 11839 17524 11851 17527
rect 12342 17524 12348 17536
rect 11839 17496 12348 17524
rect 11839 17493 11851 17496
rect 11793 17487 11851 17493
rect 12342 17484 12348 17496
rect 12400 17484 12406 17536
rect 13372 17533 13400 17564
rect 13446 17552 13452 17604
rect 13504 17592 13510 17604
rect 15028 17592 15056 17632
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15289 17663 15347 17669
rect 15289 17660 15301 17663
rect 15151 17632 15301 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 15289 17629 15301 17632
rect 15335 17629 15347 17663
rect 15289 17623 15347 17629
rect 15381 17663 15439 17669
rect 15381 17629 15393 17663
rect 15427 17660 15439 17663
rect 15654 17660 15660 17672
rect 15427 17632 15660 17660
rect 15427 17629 15439 17632
rect 15381 17623 15439 17629
rect 15654 17620 15660 17632
rect 15712 17620 15718 17672
rect 15470 17592 15476 17604
rect 13504 17564 14412 17592
rect 15028 17564 15476 17592
rect 13504 17552 13510 17564
rect 14384 17536 14412 17564
rect 15470 17552 15476 17564
rect 15528 17552 15534 17604
rect 13357 17527 13415 17533
rect 13357 17493 13369 17527
rect 13403 17493 13415 17527
rect 13357 17487 13415 17493
rect 13538 17484 13544 17536
rect 13596 17484 13602 17536
rect 13998 17484 14004 17536
rect 14056 17484 14062 17536
rect 14090 17484 14096 17536
rect 14148 17524 14154 17536
rect 14185 17527 14243 17533
rect 14185 17524 14197 17527
rect 14148 17496 14197 17524
rect 14148 17484 14154 17496
rect 14185 17493 14197 17496
rect 14231 17493 14243 17527
rect 14185 17487 14243 17493
rect 14366 17484 14372 17536
rect 14424 17484 14430 17536
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 15856 17524 15884 17691
rect 16114 17688 16120 17740
rect 16172 17728 16178 17740
rect 16301 17731 16359 17737
rect 16301 17728 16313 17731
rect 16172 17700 16313 17728
rect 16172 17688 16178 17700
rect 16301 17697 16313 17700
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17629 16451 17663
rect 16500 17660 16528 17768
rect 16666 17756 16672 17808
rect 16724 17796 16730 17808
rect 16761 17799 16819 17805
rect 16761 17796 16773 17799
rect 16724 17768 16773 17796
rect 16724 17756 16730 17768
rect 16761 17765 16773 17768
rect 16807 17796 16819 17799
rect 17925 17799 17983 17805
rect 17925 17796 17937 17799
rect 16807 17768 17937 17796
rect 16807 17765 16819 17768
rect 16761 17759 16819 17765
rect 17925 17765 17937 17768
rect 17971 17765 17983 17799
rect 17925 17759 17983 17765
rect 18046 17756 18052 17808
rect 18104 17796 18110 17808
rect 18141 17799 18199 17805
rect 18141 17796 18153 17799
rect 18104 17768 18153 17796
rect 18104 17756 18110 17768
rect 18141 17765 18153 17768
rect 18187 17765 18199 17799
rect 18141 17759 18199 17765
rect 19058 17756 19064 17808
rect 19116 17756 19122 17808
rect 21729 17799 21787 17805
rect 21729 17765 21741 17799
rect 21775 17796 21787 17799
rect 22002 17796 22008 17808
rect 21775 17768 22008 17796
rect 21775 17765 21787 17768
rect 21729 17759 21787 17765
rect 22002 17756 22008 17768
rect 22060 17756 22066 17808
rect 22741 17799 22799 17805
rect 22741 17765 22753 17799
rect 22787 17796 22799 17799
rect 23860 17796 23888 17824
rect 22787 17768 23888 17796
rect 24029 17799 24087 17805
rect 22787 17765 22799 17768
rect 22741 17759 22799 17765
rect 24029 17765 24041 17799
rect 24075 17796 24087 17799
rect 24302 17796 24308 17808
rect 24075 17768 24308 17796
rect 24075 17765 24087 17768
rect 24029 17759 24087 17765
rect 24302 17756 24308 17768
rect 24360 17756 24366 17808
rect 25038 17756 25044 17808
rect 25096 17756 25102 17808
rect 25869 17799 25927 17805
rect 25869 17796 25881 17799
rect 25424 17768 25881 17796
rect 19062 17753 19120 17756
rect 16942 17688 16948 17740
rect 17000 17688 17006 17740
rect 17586 17688 17592 17740
rect 17644 17688 17650 17740
rect 17880 17700 19012 17728
rect 19062 17719 19074 17753
rect 19108 17719 19120 17753
rect 19062 17713 19120 17719
rect 17126 17660 17132 17672
rect 16500 17632 17132 17660
rect 16393 17623 16451 17629
rect 16408 17592 16436 17623
rect 17126 17620 17132 17632
rect 17184 17620 17190 17672
rect 16482 17592 16488 17604
rect 16408 17564 16488 17592
rect 16482 17552 16488 17564
rect 16540 17552 16546 17604
rect 16850 17552 16856 17604
rect 16908 17592 16914 17604
rect 17218 17592 17224 17604
rect 16908 17564 17224 17592
rect 16908 17552 16914 17564
rect 17218 17552 17224 17564
rect 17276 17552 17282 17604
rect 17678 17552 17684 17604
rect 17736 17592 17742 17604
rect 17880 17592 17908 17700
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 18877 17663 18935 17669
rect 18877 17660 18889 17663
rect 18012 17632 18889 17660
rect 18012 17620 18018 17632
rect 18877 17629 18889 17632
rect 18923 17629 18935 17663
rect 18984 17660 19012 17700
rect 19426 17688 19432 17740
rect 19484 17688 19490 17740
rect 20622 17688 20628 17740
rect 20680 17688 20686 17740
rect 19153 17663 19211 17669
rect 19153 17660 19165 17663
rect 18984 17632 19165 17660
rect 18877 17623 18935 17629
rect 19153 17629 19165 17632
rect 19199 17629 19211 17663
rect 19153 17623 19211 17629
rect 19337 17663 19395 17669
rect 19337 17629 19349 17663
rect 19383 17660 19395 17663
rect 19444 17660 19472 17688
rect 25424 17672 25452 17768
rect 25869 17765 25881 17768
rect 25915 17796 25927 17799
rect 26896 17796 26924 17836
rect 28718 17824 28724 17836
rect 28776 17824 28782 17876
rect 28810 17824 28816 17876
rect 28868 17864 28874 17876
rect 30009 17867 30067 17873
rect 30009 17864 30021 17867
rect 28868 17836 30021 17864
rect 28868 17824 28874 17836
rect 30009 17833 30021 17836
rect 30055 17833 30067 17867
rect 30009 17827 30067 17833
rect 27890 17796 27896 17808
rect 25915 17768 26924 17796
rect 27738 17768 27896 17796
rect 25915 17765 25927 17768
rect 25869 17759 25927 17765
rect 27890 17756 27896 17768
rect 27948 17756 27954 17808
rect 28074 17756 28080 17808
rect 28132 17796 28138 17808
rect 28169 17799 28227 17805
rect 28169 17796 28181 17799
rect 28132 17768 28181 17796
rect 28132 17756 28138 17768
rect 28169 17765 28181 17768
rect 28215 17765 28227 17799
rect 28169 17759 28227 17765
rect 28902 17756 28908 17808
rect 28960 17796 28966 17808
rect 29181 17799 29239 17805
rect 29181 17796 29193 17799
rect 28960 17768 29193 17796
rect 28960 17756 28966 17768
rect 29181 17765 29193 17768
rect 29227 17796 29239 17799
rect 29227 17768 29868 17796
rect 29227 17765 29239 17768
rect 29181 17759 29239 17765
rect 25682 17688 25688 17740
rect 25740 17728 25746 17740
rect 26421 17731 26479 17737
rect 26421 17728 26433 17731
rect 25740 17700 26433 17728
rect 25740 17688 25746 17700
rect 26421 17697 26433 17700
rect 26467 17728 26479 17731
rect 26878 17728 26884 17740
rect 26467 17700 26884 17728
rect 26467 17697 26479 17700
rect 26421 17691 26479 17697
rect 26878 17688 26884 17700
rect 26936 17688 26942 17740
rect 19383 17632 19472 17660
rect 19521 17663 19579 17669
rect 19383 17629 19395 17632
rect 19337 17623 19395 17629
rect 19521 17629 19533 17663
rect 19567 17660 19579 17663
rect 19610 17660 19616 17672
rect 19567 17632 19616 17660
rect 19567 17629 19579 17632
rect 19521 17623 19579 17629
rect 19610 17620 19616 17632
rect 19668 17660 19674 17672
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 19668 17632 20269 17660
rect 19668 17620 19674 17632
rect 20257 17629 20269 17632
rect 20303 17660 20315 17663
rect 21266 17660 21272 17672
rect 20303 17632 21272 17660
rect 20303 17629 20315 17632
rect 20257 17623 20315 17629
rect 21266 17620 21272 17632
rect 21324 17620 21330 17672
rect 22005 17663 22063 17669
rect 22005 17629 22017 17663
rect 22051 17660 22063 17663
rect 22094 17660 22100 17672
rect 22051 17632 22100 17660
rect 22051 17629 22063 17632
rect 22005 17623 22063 17629
rect 22094 17620 22100 17632
rect 22152 17620 22158 17672
rect 23017 17663 23075 17669
rect 23017 17629 23029 17663
rect 23063 17660 23075 17663
rect 23566 17660 23572 17672
rect 23063 17632 23572 17660
rect 23063 17629 23075 17632
rect 23017 17623 23075 17629
rect 23566 17620 23572 17632
rect 23624 17620 23630 17672
rect 23750 17620 23756 17672
rect 23808 17620 23814 17672
rect 25406 17620 25412 17672
rect 25464 17620 25470 17672
rect 25777 17663 25835 17669
rect 25777 17629 25789 17663
rect 25823 17660 25835 17663
rect 26786 17660 26792 17672
rect 25823 17632 26792 17660
rect 25823 17629 25835 17632
rect 25777 17623 25835 17629
rect 26786 17620 26792 17632
rect 26844 17620 26850 17672
rect 28445 17663 28503 17669
rect 28445 17629 28457 17663
rect 28491 17660 28503 17663
rect 28994 17660 29000 17672
rect 28491 17632 29000 17660
rect 28491 17629 28503 17632
rect 28445 17623 28503 17629
rect 28994 17620 29000 17632
rect 29052 17660 29058 17672
rect 29362 17660 29368 17672
rect 29052 17632 29368 17660
rect 29052 17620 29058 17632
rect 29362 17620 29368 17632
rect 29420 17620 29426 17672
rect 29840 17660 29868 17768
rect 29914 17688 29920 17740
rect 29972 17688 29978 17740
rect 30653 17731 30711 17737
rect 30653 17697 30665 17731
rect 30699 17728 30711 17731
rect 30834 17728 30840 17740
rect 30699 17700 30840 17728
rect 30699 17697 30711 17700
rect 30653 17691 30711 17697
rect 30834 17688 30840 17700
rect 30892 17688 30898 17740
rect 30101 17663 30159 17669
rect 30101 17660 30113 17663
rect 29840 17632 30113 17660
rect 30101 17629 30113 17632
rect 30147 17629 30159 17663
rect 30101 17623 30159 17629
rect 31665 17663 31723 17669
rect 31665 17629 31677 17663
rect 31711 17660 31723 17663
rect 33134 17660 33140 17672
rect 31711 17632 33140 17660
rect 31711 17629 31723 17632
rect 31665 17623 31723 17629
rect 33134 17620 33140 17632
rect 33192 17620 33198 17672
rect 17736 17564 17908 17592
rect 17736 17552 17742 17564
rect 18138 17552 18144 17604
rect 18196 17592 18202 17604
rect 19245 17595 19303 17601
rect 19245 17592 19257 17595
rect 18196 17564 19257 17592
rect 18196 17552 18202 17564
rect 19245 17561 19257 17564
rect 19291 17561 19303 17595
rect 19245 17555 19303 17561
rect 17310 17524 17316 17536
rect 14516 17496 17316 17524
rect 14516 17484 14522 17496
rect 17310 17484 17316 17496
rect 17368 17524 17374 17536
rect 17497 17527 17555 17533
rect 17497 17524 17509 17527
rect 17368 17496 17509 17524
rect 17368 17484 17374 17496
rect 17497 17493 17509 17496
rect 17543 17493 17555 17527
rect 17497 17487 17555 17493
rect 17773 17527 17831 17533
rect 17773 17493 17785 17527
rect 17819 17524 17831 17527
rect 17862 17524 17868 17536
rect 17819 17496 17868 17524
rect 17819 17493 17831 17496
rect 17773 17487 17831 17493
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 17954 17484 17960 17536
rect 18012 17484 18018 17536
rect 18230 17484 18236 17536
rect 18288 17524 18294 17536
rect 18325 17527 18383 17533
rect 18325 17524 18337 17527
rect 18288 17496 18337 17524
rect 18288 17484 18294 17496
rect 18325 17493 18337 17496
rect 18371 17493 18383 17527
rect 18325 17487 18383 17493
rect 20070 17484 20076 17536
rect 20128 17484 20134 17536
rect 26326 17484 26332 17536
rect 26384 17484 26390 17536
rect 29546 17484 29552 17536
rect 29604 17484 29610 17536
rect 2760 17434 32200 17456
rect 2760 17382 6286 17434
rect 6338 17382 6350 17434
rect 6402 17382 6414 17434
rect 6466 17382 6478 17434
rect 6530 17382 6542 17434
rect 6594 17382 13646 17434
rect 13698 17382 13710 17434
rect 13762 17382 13774 17434
rect 13826 17382 13838 17434
rect 13890 17382 13902 17434
rect 13954 17382 21006 17434
rect 21058 17382 21070 17434
rect 21122 17382 21134 17434
rect 21186 17382 21198 17434
rect 21250 17382 21262 17434
rect 21314 17382 28366 17434
rect 28418 17382 28430 17434
rect 28482 17382 28494 17434
rect 28546 17382 28558 17434
rect 28610 17382 28622 17434
rect 28674 17382 32200 17434
rect 2760 17360 32200 17382
rect 8294 17280 8300 17332
rect 8352 17320 8358 17332
rect 9309 17323 9367 17329
rect 9309 17320 9321 17323
rect 8352 17292 9321 17320
rect 8352 17280 8358 17292
rect 9309 17289 9321 17292
rect 9355 17289 9367 17323
rect 9309 17283 9367 17289
rect 10594 17280 10600 17332
rect 10652 17280 10658 17332
rect 11698 17280 11704 17332
rect 11756 17320 11762 17332
rect 11885 17323 11943 17329
rect 11885 17320 11897 17323
rect 11756 17292 11897 17320
rect 11756 17280 11762 17292
rect 11885 17289 11897 17292
rect 11931 17289 11943 17323
rect 11885 17283 11943 17289
rect 12986 17280 12992 17332
rect 13044 17320 13050 17332
rect 13081 17323 13139 17329
rect 13081 17320 13093 17323
rect 13044 17292 13093 17320
rect 13044 17280 13050 17292
rect 13081 17289 13093 17292
rect 13127 17289 13139 17323
rect 13081 17283 13139 17289
rect 13262 17280 13268 17332
rect 13320 17280 13326 17332
rect 13538 17280 13544 17332
rect 13596 17280 13602 17332
rect 13909 17323 13967 17329
rect 13909 17289 13921 17323
rect 13955 17289 13967 17323
rect 13909 17283 13967 17289
rect 9217 17255 9275 17261
rect 9217 17221 9229 17255
rect 9263 17252 9275 17255
rect 10612 17252 10640 17280
rect 9263 17224 10640 17252
rect 9263 17221 9275 17224
rect 9217 17215 9275 17221
rect 7745 17187 7803 17193
rect 7745 17153 7757 17187
rect 7791 17184 7803 17187
rect 8110 17184 8116 17196
rect 7791 17156 8116 17184
rect 7791 17153 7803 17156
rect 7745 17147 7803 17153
rect 8110 17144 8116 17156
rect 8168 17144 8174 17196
rect 9766 17144 9772 17196
rect 9824 17144 9830 17196
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17184 10011 17187
rect 10042 17184 10048 17196
rect 9999 17156 10048 17184
rect 9999 17153 10011 17156
rect 9953 17147 10011 17153
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 12158 17144 12164 17196
rect 12216 17144 12222 17196
rect 7282 17076 7288 17128
rect 7340 17116 7346 17128
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 7340 17088 7481 17116
rect 7340 17076 7346 17088
rect 7469 17085 7481 17088
rect 7515 17085 7527 17119
rect 7469 17079 7527 17085
rect 9674 17076 9680 17128
rect 9732 17076 9738 17128
rect 10962 17076 10968 17128
rect 11020 17076 11026 17128
rect 11977 17119 12035 17125
rect 11977 17085 11989 17119
rect 12023 17116 12035 17119
rect 12176 17116 12204 17144
rect 12023 17088 12204 17116
rect 12023 17085 12035 17088
rect 11977 17079 12035 17085
rect 12250 17076 12256 17128
rect 12308 17076 12314 17128
rect 12342 17076 12348 17128
rect 12400 17116 12406 17128
rect 12897 17119 12955 17125
rect 12400 17088 12445 17116
rect 12400 17076 12406 17088
rect 12897 17085 12909 17119
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 8478 17008 8484 17060
rect 8536 17008 8542 17060
rect 9692 17048 9720 17076
rect 9950 17048 9956 17060
rect 9692 17020 9956 17048
rect 9950 17008 9956 17020
rect 10008 17048 10014 17060
rect 11333 17051 11391 17057
rect 11333 17048 11345 17051
rect 10008 17020 11345 17048
rect 10008 17008 10014 17020
rect 11333 17017 11345 17020
rect 11379 17017 11391 17051
rect 11333 17011 11391 17017
rect 11425 17051 11483 17057
rect 11425 17017 11437 17051
rect 11471 17048 11483 17051
rect 11514 17048 11520 17060
rect 11471 17020 11520 17048
rect 11471 17017 11483 17020
rect 11425 17011 11483 17017
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 12161 17051 12219 17057
rect 12161 17048 12173 17051
rect 11992 17020 12173 17048
rect 11992 16992 12020 17020
rect 12161 17017 12173 17020
rect 12207 17048 12219 17051
rect 12912 17048 12940 17079
rect 12207 17020 12940 17048
rect 13280 17048 13308 17280
rect 13556 17184 13584 17280
rect 13464 17156 13584 17184
rect 13924 17184 13952 17283
rect 13998 17280 14004 17332
rect 14056 17280 14062 17332
rect 14185 17323 14243 17329
rect 14185 17289 14197 17323
rect 14231 17320 14243 17323
rect 14366 17320 14372 17332
rect 14231 17292 14372 17320
rect 14231 17289 14243 17292
rect 14185 17283 14243 17289
rect 14366 17280 14372 17292
rect 14424 17320 14430 17332
rect 16022 17320 16028 17332
rect 14424 17292 16028 17320
rect 14424 17280 14430 17292
rect 16022 17280 16028 17292
rect 16080 17280 16086 17332
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16301 17323 16359 17329
rect 16301 17320 16313 17323
rect 16264 17292 16313 17320
rect 16264 17280 16270 17292
rect 16301 17289 16313 17292
rect 16347 17289 16359 17323
rect 16301 17283 16359 17289
rect 16390 17280 16396 17332
rect 16448 17280 16454 17332
rect 17586 17280 17592 17332
rect 17644 17320 17650 17332
rect 18877 17323 18935 17329
rect 18877 17320 18889 17323
rect 17644 17292 18889 17320
rect 17644 17280 17650 17292
rect 18877 17289 18889 17292
rect 18923 17289 18935 17323
rect 18877 17283 18935 17289
rect 20622 17280 20628 17332
rect 20680 17320 20686 17332
rect 20993 17323 21051 17329
rect 20993 17320 21005 17323
rect 20680 17292 21005 17320
rect 20680 17280 20686 17292
rect 20993 17289 21005 17292
rect 21039 17289 21051 17323
rect 20993 17283 21051 17289
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 25038 17320 25044 17332
rect 24903 17292 25044 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 25038 17280 25044 17292
rect 25096 17280 25102 17332
rect 28813 17323 28871 17329
rect 28813 17289 28825 17323
rect 28859 17320 28871 17323
rect 28902 17320 28908 17332
rect 28859 17292 28908 17320
rect 28859 17289 28871 17292
rect 28813 17283 28871 17289
rect 28902 17280 28908 17292
rect 28960 17280 28966 17332
rect 29227 17323 29285 17329
rect 29227 17289 29239 17323
rect 29273 17320 29285 17323
rect 29454 17320 29460 17332
rect 29273 17292 29460 17320
rect 29273 17289 29285 17292
rect 29227 17283 29285 17289
rect 29454 17280 29460 17292
rect 29512 17280 29518 17332
rect 29914 17280 29920 17332
rect 29972 17320 29978 17332
rect 31205 17323 31263 17329
rect 31205 17320 31217 17323
rect 29972 17292 31217 17320
rect 29972 17280 29978 17292
rect 31205 17289 31217 17292
rect 31251 17289 31263 17323
rect 31205 17283 31263 17289
rect 14016 17252 14044 17280
rect 14550 17252 14556 17264
rect 14016 17224 14556 17252
rect 14550 17212 14556 17224
rect 14608 17212 14614 17264
rect 16114 17252 16120 17264
rect 14936 17224 16120 17252
rect 14274 17184 14280 17196
rect 13924 17156 14280 17184
rect 13354 17076 13360 17128
rect 13412 17076 13418 17128
rect 13464 17125 13492 17156
rect 14274 17144 14280 17156
rect 14332 17144 14338 17196
rect 14936 17184 14964 17224
rect 16114 17212 16120 17224
rect 16172 17212 16178 17264
rect 16408 17252 16436 17280
rect 16853 17255 16911 17261
rect 16853 17252 16865 17255
rect 16408 17224 16865 17252
rect 16853 17221 16865 17224
rect 16899 17252 16911 17255
rect 17954 17252 17960 17264
rect 16899 17224 17960 17252
rect 16899 17221 16911 17224
rect 16853 17215 16911 17221
rect 17954 17212 17960 17224
rect 18012 17212 18018 17264
rect 18138 17212 18144 17264
rect 18196 17212 18202 17264
rect 14568 17156 14964 17184
rect 13449 17119 13507 17125
rect 13449 17085 13461 17119
rect 13495 17085 13507 17119
rect 13449 17079 13507 17085
rect 13538 17076 13544 17128
rect 13596 17076 13602 17128
rect 13998 17076 14004 17128
rect 14056 17116 14062 17128
rect 14458 17125 14464 17128
rect 14441 17119 14464 17125
rect 14441 17118 14453 17119
rect 14056 17112 14353 17116
rect 14430 17112 14453 17118
rect 14056 17088 14453 17112
rect 14056 17076 14062 17088
rect 14325 17085 14453 17088
rect 14325 17084 14464 17085
rect 14441 17079 14464 17084
rect 14458 17076 14464 17079
rect 14516 17076 14522 17128
rect 14568 17122 14596 17156
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15068 17156 15231 17184
rect 15068 17144 15074 17156
rect 14553 17116 14611 17122
rect 14553 17082 14565 17116
rect 14599 17082 14611 17116
rect 14553 17076 14611 17082
rect 14645 17116 14703 17122
rect 14645 17082 14657 17116
rect 14691 17082 14703 17116
rect 14645 17076 14703 17082
rect 14823 17119 14881 17125
rect 14823 17085 14835 17119
rect 14869 17085 14881 17119
rect 14823 17079 14881 17085
rect 13280 17020 14136 17048
rect 12207 17017 12219 17020
rect 12161 17011 12219 17017
rect 9677 16983 9735 16989
rect 9677 16949 9689 16983
rect 9723 16980 9735 16983
rect 10226 16980 10232 16992
rect 9723 16952 10232 16980
rect 9723 16949 9735 16952
rect 9677 16943 9735 16949
rect 10226 16940 10232 16952
rect 10284 16980 10290 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 10284 16952 10333 16980
rect 10284 16940 10290 16952
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 10321 16943 10379 16949
rect 11974 16940 11980 16992
rect 12032 16940 12038 16992
rect 12618 16940 12624 16992
rect 12676 16940 12682 16992
rect 12802 16940 12808 16992
rect 12860 16940 12866 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 14108 16989 14136 17020
rect 13909 16983 13967 16989
rect 13909 16980 13921 16983
rect 13596 16952 13921 16980
rect 13596 16940 13602 16952
rect 13909 16949 13921 16952
rect 13955 16949 13967 16983
rect 13909 16943 13967 16949
rect 14093 16983 14151 16989
rect 14093 16949 14105 16983
rect 14139 16949 14151 16983
rect 14660 16980 14688 17076
rect 14844 17048 14872 17079
rect 14918 17076 14924 17128
rect 14976 17076 14982 17128
rect 15102 17076 15108 17128
rect 15160 17076 15166 17128
rect 15203 17116 15231 17156
rect 15746 17144 15752 17196
rect 15804 17184 15810 17196
rect 16298 17184 16304 17196
rect 15804 17156 16304 17184
rect 15804 17144 15810 17156
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 17034 17144 17040 17196
rect 17092 17144 17098 17196
rect 17126 17144 17132 17196
rect 17184 17184 17190 17196
rect 18046 17184 18052 17196
rect 17184 17156 18052 17184
rect 17184 17144 17190 17156
rect 18046 17144 18052 17156
rect 18104 17144 18110 17196
rect 16025 17119 16083 17125
rect 16025 17116 16037 17119
rect 15203 17088 16037 17116
rect 16025 17085 16037 17088
rect 16071 17085 16083 17119
rect 16025 17079 16083 17085
rect 16209 17119 16267 17125
rect 16209 17085 16221 17119
rect 16255 17116 16267 17119
rect 16574 17116 16580 17128
rect 16255 17088 16580 17116
rect 16255 17085 16267 17088
rect 16209 17079 16267 17085
rect 15120 17048 15148 17076
rect 16224 17048 16252 17079
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 16758 17076 16764 17128
rect 16816 17076 16822 17128
rect 17052 17116 17080 17144
rect 17221 17119 17279 17125
rect 17221 17116 17233 17119
rect 17052 17088 17233 17116
rect 17221 17085 17233 17088
rect 17267 17085 17279 17119
rect 17221 17079 17279 17085
rect 17310 17076 17316 17128
rect 17368 17116 17374 17128
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 17368 17088 17509 17116
rect 17368 17076 17374 17088
rect 17497 17085 17509 17088
rect 17543 17085 17555 17119
rect 17497 17079 17555 17085
rect 17586 17076 17592 17128
rect 17644 17076 17650 17128
rect 18156 17116 18184 17212
rect 19334 17144 19340 17196
rect 19392 17184 19398 17196
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 19392 17156 20637 17184
rect 19392 17144 19398 17156
rect 20625 17153 20637 17156
rect 20671 17184 20683 17187
rect 22094 17184 22100 17196
rect 20671 17156 22100 17184
rect 20671 17153 20683 17156
rect 20625 17147 20683 17153
rect 22094 17144 22100 17156
rect 22152 17184 22158 17196
rect 23017 17187 23075 17193
rect 23017 17184 23029 17187
rect 22152 17156 23029 17184
rect 22152 17144 22158 17156
rect 23017 17153 23029 17156
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 28169 17187 28227 17193
rect 28169 17153 28181 17187
rect 28215 17184 28227 17187
rect 28994 17184 29000 17196
rect 28215 17156 29000 17184
rect 28215 17153 28227 17156
rect 28169 17147 28227 17153
rect 28994 17144 29000 17156
rect 29052 17184 29058 17196
rect 31021 17187 31079 17193
rect 31021 17184 31033 17187
rect 29052 17156 31033 17184
rect 29052 17144 29058 17156
rect 31021 17153 31033 17156
rect 31067 17153 31079 17187
rect 31021 17147 31079 17153
rect 17972 17088 18184 17116
rect 14844 17020 15148 17048
rect 15304 17020 16252 17048
rect 15304 16992 15332 17020
rect 17034 17008 17040 17060
rect 17092 17008 17098 17060
rect 17129 17051 17187 17057
rect 17129 17017 17141 17051
rect 17175 17048 17187 17051
rect 17972 17048 18000 17088
rect 18506 17076 18512 17128
rect 18564 17116 18570 17128
rect 18693 17119 18751 17125
rect 18693 17116 18705 17119
rect 18564 17088 18705 17116
rect 18564 17076 18570 17088
rect 18693 17085 18705 17088
rect 18739 17085 18751 17119
rect 18693 17079 18751 17085
rect 19242 17076 19248 17128
rect 19300 17076 19306 17128
rect 21085 17119 21143 17125
rect 21085 17085 21097 17119
rect 21131 17116 21143 17119
rect 21450 17116 21456 17128
rect 21131 17088 21456 17116
rect 21131 17085 21143 17088
rect 21085 17079 21143 17085
rect 21450 17076 21456 17088
rect 21508 17076 21514 17128
rect 23106 17076 23112 17128
rect 23164 17076 23170 17128
rect 23293 17119 23351 17125
rect 23293 17085 23305 17119
rect 23339 17085 23351 17119
rect 23293 17079 23351 17085
rect 17175 17020 18000 17048
rect 17175 17017 17187 17020
rect 17129 17011 17187 17017
rect 18046 17008 18052 17060
rect 18104 17008 18110 17060
rect 20346 17008 20352 17060
rect 20404 17008 20410 17060
rect 22741 17051 22799 17057
rect 22310 17020 22692 17048
rect 14826 16980 14832 16992
rect 14660 16952 14832 16980
rect 14093 16943 14151 16949
rect 14826 16940 14832 16952
rect 14884 16940 14890 16992
rect 15010 16940 15016 16992
rect 15068 16980 15074 16992
rect 15105 16983 15163 16989
rect 15105 16980 15117 16983
rect 15068 16952 15117 16980
rect 15068 16940 15074 16952
rect 15105 16949 15117 16952
rect 15151 16949 15163 16983
rect 15105 16943 15163 16949
rect 15286 16940 15292 16992
rect 15344 16940 15350 16992
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15841 16983 15899 16989
rect 15841 16980 15853 16983
rect 15436 16952 15853 16980
rect 15436 16940 15442 16952
rect 15841 16949 15853 16952
rect 15887 16949 15899 16983
rect 15841 16943 15899 16949
rect 15930 16940 15936 16992
rect 15988 16980 15994 16992
rect 16577 16983 16635 16989
rect 16577 16980 16589 16983
rect 15988 16952 16589 16980
rect 15988 16940 15994 16952
rect 16577 16949 16589 16952
rect 16623 16980 16635 16983
rect 16666 16980 16672 16992
rect 16623 16952 16672 16980
rect 16623 16949 16635 16952
rect 16577 16943 16635 16949
rect 16666 16940 16672 16952
rect 16724 16980 16730 16992
rect 17310 16980 17316 16992
rect 16724 16952 17316 16980
rect 16724 16940 16730 16952
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17405 16983 17463 16989
rect 17405 16949 17417 16983
rect 17451 16980 17463 16983
rect 17862 16980 17868 16992
rect 17451 16952 17868 16980
rect 17451 16949 17463 16952
rect 17405 16943 17463 16949
rect 17862 16940 17868 16952
rect 17920 16940 17926 16992
rect 17954 16940 17960 16992
rect 18012 16980 18018 16992
rect 18141 16983 18199 16989
rect 18141 16980 18153 16983
rect 18012 16952 18153 16980
rect 18012 16940 18018 16952
rect 18141 16949 18153 16952
rect 18187 16949 18199 16983
rect 18141 16943 18199 16949
rect 21266 16940 21272 16992
rect 21324 16940 21330 16992
rect 22664 16980 22692 17020
rect 22741 17017 22753 17051
rect 22787 17048 22799 17051
rect 23124 17048 23152 17076
rect 22787 17020 23152 17048
rect 23201 17051 23259 17057
rect 22787 17017 22799 17020
rect 22741 17011 22799 17017
rect 23201 17017 23213 17051
rect 23247 17017 23259 17051
rect 23308 17048 23336 17079
rect 24946 17076 24952 17128
rect 25004 17076 25010 17128
rect 28905 17119 28963 17125
rect 28905 17085 28917 17119
rect 28951 17085 28963 17119
rect 28905 17079 28963 17085
rect 23658 17048 23664 17060
rect 23308 17020 23664 17048
rect 23201 17011 23259 17017
rect 23216 16980 23244 17011
rect 23658 17008 23664 17020
rect 23716 17048 23722 17060
rect 23716 17020 26556 17048
rect 23716 17008 23722 17020
rect 26528 16992 26556 17020
rect 27338 17008 27344 17060
rect 27396 17008 27402 17060
rect 27893 17051 27951 17057
rect 27893 17017 27905 17051
rect 27939 17017 27951 17051
rect 27893 17011 27951 17017
rect 22664 16952 23244 16980
rect 25406 16940 25412 16992
rect 25464 16940 25470 16992
rect 25498 16940 25504 16992
rect 25556 16980 25562 16992
rect 26421 16983 26479 16989
rect 26421 16980 26433 16983
rect 25556 16952 26433 16980
rect 25556 16940 25562 16952
rect 26421 16949 26433 16952
rect 26467 16949 26479 16983
rect 26421 16943 26479 16949
rect 26510 16940 26516 16992
rect 26568 16940 26574 16992
rect 27062 16940 27068 16992
rect 27120 16980 27126 16992
rect 27908 16980 27936 17011
rect 28920 16992 28948 17079
rect 30650 17076 30656 17128
rect 30708 17076 30714 17128
rect 30926 17076 30932 17128
rect 30984 17116 30990 17128
rect 31757 17119 31815 17125
rect 31757 17116 31769 17119
rect 30984 17088 31769 17116
rect 30984 17076 30990 17088
rect 31757 17085 31769 17088
rect 31803 17085 31815 17119
rect 31757 17079 31815 17085
rect 28997 17051 29055 17057
rect 28997 17017 29009 17051
rect 29043 17048 29055 17051
rect 29043 17020 29670 17048
rect 29043 17017 29055 17020
rect 28997 17011 29055 17017
rect 27120 16952 27936 16980
rect 27120 16940 27126 16952
rect 28902 16940 28908 16992
rect 28960 16980 28966 16992
rect 30374 16980 30380 16992
rect 28960 16952 30380 16980
rect 28960 16940 28966 16952
rect 30374 16940 30380 16952
rect 30432 16940 30438 16992
rect 2760 16890 32200 16912
rect 2760 16838 6946 16890
rect 6998 16838 7010 16890
rect 7062 16838 7074 16890
rect 7126 16838 7138 16890
rect 7190 16838 7202 16890
rect 7254 16838 14306 16890
rect 14358 16838 14370 16890
rect 14422 16838 14434 16890
rect 14486 16838 14498 16890
rect 14550 16838 14562 16890
rect 14614 16838 21666 16890
rect 21718 16838 21730 16890
rect 21782 16838 21794 16890
rect 21846 16838 21858 16890
rect 21910 16838 21922 16890
rect 21974 16838 29026 16890
rect 29078 16838 29090 16890
rect 29142 16838 29154 16890
rect 29206 16838 29218 16890
rect 29270 16838 29282 16890
rect 29334 16838 32200 16890
rect 2760 16816 32200 16838
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 7984 16748 8217 16776
rect 7984 16736 7990 16748
rect 8205 16745 8217 16748
rect 8251 16745 8263 16779
rect 8205 16739 8263 16745
rect 8294 16736 8300 16788
rect 8352 16736 8358 16788
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 8573 16779 8631 16785
rect 8573 16776 8585 16779
rect 8536 16748 8585 16776
rect 8536 16736 8542 16748
rect 8573 16745 8585 16748
rect 8619 16745 8631 16779
rect 8573 16739 8631 16745
rect 8846 16736 8852 16788
rect 8904 16736 8910 16788
rect 9122 16736 9128 16788
rect 9180 16736 9186 16788
rect 10962 16736 10968 16788
rect 11020 16776 11026 16788
rect 11793 16779 11851 16785
rect 11793 16776 11805 16779
rect 11020 16748 11805 16776
rect 11020 16736 11026 16748
rect 11793 16745 11805 16748
rect 11839 16776 11851 16779
rect 13078 16776 13084 16788
rect 11839 16748 13084 16776
rect 11839 16745 11851 16748
rect 11793 16739 11851 16745
rect 5902 16600 5908 16652
rect 5960 16600 5966 16652
rect 8312 16649 8340 16736
rect 10428 16680 11744 16708
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16640 8355 16643
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 8343 16612 8493 16640
rect 8343 16609 8355 16612
rect 8297 16603 8355 16609
rect 8481 16609 8493 16612
rect 8527 16640 8539 16643
rect 8757 16643 8815 16649
rect 8757 16640 8769 16643
rect 8527 16612 8769 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 8757 16609 8769 16612
rect 8803 16640 8815 16643
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8803 16612 9045 16640
rect 8803 16609 8815 16612
rect 8757 16603 8815 16609
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 9033 16603 9091 16609
rect 10134 16600 10140 16652
rect 10192 16640 10198 16652
rect 10428 16649 10456 16680
rect 11716 16652 11744 16680
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 10192 16612 10241 16640
rect 10192 16600 10198 16612
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 10413 16643 10471 16649
rect 10413 16609 10425 16643
rect 10459 16609 10471 16643
rect 10413 16603 10471 16609
rect 10962 16600 10968 16652
rect 11020 16600 11026 16652
rect 11333 16643 11391 16649
rect 11333 16609 11345 16643
rect 11379 16640 11391 16643
rect 11606 16640 11612 16652
rect 11379 16612 11612 16640
rect 11379 16609 11391 16612
rect 11333 16603 11391 16609
rect 11606 16600 11612 16612
rect 11664 16600 11670 16652
rect 11698 16600 11704 16652
rect 11756 16600 11762 16652
rect 11808 16640 11836 16739
rect 13078 16736 13084 16748
rect 13136 16736 13142 16788
rect 14090 16736 14096 16788
rect 14148 16736 14154 16788
rect 14826 16736 14832 16788
rect 14884 16776 14890 16788
rect 15013 16779 15071 16785
rect 15013 16776 15025 16779
rect 14884 16748 15025 16776
rect 14884 16736 14890 16748
rect 15013 16745 15025 16748
rect 15059 16745 15071 16779
rect 15013 16739 15071 16745
rect 15562 16736 15568 16788
rect 15620 16776 15626 16788
rect 15841 16779 15899 16785
rect 15841 16776 15853 16779
rect 15620 16748 15853 16776
rect 15620 16736 15626 16748
rect 15841 16745 15853 16748
rect 15887 16745 15899 16779
rect 15841 16739 15899 16745
rect 16025 16779 16083 16785
rect 16025 16745 16037 16779
rect 16071 16776 16083 16779
rect 16071 16748 16160 16776
rect 16071 16745 16083 16748
rect 16025 16739 16083 16745
rect 12820 16680 13492 16708
rect 12820 16652 12848 16680
rect 12069 16643 12127 16649
rect 12069 16640 12081 16643
rect 11808 16612 12081 16640
rect 12069 16609 12081 16612
rect 12115 16609 12127 16643
rect 12069 16603 12127 16609
rect 12621 16643 12679 16649
rect 12621 16609 12633 16643
rect 12667 16640 12679 16643
rect 12802 16640 12808 16652
rect 12667 16612 12808 16640
rect 12667 16609 12679 16612
rect 12621 16603 12679 16609
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13354 16640 13360 16652
rect 13311 16612 13360 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13354 16600 13360 16612
rect 13412 16600 13418 16652
rect 13464 16649 13492 16680
rect 13998 16668 14004 16720
rect 14056 16708 14062 16720
rect 14369 16711 14427 16717
rect 14369 16708 14381 16711
rect 14056 16680 14381 16708
rect 14056 16668 14062 16680
rect 14369 16677 14381 16680
rect 14415 16677 14427 16711
rect 14369 16671 14427 16677
rect 14752 16680 15148 16708
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16609 13507 16643
rect 13449 16603 13507 16609
rect 13541 16643 13599 16649
rect 13541 16609 13553 16643
rect 13587 16609 13599 16643
rect 13541 16603 13599 16609
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 14752 16640 14780 16680
rect 15120 16649 15148 16680
rect 14921 16643 14979 16649
rect 14921 16640 14933 16643
rect 13771 16612 14780 16640
rect 14844 16612 14933 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 10321 16575 10379 16581
rect 10321 16541 10333 16575
rect 10367 16572 10379 16575
rect 11425 16575 11483 16581
rect 10367 16544 10456 16572
rect 10367 16541 10379 16544
rect 10321 16535 10379 16541
rect 10428 16516 10456 16544
rect 11425 16541 11437 16575
rect 11471 16572 11483 16575
rect 11514 16572 11520 16584
rect 11471 16544 11520 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 11514 16532 11520 16544
rect 11572 16532 11578 16584
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 12084 16544 12265 16572
rect 12084 16516 12112 16544
rect 12253 16541 12265 16544
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 12529 16575 12587 16581
rect 12529 16541 12541 16575
rect 12575 16572 12587 16575
rect 13556 16572 13584 16603
rect 14844 16572 14872 16612
rect 14921 16609 14933 16612
rect 14967 16609 14979 16643
rect 14921 16603 14979 16609
rect 15105 16643 15163 16649
rect 15105 16609 15117 16643
rect 15151 16609 15163 16643
rect 15105 16603 15163 16609
rect 15194 16600 15200 16652
rect 15252 16640 15258 16652
rect 15381 16643 15439 16649
rect 15381 16640 15393 16643
rect 15252 16612 15393 16640
rect 15252 16600 15258 16612
rect 15381 16609 15393 16612
rect 15427 16640 15439 16643
rect 15966 16643 16024 16649
rect 15966 16640 15978 16643
rect 15427 16612 15978 16640
rect 15427 16609 15439 16612
rect 15381 16603 15439 16609
rect 15966 16609 15978 16612
rect 16012 16609 16024 16643
rect 15966 16603 16024 16609
rect 12575 16544 13584 16572
rect 14660 16544 14872 16572
rect 15028 16544 15700 16572
rect 12575 16541 12587 16544
rect 12529 16535 12587 16541
rect 6730 16464 6736 16516
rect 6788 16504 6794 16516
rect 6788 16476 10364 16504
rect 6788 16464 6794 16476
rect 5258 16396 5264 16448
rect 5316 16396 5322 16448
rect 10336 16436 10364 16476
rect 10410 16464 10416 16516
rect 10468 16464 10474 16516
rect 12066 16464 12072 16516
rect 12124 16464 12130 16516
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12544 16504 12572 16535
rect 12216 16476 12572 16504
rect 13357 16507 13415 16513
rect 12216 16464 12222 16476
rect 13357 16473 13369 16507
rect 13403 16473 13415 16507
rect 13357 16467 13415 16473
rect 12526 16436 12532 16448
rect 10336 16408 12532 16436
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 13372 16436 13400 16467
rect 12676 16408 13400 16436
rect 14660 16436 14688 16544
rect 14737 16507 14795 16513
rect 14737 16473 14749 16507
rect 14783 16504 14795 16507
rect 15028 16504 15056 16544
rect 14783 16476 15056 16504
rect 15672 16504 15700 16544
rect 15746 16532 15752 16584
rect 15804 16572 15810 16584
rect 16132 16572 16160 16748
rect 16482 16736 16488 16788
rect 16540 16776 16546 16788
rect 17221 16779 17279 16785
rect 17221 16776 17233 16779
rect 16540 16748 17233 16776
rect 16540 16736 16546 16748
rect 17221 16745 17233 16748
rect 17267 16776 17279 16779
rect 18785 16779 18843 16785
rect 18785 16776 18797 16779
rect 17267 16748 18797 16776
rect 17267 16745 17279 16748
rect 17221 16739 17279 16745
rect 18785 16745 18797 16748
rect 18831 16745 18843 16779
rect 18785 16739 18843 16745
rect 20070 16736 20076 16788
rect 20128 16736 20134 16788
rect 21266 16736 21272 16788
rect 21324 16776 21330 16788
rect 21324 16748 22094 16776
rect 21324 16736 21330 16748
rect 17586 16708 17592 16720
rect 16684 16680 17592 16708
rect 16684 16652 16712 16680
rect 17586 16668 17592 16680
rect 17644 16668 17650 16720
rect 17770 16708 17776 16720
rect 17696 16680 17776 16708
rect 16206 16600 16212 16652
rect 16264 16640 16270 16652
rect 16393 16643 16451 16649
rect 16393 16640 16405 16643
rect 16264 16612 16405 16640
rect 16264 16600 16270 16612
rect 16393 16609 16405 16612
rect 16439 16609 16451 16643
rect 16393 16603 16451 16609
rect 16574 16600 16580 16652
rect 16632 16600 16638 16652
rect 16666 16600 16672 16652
rect 16724 16600 16730 16652
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 16776 16612 17417 16640
rect 15804 16544 16160 16572
rect 16485 16575 16543 16581
rect 15804 16532 15810 16544
rect 16485 16541 16497 16575
rect 16531 16541 16543 16575
rect 16592 16572 16620 16600
rect 16776 16572 16804 16612
rect 17405 16609 17417 16612
rect 17451 16609 17463 16643
rect 17405 16603 17463 16609
rect 17497 16643 17555 16649
rect 17497 16609 17509 16643
rect 17543 16640 17555 16643
rect 17696 16640 17724 16680
rect 17770 16668 17776 16680
rect 17828 16708 17834 16720
rect 20088 16708 20116 16736
rect 20257 16711 20315 16717
rect 20257 16708 20269 16711
rect 17828 16680 19472 16708
rect 20088 16680 20269 16708
rect 17828 16668 17834 16680
rect 19444 16652 19472 16680
rect 20257 16677 20269 16680
rect 20303 16677 20315 16711
rect 20257 16671 20315 16677
rect 17543 16612 17724 16640
rect 18693 16643 18751 16649
rect 17543 16609 17555 16612
rect 17497 16603 17555 16609
rect 18693 16609 18705 16643
rect 18739 16640 18751 16643
rect 19337 16643 19395 16649
rect 19337 16640 19349 16643
rect 18739 16612 19349 16640
rect 18739 16609 18751 16612
rect 18693 16603 18751 16609
rect 19337 16609 19349 16612
rect 19383 16609 19395 16643
rect 19337 16603 19395 16609
rect 16592 16544 16804 16572
rect 16485 16535 16543 16541
rect 16500 16504 16528 16535
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17512 16572 17540 16603
rect 19426 16600 19432 16652
rect 19484 16600 19490 16652
rect 19518 16600 19524 16652
rect 19576 16640 19582 16652
rect 20073 16643 20131 16649
rect 20073 16640 20085 16643
rect 19576 16612 20085 16640
rect 19576 16600 19582 16612
rect 20073 16609 20085 16612
rect 20119 16609 20131 16643
rect 22066 16640 22094 16748
rect 22830 16736 22836 16788
rect 22888 16736 22894 16788
rect 26326 16736 26332 16788
rect 26384 16736 26390 16788
rect 27062 16736 27068 16788
rect 27120 16736 27126 16788
rect 27338 16736 27344 16788
rect 27396 16736 27402 16788
rect 30650 16736 30656 16788
rect 30708 16776 30714 16788
rect 31205 16779 31263 16785
rect 31205 16776 31217 16779
rect 30708 16748 31217 16776
rect 30708 16736 30714 16748
rect 31205 16745 31217 16748
rect 31251 16745 31263 16779
rect 31205 16739 31263 16745
rect 22189 16643 22247 16649
rect 22189 16640 22201 16643
rect 22066 16612 22201 16640
rect 20073 16603 20131 16609
rect 22189 16609 22201 16612
rect 22235 16609 22247 16643
rect 26344 16640 26372 16736
rect 26510 16668 26516 16720
rect 26568 16708 26574 16720
rect 28902 16708 28908 16720
rect 26568 16680 28908 16708
rect 26568 16668 26574 16680
rect 27448 16649 27476 16680
rect 28902 16668 28908 16680
rect 28960 16668 28966 16720
rect 29546 16668 29552 16720
rect 29604 16708 29610 16720
rect 29641 16711 29699 16717
rect 29641 16708 29653 16711
rect 29604 16680 29653 16708
rect 29604 16668 29610 16680
rect 29641 16677 29653 16680
rect 29687 16677 29699 16711
rect 31294 16708 31300 16720
rect 30866 16680 31300 16708
rect 29641 16671 29699 16677
rect 31294 16668 31300 16680
rect 31352 16668 31358 16720
rect 26421 16643 26479 16649
rect 26421 16640 26433 16643
rect 26344 16612 26433 16640
rect 22189 16603 22247 16609
rect 26421 16609 26433 16612
rect 26467 16609 26479 16643
rect 26421 16603 26479 16609
rect 27433 16643 27491 16649
rect 27433 16609 27445 16643
rect 27479 16609 27491 16643
rect 27433 16603 27491 16609
rect 17368 16544 17540 16572
rect 17368 16532 17374 16544
rect 17862 16532 17868 16584
rect 17920 16532 17926 16584
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16541 18935 16575
rect 18877 16535 18935 16541
rect 16942 16504 16948 16516
rect 15672 16476 16948 16504
rect 14783 16473 14795 16476
rect 14737 16467 14795 16473
rect 16942 16464 16948 16476
rect 17000 16464 17006 16516
rect 17773 16507 17831 16513
rect 17773 16504 17785 16507
rect 17052 16476 17785 16504
rect 14829 16439 14887 16445
rect 14829 16436 14841 16439
rect 14660 16408 14841 16436
rect 12676 16396 12682 16408
rect 14829 16405 14841 16408
rect 14875 16436 14887 16439
rect 15562 16436 15568 16448
rect 14875 16408 15568 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 15654 16396 15660 16448
rect 15712 16436 15718 16448
rect 15930 16436 15936 16448
rect 15712 16408 15936 16436
rect 15712 16396 15718 16408
rect 15930 16396 15936 16408
rect 15988 16396 15994 16448
rect 16114 16396 16120 16448
rect 16172 16436 16178 16448
rect 17052 16436 17080 16476
rect 17773 16473 17785 16476
rect 17819 16473 17831 16507
rect 17880 16504 17908 16532
rect 18892 16504 18920 16535
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20036 16544 22094 16572
rect 20036 16532 20042 16544
rect 17880 16476 18920 16504
rect 17773 16467 17831 16473
rect 16172 16408 17080 16436
rect 16172 16396 16178 16408
rect 17402 16396 17408 16448
rect 17460 16396 17466 16448
rect 18325 16439 18383 16445
rect 18325 16405 18337 16439
rect 18371 16436 18383 16439
rect 18414 16436 18420 16448
rect 18371 16408 18420 16436
rect 18371 16405 18383 16408
rect 18325 16399 18383 16405
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 22066 16436 22094 16544
rect 29362 16532 29368 16584
rect 29420 16532 29426 16584
rect 31846 16532 31852 16584
rect 31904 16532 31910 16584
rect 30834 16464 30840 16516
rect 30892 16464 30898 16516
rect 30374 16436 30380 16448
rect 22066 16408 30380 16436
rect 30374 16396 30380 16408
rect 30432 16396 30438 16448
rect 30852 16436 30880 16464
rect 31113 16439 31171 16445
rect 31113 16436 31125 16439
rect 30852 16408 31125 16436
rect 31113 16405 31125 16408
rect 31159 16405 31171 16439
rect 31113 16399 31171 16405
rect 2760 16346 32200 16368
rect 2760 16294 6286 16346
rect 6338 16294 6350 16346
rect 6402 16294 6414 16346
rect 6466 16294 6478 16346
rect 6530 16294 6542 16346
rect 6594 16294 13646 16346
rect 13698 16294 13710 16346
rect 13762 16294 13774 16346
rect 13826 16294 13838 16346
rect 13890 16294 13902 16346
rect 13954 16294 21006 16346
rect 21058 16294 21070 16346
rect 21122 16294 21134 16346
rect 21186 16294 21198 16346
rect 21250 16294 21262 16346
rect 21314 16294 28366 16346
rect 28418 16294 28430 16346
rect 28482 16294 28494 16346
rect 28546 16294 28558 16346
rect 28610 16294 28622 16346
rect 28674 16294 32200 16346
rect 2760 16272 32200 16294
rect 11793 16235 11851 16241
rect 11793 16201 11805 16235
rect 11839 16232 11851 16235
rect 12158 16232 12164 16244
rect 11839 16204 12164 16232
rect 11839 16201 11851 16204
rect 11793 16195 11851 16201
rect 12158 16192 12164 16204
rect 12216 16192 12222 16244
rect 13078 16192 13084 16244
rect 13136 16192 13142 16244
rect 13170 16192 13176 16244
rect 13228 16232 13234 16244
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 13228 16204 13645 16232
rect 13228 16192 13234 16204
rect 13633 16201 13645 16204
rect 13679 16201 13691 16235
rect 13633 16195 13691 16201
rect 14182 16192 14188 16244
rect 14240 16192 14246 16244
rect 15010 16232 15016 16244
rect 14384 16204 15016 16232
rect 8297 16167 8355 16173
rect 8297 16164 8309 16167
rect 8220 16136 8309 16164
rect 5626 16056 5632 16108
rect 5684 16096 5690 16108
rect 6181 16099 6239 16105
rect 6181 16096 6193 16099
rect 5684 16068 6193 16096
rect 5684 16056 5690 16068
rect 6181 16065 6193 16068
rect 6227 16096 6239 16099
rect 6638 16096 6644 16108
rect 6227 16068 6644 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 6638 16056 6644 16068
rect 6696 16056 6702 16108
rect 8220 16105 8248 16136
rect 8297 16133 8309 16136
rect 8343 16133 8355 16167
rect 12342 16164 12348 16176
rect 8297 16127 8355 16133
rect 11348 16136 12348 16164
rect 8205 16099 8263 16105
rect 8205 16065 8217 16099
rect 8251 16065 8263 16099
rect 9125 16099 9183 16105
rect 9125 16096 9137 16099
rect 8205 16059 8263 16065
rect 8496 16068 9137 16096
rect 8496 16040 8524 16068
rect 9125 16065 9137 16068
rect 9171 16065 9183 16099
rect 9125 16059 9183 16065
rect 4249 16031 4307 16037
rect 4249 16028 4261 16031
rect 3436 16000 4261 16028
rect 1302 15920 1308 15972
rect 1360 15960 1366 15972
rect 3237 15963 3295 15969
rect 3237 15960 3249 15963
rect 1360 15932 3249 15960
rect 1360 15920 1366 15932
rect 3237 15929 3249 15932
rect 3283 15929 3295 15963
rect 3237 15923 3295 15929
rect 3436 15904 3464 16000
rect 4249 15997 4261 16000
rect 4295 16028 4307 16031
rect 4617 16031 4675 16037
rect 4617 16028 4629 16031
rect 4295 16000 4629 16028
rect 4295 15997 4307 16000
rect 4249 15991 4307 15997
rect 4617 15997 4629 16000
rect 4663 15997 4675 16031
rect 4617 15991 4675 15997
rect 6457 16031 6515 16037
rect 6457 15997 6469 16031
rect 6503 16028 6515 16031
rect 6730 16028 6736 16040
rect 6503 16000 6736 16028
rect 6503 15997 6515 16000
rect 6457 15991 6515 15997
rect 6730 15988 6736 16000
rect 6788 15988 6794 16040
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 6871 16000 7297 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 5261 15963 5319 15969
rect 5261 15929 5273 15963
rect 5307 15960 5319 15963
rect 5810 15960 5816 15972
rect 5307 15932 5816 15960
rect 5307 15929 5319 15932
rect 5261 15923 5319 15929
rect 5810 15920 5816 15932
rect 5868 15920 5874 15972
rect 6178 15920 6184 15972
rect 6236 15960 6242 15972
rect 6840 15960 6868 15991
rect 6236 15932 6868 15960
rect 7300 15960 7328 15991
rect 8478 15988 8484 16040
rect 8536 15988 8542 16040
rect 8849 16031 8907 16037
rect 8849 15997 8861 16031
rect 8895 16028 8907 16031
rect 10962 16028 10968 16040
rect 8895 16000 10968 16028
rect 8895 15997 8907 16000
rect 8849 15991 8907 15997
rect 10962 15988 10968 16000
rect 11020 15988 11026 16040
rect 11348 16037 11376 16136
rect 12342 16124 12348 16136
rect 12400 16124 12406 16176
rect 12526 16124 12532 16176
rect 12584 16124 12590 16176
rect 13817 16167 13875 16173
rect 13817 16133 13829 16167
rect 13863 16164 13875 16167
rect 14200 16164 14228 16192
rect 14384 16173 14412 16204
rect 15010 16192 15016 16204
rect 15068 16232 15074 16244
rect 15289 16235 15347 16241
rect 15289 16232 15301 16235
rect 15068 16204 15301 16232
rect 15068 16192 15074 16204
rect 15289 16201 15301 16204
rect 15335 16201 15347 16235
rect 15289 16195 15347 16201
rect 13863 16136 14228 16164
rect 14369 16167 14427 16173
rect 13863 16133 13875 16136
rect 13817 16127 13875 16133
rect 14369 16133 14381 16167
rect 14415 16133 14427 16167
rect 15304 16164 15332 16195
rect 15470 16192 15476 16244
rect 15528 16232 15534 16244
rect 16666 16232 16672 16244
rect 15528 16204 16672 16232
rect 15528 16192 15534 16204
rect 16666 16192 16672 16204
rect 16724 16192 16730 16244
rect 17402 16232 17408 16244
rect 16776 16204 17408 16232
rect 16776 16164 16804 16204
rect 17402 16192 17408 16204
rect 17460 16192 17466 16244
rect 17589 16235 17647 16241
rect 17589 16201 17601 16235
rect 17635 16232 17647 16235
rect 17678 16232 17684 16244
rect 17635 16204 17684 16232
rect 17635 16201 17647 16204
rect 17589 16195 17647 16201
rect 17678 16192 17684 16204
rect 17736 16192 17742 16244
rect 19889 16235 19947 16241
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 19978 16232 19984 16244
rect 19935 16204 19984 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 22925 16235 22983 16241
rect 22925 16232 22937 16235
rect 22066 16204 22937 16232
rect 15304 16136 16804 16164
rect 14369 16127 14427 16133
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 12253 16099 12311 16105
rect 12253 16096 12265 16099
rect 12124 16068 12265 16096
rect 12124 16056 12130 16068
rect 12253 16065 12265 16068
rect 12299 16096 12311 16099
rect 12299 16068 12572 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 11333 16031 11391 16037
rect 11333 16028 11345 16031
rect 11164 16000 11345 16028
rect 7300 15932 7972 15960
rect 6236 15920 6242 15932
rect 7944 15904 7972 15932
rect 8570 15920 8576 15972
rect 8628 15920 8634 15972
rect 8665 15963 8723 15969
rect 8665 15929 8677 15963
rect 8711 15960 8723 15963
rect 10410 15960 10416 15972
rect 8711 15932 10416 15960
rect 8711 15929 8723 15932
rect 8665 15923 8723 15929
rect 10410 15920 10416 15932
rect 10468 15920 10474 15972
rect 3418 15852 3424 15904
rect 3476 15852 3482 15904
rect 5442 15852 5448 15904
rect 5500 15892 5506 15904
rect 6733 15895 6791 15901
rect 6733 15892 6745 15895
rect 5500 15864 6745 15892
rect 5500 15852 5506 15864
rect 6733 15861 6745 15864
rect 6779 15861 6791 15895
rect 6733 15855 6791 15861
rect 6822 15852 6828 15904
rect 6880 15892 6886 15904
rect 7193 15895 7251 15901
rect 7193 15892 7205 15895
rect 6880 15864 7205 15892
rect 6880 15852 6886 15864
rect 7193 15861 7205 15864
rect 7239 15861 7251 15895
rect 7193 15855 7251 15861
rect 7558 15852 7564 15904
rect 7616 15852 7622 15904
rect 7926 15852 7932 15904
rect 7984 15852 7990 15904
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 11164 15901 11192 16000
rect 11333 15997 11345 16000
rect 11379 15997 11391 16031
rect 11333 15991 11391 15997
rect 11701 16031 11759 16037
rect 11701 15997 11713 16031
rect 11747 16028 11759 16031
rect 11882 16028 11888 16040
rect 11747 16000 11888 16028
rect 11747 15997 11759 16000
rect 11701 15991 11759 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 11977 16031 12035 16037
rect 11977 15997 11989 16031
rect 12023 16028 12035 16031
rect 12434 16028 12440 16040
rect 12023 16000 12440 16028
rect 12023 15997 12035 16000
rect 11977 15991 12035 15997
rect 12434 15988 12440 16000
rect 12492 15988 12498 16040
rect 12544 16037 12572 16068
rect 13446 16056 13452 16108
rect 13504 16096 13510 16108
rect 14384 16096 14412 16127
rect 17126 16124 17132 16176
rect 17184 16124 17190 16176
rect 19794 16124 19800 16176
rect 19852 16164 19858 16176
rect 22066 16164 22094 16204
rect 22925 16201 22937 16204
rect 22971 16201 22983 16235
rect 30006 16232 30012 16244
rect 22925 16195 22983 16201
rect 23492 16204 30012 16232
rect 19852 16136 22094 16164
rect 22557 16167 22615 16173
rect 19852 16124 19858 16136
rect 22557 16133 22569 16167
rect 22603 16164 22615 16167
rect 23106 16164 23112 16176
rect 22603 16136 23112 16164
rect 22603 16133 22615 16136
rect 22557 16127 22615 16133
rect 23106 16124 23112 16136
rect 23164 16124 23170 16176
rect 13504 16068 14412 16096
rect 13504 16056 13510 16068
rect 14642 16056 14648 16108
rect 14700 16096 14706 16108
rect 15286 16096 15292 16108
rect 14700 16068 15292 16096
rect 14700 16056 14706 16068
rect 15286 16056 15292 16068
rect 15344 16056 15350 16108
rect 15488 16068 16160 16096
rect 12529 16031 12587 16037
rect 12529 15997 12541 16031
rect 12575 15997 12587 16031
rect 12529 15991 12587 15997
rect 12618 15988 12624 16040
rect 12676 16028 12682 16040
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 12676 16000 12725 16028
rect 12676 15988 12682 16000
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 13354 15988 13360 16040
rect 13412 16028 13418 16040
rect 13998 16028 14004 16040
rect 13412 16000 14004 16028
rect 13412 15988 13418 16000
rect 13998 15988 14004 16000
rect 14056 15988 14062 16040
rect 13538 15920 13544 15972
rect 13596 15960 13602 15972
rect 14093 15963 14151 15969
rect 14093 15960 14105 15963
rect 13596 15932 14105 15960
rect 13596 15920 13602 15932
rect 14093 15929 14105 15932
rect 14139 15960 14151 15963
rect 14642 15960 14648 15972
rect 14139 15932 14648 15960
rect 14139 15929 14151 15932
rect 14093 15923 14151 15929
rect 14642 15920 14648 15932
rect 14700 15960 14706 15972
rect 15313 15969 15341 16056
rect 15488 16040 15516 16068
rect 15470 15988 15476 16040
rect 15528 15988 15534 16040
rect 15654 15988 15660 16040
rect 15712 15988 15718 16040
rect 16132 16037 16160 16068
rect 16850 16056 16856 16108
rect 16908 16056 16914 16108
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 20956 16068 23397 16096
rect 20956 16056 20962 16068
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 15933 16031 15991 16037
rect 15933 15997 15945 16031
rect 15979 15997 15991 16031
rect 15933 15991 15991 15997
rect 16117 16031 16175 16037
rect 16117 15997 16129 16031
rect 16163 16028 16175 16031
rect 16574 16028 16580 16040
rect 16163 16000 16580 16028
rect 16163 15997 16175 16000
rect 16117 15991 16175 15997
rect 14921 15963 14979 15969
rect 14921 15960 14933 15963
rect 14700 15932 14933 15960
rect 14700 15920 14706 15932
rect 14921 15929 14933 15932
rect 14967 15929 14979 15963
rect 14921 15923 14979 15929
rect 15298 15963 15356 15969
rect 15298 15929 15310 15963
rect 15344 15929 15356 15963
rect 15298 15923 15356 15929
rect 11149 15895 11207 15901
rect 11149 15892 11161 15895
rect 10744 15864 11161 15892
rect 10744 15852 10750 15864
rect 11149 15861 11161 15864
rect 11195 15861 11207 15895
rect 11149 15855 11207 15861
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 12342 15892 12348 15904
rect 11572 15864 12348 15892
rect 11572 15852 11578 15864
rect 12342 15852 12348 15864
rect 12400 15852 12406 15904
rect 14936 15892 14964 15923
rect 15010 15892 15016 15904
rect 14936 15864 15016 15892
rect 15010 15852 15016 15864
rect 15068 15892 15074 15904
rect 15672 15892 15700 15988
rect 15068 15864 15700 15892
rect 15948 15892 15976 15991
rect 16574 15988 16580 16000
rect 16632 15988 16638 16040
rect 16666 15988 16672 16040
rect 16724 16028 16730 16040
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 16724 16000 16957 16028
rect 16724 15988 16730 16000
rect 16945 15997 16957 16000
rect 16991 16028 17003 16031
rect 17865 16031 17923 16037
rect 17865 16028 17877 16031
rect 16991 16000 17877 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17865 15997 17877 16000
rect 17911 15997 17923 16031
rect 17865 15991 17923 15997
rect 18138 15988 18144 16040
rect 18196 15988 18202 16040
rect 23492 16028 23520 16204
rect 30006 16192 30012 16204
rect 30064 16192 30070 16244
rect 31846 16192 31852 16244
rect 31904 16192 31910 16244
rect 24029 16099 24087 16105
rect 24029 16065 24041 16099
rect 24075 16096 24087 16099
rect 25498 16096 25504 16108
rect 24075 16068 25504 16096
rect 24075 16065 24087 16068
rect 24029 16059 24087 16065
rect 25498 16056 25504 16068
rect 25556 16056 25562 16108
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16096 29147 16099
rect 29362 16096 29368 16108
rect 29135 16068 29368 16096
rect 29135 16065 29147 16068
rect 29089 16059 29147 16065
rect 29362 16056 29368 16068
rect 29420 16056 29426 16108
rect 29822 16096 29828 16108
rect 29472 16068 29828 16096
rect 22940 16000 23520 16028
rect 16298 15920 16304 15972
rect 16356 15960 16362 15972
rect 17221 15963 17279 15969
rect 17221 15960 17233 15963
rect 16356 15932 17233 15960
rect 16356 15920 16362 15932
rect 17221 15929 17233 15932
rect 17267 15929 17279 15963
rect 17221 15923 17279 15929
rect 17635 15963 17693 15969
rect 17635 15929 17647 15963
rect 17681 15960 17693 15963
rect 17770 15960 17776 15972
rect 17681 15932 17776 15960
rect 17681 15929 17693 15932
rect 17635 15923 17693 15929
rect 17770 15920 17776 15932
rect 17828 15920 17834 15972
rect 19150 15920 19156 15972
rect 19208 15920 19214 15972
rect 17034 15892 17040 15904
rect 15948 15864 17040 15892
rect 15068 15852 15074 15864
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 22940 15901 22968 16000
rect 24118 15988 24124 16040
rect 24176 15988 24182 16040
rect 26602 15988 26608 16040
rect 26660 16028 26666 16040
rect 29472 16037 29500 16068
rect 29822 16056 29828 16068
rect 29880 16056 29886 16108
rect 26881 16031 26939 16037
rect 26881 16028 26893 16031
rect 26660 16000 26893 16028
rect 26660 15988 26666 16000
rect 26881 15997 26893 16000
rect 26927 15997 26939 16031
rect 26881 15991 26939 15997
rect 29457 16031 29515 16037
rect 29457 15997 29469 16031
rect 29503 15997 29515 16031
rect 29457 15991 29515 15997
rect 30883 16031 30941 16037
rect 30883 15997 30895 16031
rect 30929 16028 30941 16031
rect 31205 16031 31263 16037
rect 31205 16028 31217 16031
rect 30929 16000 31217 16028
rect 30929 15997 30941 16000
rect 30883 15991 30941 15997
rect 31205 15997 31217 16000
rect 31251 15997 31263 16031
rect 31205 15991 31263 15997
rect 30190 15920 30196 15972
rect 30248 15920 30254 15972
rect 22925 15895 22983 15901
rect 22925 15861 22937 15895
rect 22971 15861 22983 15895
rect 22925 15855 22983 15861
rect 23109 15895 23167 15901
rect 23109 15861 23121 15895
rect 23155 15892 23167 15895
rect 24394 15892 24400 15904
rect 23155 15864 24400 15892
rect 23155 15861 23167 15864
rect 23109 15855 23167 15861
rect 24394 15852 24400 15864
rect 24452 15852 24458 15904
rect 24578 15852 24584 15904
rect 24636 15892 24642 15904
rect 24765 15895 24823 15901
rect 24765 15892 24777 15895
rect 24636 15864 24777 15892
rect 24636 15852 24642 15864
rect 24765 15861 24777 15864
rect 24811 15861 24823 15895
rect 24765 15855 24823 15861
rect 26326 15852 26332 15904
rect 26384 15852 26390 15904
rect 2760 15802 32200 15824
rect 2760 15750 6946 15802
rect 6998 15750 7010 15802
rect 7062 15750 7074 15802
rect 7126 15750 7138 15802
rect 7190 15750 7202 15802
rect 7254 15750 14306 15802
rect 14358 15750 14370 15802
rect 14422 15750 14434 15802
rect 14486 15750 14498 15802
rect 14550 15750 14562 15802
rect 14614 15750 21666 15802
rect 21718 15750 21730 15802
rect 21782 15750 21794 15802
rect 21846 15750 21858 15802
rect 21910 15750 21922 15802
rect 21974 15750 29026 15802
rect 29078 15750 29090 15802
rect 29142 15750 29154 15802
rect 29206 15750 29218 15802
rect 29270 15750 29282 15802
rect 29334 15750 32200 15802
rect 2760 15728 32200 15750
rect 3418 15648 3424 15700
rect 3476 15648 3482 15700
rect 5442 15688 5448 15700
rect 4816 15660 5448 15688
rect 4816 15620 4844 15660
rect 5442 15648 5448 15660
rect 5500 15648 5506 15700
rect 6822 15688 6828 15700
rect 6380 15660 6828 15688
rect 4462 15592 4844 15620
rect 4893 15623 4951 15629
rect 4893 15589 4905 15623
rect 4939 15620 4951 15623
rect 5258 15620 5264 15632
rect 4939 15592 5264 15620
rect 4939 15589 4951 15592
rect 4893 15583 4951 15589
rect 5258 15580 5264 15592
rect 5316 15580 5322 15632
rect 6380 15620 6408 15660
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 12069 15691 12127 15697
rect 12069 15657 12081 15691
rect 12115 15688 12127 15691
rect 12250 15688 12256 15700
rect 12115 15660 12256 15688
rect 12115 15657 12127 15660
rect 12069 15651 12127 15657
rect 12250 15648 12256 15660
rect 12308 15648 12314 15700
rect 12342 15648 12348 15700
rect 12400 15688 12406 15700
rect 12400 15660 13124 15688
rect 12400 15648 12406 15660
rect 6302 15592 6408 15620
rect 6733 15623 6791 15629
rect 6733 15589 6745 15623
rect 6779 15620 6791 15623
rect 7101 15623 7159 15629
rect 7101 15620 7113 15623
rect 6779 15592 7113 15620
rect 6779 15589 6791 15592
rect 6733 15583 6791 15589
rect 7101 15589 7113 15592
rect 7147 15589 7159 15623
rect 7101 15583 7159 15589
rect 12158 15580 12164 15632
rect 12216 15620 12222 15632
rect 12216 15592 12664 15620
rect 12216 15580 12222 15592
rect 12636 15564 12664 15592
rect 11054 15512 11060 15564
rect 11112 15512 11118 15564
rect 11146 15512 11152 15564
rect 11204 15512 11210 15564
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15552 11391 15555
rect 12342 15552 12348 15564
rect 11379 15524 12348 15552
rect 11379 15521 11391 15524
rect 11333 15515 11391 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 12618 15512 12624 15564
rect 12676 15512 12682 15564
rect 12802 15512 12808 15564
rect 12860 15512 12866 15564
rect 12894 15512 12900 15564
rect 12952 15512 12958 15564
rect 5169 15487 5227 15493
rect 5169 15453 5181 15487
rect 5215 15484 5227 15487
rect 5442 15484 5448 15496
rect 5215 15456 5448 15484
rect 5215 15453 5227 15456
rect 5169 15447 5227 15453
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 7282 15484 7288 15496
rect 7055 15456 7288 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 7282 15444 7288 15456
rect 7340 15444 7346 15496
rect 7650 15444 7656 15496
rect 7708 15444 7714 15496
rect 9030 15444 9036 15496
rect 9088 15444 9094 15496
rect 11517 15487 11575 15493
rect 11517 15453 11529 15487
rect 11563 15484 11575 15487
rect 11790 15484 11796 15496
rect 11563 15456 11796 15484
rect 11563 15453 11575 15456
rect 11517 15447 11575 15453
rect 11790 15444 11796 15456
rect 11848 15484 11854 15496
rect 12526 15484 12532 15496
rect 11848 15456 12532 15484
rect 11848 15444 11854 15456
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 12820 15416 12848 15512
rect 13096 15484 13124 15660
rect 13170 15648 13176 15700
rect 13228 15648 13234 15700
rect 14182 15648 14188 15700
rect 14240 15648 14246 15700
rect 14642 15648 14648 15700
rect 14700 15648 14706 15700
rect 15286 15648 15292 15700
rect 15344 15648 15350 15700
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 17773 15691 17831 15697
rect 17773 15688 17785 15691
rect 17552 15660 17785 15688
rect 17552 15648 17558 15660
rect 17773 15657 17785 15660
rect 17819 15657 17831 15691
rect 17773 15651 17831 15657
rect 19150 15648 19156 15700
rect 19208 15688 19214 15700
rect 19245 15691 19303 15697
rect 19245 15688 19257 15691
rect 19208 15660 19257 15688
rect 19208 15648 19214 15660
rect 19245 15657 19257 15660
rect 19291 15657 19303 15691
rect 19245 15651 19303 15657
rect 19981 15691 20039 15697
rect 19981 15657 19993 15691
rect 20027 15657 20039 15691
rect 23106 15688 23112 15700
rect 19981 15651 20039 15657
rect 21192 15660 23112 15688
rect 13188 15561 13216 15648
rect 13262 15580 13268 15632
rect 13320 15580 13326 15632
rect 13909 15623 13967 15629
rect 13909 15589 13921 15623
rect 13955 15620 13967 15623
rect 14200 15620 14228 15648
rect 14660 15620 14688 15648
rect 13955 15592 14136 15620
rect 14200 15592 14320 15620
rect 13955 15589 13967 15592
rect 13909 15583 13967 15589
rect 14108 15564 14136 15592
rect 13173 15555 13231 15561
rect 13173 15521 13185 15555
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 13372 15484 13400 15515
rect 13998 15512 14004 15564
rect 14056 15512 14062 15564
rect 14090 15512 14096 15564
rect 14148 15512 14154 15564
rect 14182 15512 14188 15564
rect 14240 15512 14246 15564
rect 14292 15561 14320 15592
rect 14568 15592 14688 15620
rect 15304 15620 15332 15648
rect 15654 15620 15660 15632
rect 15304 15592 15660 15620
rect 14568 15561 14596 15592
rect 15654 15580 15660 15592
rect 15712 15620 15718 15632
rect 15712 15592 15976 15620
rect 15712 15580 15718 15592
rect 14277 15555 14335 15561
rect 14277 15521 14289 15555
rect 14323 15521 14335 15555
rect 14277 15515 14335 15521
rect 14553 15555 14611 15561
rect 14553 15521 14565 15555
rect 14599 15521 14611 15555
rect 14553 15515 14611 15521
rect 14645 15555 14703 15561
rect 14645 15521 14657 15555
rect 14691 15552 14703 15555
rect 14826 15552 14832 15564
rect 14691 15524 14832 15552
rect 14691 15521 14703 15524
rect 14645 15515 14703 15521
rect 14826 15512 14832 15524
rect 14884 15512 14890 15564
rect 15013 15555 15071 15561
rect 15013 15521 15025 15555
rect 15059 15552 15071 15555
rect 15059 15524 15332 15552
rect 15059 15521 15071 15524
rect 15013 15515 15071 15521
rect 15194 15484 15200 15496
rect 13096 15456 15200 15484
rect 15194 15444 15200 15456
rect 15252 15444 15258 15496
rect 15304 15484 15332 15524
rect 15378 15512 15384 15564
rect 15436 15512 15442 15564
rect 15562 15512 15568 15564
rect 15620 15512 15626 15564
rect 15948 15561 15976 15592
rect 16132 15592 16804 15620
rect 16132 15564 16160 15592
rect 15933 15555 15991 15561
rect 15933 15521 15945 15555
rect 15979 15521 15991 15555
rect 15933 15515 15991 15521
rect 16114 15512 16120 15564
rect 16172 15512 16178 15564
rect 16666 15512 16672 15564
rect 16724 15512 16730 15564
rect 16776 15552 16804 15592
rect 17034 15580 17040 15632
rect 17092 15620 17098 15632
rect 19797 15623 19855 15629
rect 17092 15592 17724 15620
rect 17092 15580 17098 15592
rect 17129 15555 17187 15561
rect 17129 15552 17141 15555
rect 16776 15524 17141 15552
rect 17129 15521 17141 15524
rect 17175 15521 17187 15555
rect 17129 15515 17187 15521
rect 17218 15512 17224 15564
rect 17276 15512 17282 15564
rect 15838 15484 15844 15496
rect 15304 15456 15844 15484
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16574 15444 16580 15496
rect 16632 15444 16638 15496
rect 17017 15487 17075 15493
rect 17017 15453 17029 15487
rect 17063 15484 17075 15487
rect 17236 15484 17264 15512
rect 17063 15456 17264 15484
rect 17405 15487 17463 15493
rect 17063 15453 17075 15456
rect 17017 15447 17075 15453
rect 17405 15453 17417 15487
rect 17451 15453 17463 15487
rect 17405 15447 17463 15453
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15484 17555 15487
rect 17696 15484 17724 15592
rect 19797 15589 19809 15623
rect 19843 15589 19855 15623
rect 19797 15583 19855 15589
rect 19153 15555 19211 15561
rect 19153 15521 19165 15555
rect 19199 15521 19211 15555
rect 19153 15515 19211 15521
rect 17543 15456 17724 15484
rect 17543 15453 17555 15456
rect 17497 15447 17555 15453
rect 14829 15419 14887 15425
rect 14829 15416 14841 15419
rect 12820 15388 14841 15416
rect 14829 15385 14841 15388
rect 14875 15416 14887 15419
rect 15562 15416 15568 15428
rect 14875 15388 15568 15416
rect 14875 15385 14887 15388
rect 14829 15379 14887 15385
rect 15562 15376 15568 15388
rect 15620 15376 15626 15428
rect 5261 15351 5319 15357
rect 5261 15317 5273 15351
rect 5307 15348 5319 15351
rect 5718 15348 5724 15360
rect 5307 15320 5724 15348
rect 5307 15317 5319 15320
rect 5261 15311 5319 15317
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 8481 15351 8539 15357
rect 8481 15317 8493 15351
rect 8527 15348 8539 15351
rect 8570 15348 8576 15360
rect 8527 15320 8576 15348
rect 8527 15317 8539 15320
rect 8481 15311 8539 15317
rect 8570 15308 8576 15320
rect 8628 15348 8634 15360
rect 8938 15348 8944 15360
rect 8628 15320 8944 15348
rect 8628 15308 8634 15320
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 10873 15351 10931 15357
rect 10873 15348 10885 15351
rect 10744 15320 10885 15348
rect 10744 15308 10750 15320
rect 10873 15317 10885 15320
rect 10919 15317 10931 15351
rect 10873 15311 10931 15317
rect 10962 15308 10968 15360
rect 11020 15348 11026 15360
rect 11333 15351 11391 15357
rect 11333 15348 11345 15351
rect 11020 15320 11345 15348
rect 11020 15308 11026 15320
rect 11333 15317 11345 15320
rect 11379 15317 11391 15351
rect 11333 15311 11391 15317
rect 11790 15308 11796 15360
rect 11848 15348 11854 15360
rect 11974 15348 11980 15360
rect 11848 15320 11980 15348
rect 11848 15308 11854 15320
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12158 15308 12164 15360
rect 12216 15348 12222 15360
rect 12437 15351 12495 15357
rect 12437 15348 12449 15351
rect 12216 15320 12449 15348
rect 12216 15308 12222 15320
rect 12437 15317 12449 15320
rect 12483 15317 12495 15351
rect 12437 15311 12495 15317
rect 13998 15308 14004 15360
rect 14056 15308 14062 15360
rect 14182 15308 14188 15360
rect 14240 15348 14246 15360
rect 15470 15348 15476 15360
rect 14240 15320 15476 15348
rect 14240 15308 14246 15320
rect 15470 15308 15476 15320
rect 15528 15308 15534 15360
rect 15856 15348 15884 15444
rect 16592 15416 16620 15444
rect 17420 15416 17448 15447
rect 16592 15388 17448 15416
rect 17512 15416 17540 15447
rect 19168 15428 19196 15515
rect 19812 15484 19840 15583
rect 19996 15552 20024 15651
rect 21085 15555 21143 15561
rect 21085 15552 21097 15555
rect 19996 15524 21097 15552
rect 21085 15521 21097 15524
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 21192 15552 21220 15660
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 23293 15691 23351 15697
rect 23293 15657 23305 15691
rect 23339 15688 23351 15691
rect 24118 15688 24124 15700
rect 23339 15660 24124 15688
rect 23339 15657 23351 15660
rect 23293 15651 23351 15657
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 24394 15648 24400 15700
rect 24452 15648 24458 15700
rect 30190 15648 30196 15700
rect 30248 15648 30254 15700
rect 30466 15648 30472 15700
rect 30524 15648 30530 15700
rect 21269 15623 21327 15629
rect 21269 15589 21281 15623
rect 21315 15620 21327 15623
rect 21542 15620 21548 15632
rect 21315 15592 21548 15620
rect 21315 15589 21327 15592
rect 21269 15583 21327 15589
rect 21542 15580 21548 15592
rect 21600 15580 21606 15632
rect 23566 15620 23572 15632
rect 23046 15592 23572 15620
rect 23566 15580 23572 15592
rect 23624 15580 23630 15632
rect 21361 15555 21419 15561
rect 21361 15552 21373 15555
rect 21192 15524 21373 15552
rect 20530 15484 20536 15496
rect 19812 15456 20536 15484
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 20763 15456 20913 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 20901 15453 20913 15456
rect 20947 15453 20959 15487
rect 20901 15447 20959 15453
rect 17586 15416 17592 15428
rect 17512 15388 17592 15416
rect 17586 15376 17592 15388
rect 17644 15376 17650 15428
rect 19150 15376 19156 15428
rect 19208 15376 19214 15428
rect 19429 15419 19487 15425
rect 19429 15416 19441 15419
rect 19306 15388 19441 15416
rect 16853 15351 16911 15357
rect 16853 15348 16865 15351
rect 15856 15320 16865 15348
rect 16853 15317 16865 15320
rect 16899 15317 16911 15351
rect 16853 15311 16911 15317
rect 17494 15308 17500 15360
rect 17552 15348 17558 15360
rect 19306 15348 19334 15388
rect 19429 15385 19441 15388
rect 19475 15416 19487 15419
rect 21192 15416 21220 15524
rect 21361 15521 21373 15524
rect 21407 15521 21419 15555
rect 21361 15515 21419 15521
rect 23106 15512 23112 15564
rect 23164 15552 23170 15564
rect 24412 15561 24440 15648
rect 26050 15620 26056 15632
rect 25884 15592 26056 15620
rect 24397 15555 24455 15561
rect 23164 15524 24348 15552
rect 23164 15512 23170 15524
rect 21545 15487 21603 15493
rect 21545 15484 21557 15487
rect 19475 15388 21220 15416
rect 21376 15456 21557 15484
rect 19475 15385 19487 15388
rect 19429 15379 19487 15385
rect 21376 15360 21404 15456
rect 21545 15453 21557 15456
rect 21591 15453 21603 15487
rect 21545 15447 21603 15453
rect 21821 15487 21879 15493
rect 21821 15453 21833 15487
rect 21867 15484 21879 15487
rect 23477 15487 23535 15493
rect 23477 15484 23489 15487
rect 21867 15456 23489 15484
rect 21867 15453 21879 15456
rect 21821 15447 21879 15453
rect 23477 15453 23489 15456
rect 23523 15453 23535 15487
rect 23477 15447 23535 15453
rect 24121 15487 24179 15493
rect 24121 15453 24133 15487
rect 24167 15484 24179 15487
rect 24213 15487 24271 15493
rect 24213 15484 24225 15487
rect 24167 15456 24225 15484
rect 24167 15453 24179 15456
rect 24121 15447 24179 15453
rect 24213 15453 24225 15456
rect 24259 15453 24271 15487
rect 24320 15484 24348 15524
rect 24397 15521 24409 15555
rect 24443 15521 24455 15555
rect 24397 15515 24455 15521
rect 24578 15512 24584 15564
rect 24636 15512 24642 15564
rect 25884 15561 25912 15592
rect 26050 15580 26056 15592
rect 26108 15580 26114 15632
rect 27798 15620 27804 15632
rect 27370 15592 27804 15620
rect 27798 15580 27804 15592
rect 27856 15580 27862 15632
rect 30484 15620 30512 15648
rect 30742 15620 30748 15632
rect 30300 15592 30748 15620
rect 30300 15561 30328 15592
rect 30742 15580 30748 15592
rect 30800 15580 30806 15632
rect 31665 15623 31723 15629
rect 31665 15589 31677 15623
rect 31711 15620 31723 15623
rect 33134 15620 33140 15632
rect 31711 15592 33140 15620
rect 31711 15589 31723 15592
rect 31665 15583 31723 15589
rect 33134 15580 33140 15592
rect 33192 15580 33198 15632
rect 24673 15555 24731 15561
rect 24673 15521 24685 15555
rect 24719 15521 24731 15555
rect 24673 15515 24731 15521
rect 25869 15555 25927 15561
rect 25869 15521 25881 15555
rect 25915 15521 25927 15555
rect 25869 15515 25927 15521
rect 27709 15555 27767 15561
rect 27709 15521 27721 15555
rect 27755 15521 27767 15555
rect 27709 15515 27767 15521
rect 30285 15555 30343 15561
rect 30285 15521 30297 15555
rect 30331 15521 30343 15555
rect 30285 15515 30343 15521
rect 24688 15484 24716 15515
rect 24320 15456 24716 15484
rect 26145 15487 26203 15493
rect 24213 15447 24271 15453
rect 26145 15453 26157 15487
rect 26191 15484 26203 15487
rect 26878 15484 26884 15496
rect 26191 15456 26884 15484
rect 26191 15453 26203 15456
rect 26145 15447 26203 15453
rect 26878 15444 26884 15456
rect 26936 15444 26942 15496
rect 27617 15419 27675 15425
rect 27617 15385 27629 15419
rect 27663 15416 27675 15419
rect 27724 15416 27752 15515
rect 30374 15512 30380 15564
rect 30432 15552 30438 15564
rect 30469 15555 30527 15561
rect 30469 15552 30481 15555
rect 30432 15524 30481 15552
rect 30432 15512 30438 15524
rect 30469 15521 30481 15524
rect 30515 15521 30527 15555
rect 30469 15515 30527 15521
rect 27663 15388 28212 15416
rect 27663 15385 27675 15388
rect 27617 15379 27675 15385
rect 28184 15360 28212 15388
rect 17552 15320 19334 15348
rect 17552 15308 17558 15320
rect 19518 15308 19524 15360
rect 19576 15348 19582 15360
rect 19794 15348 19800 15360
rect 19576 15320 19800 15348
rect 19576 15308 19582 15320
rect 19794 15308 19800 15320
rect 19852 15308 19858 15360
rect 19886 15308 19892 15360
rect 19944 15348 19950 15360
rect 20073 15351 20131 15357
rect 20073 15348 20085 15351
rect 19944 15320 20085 15348
rect 19944 15308 19950 15320
rect 20073 15317 20085 15320
rect 20119 15317 20131 15351
rect 20073 15311 20131 15317
rect 21358 15308 21364 15360
rect 21416 15308 21422 15360
rect 22462 15308 22468 15360
rect 22520 15348 22526 15360
rect 24578 15348 24584 15360
rect 22520 15320 24584 15348
rect 22520 15308 22526 15320
rect 24578 15308 24584 15320
rect 24636 15308 24642 15360
rect 27893 15351 27951 15357
rect 27893 15317 27905 15351
rect 27939 15348 27951 15351
rect 27982 15348 27988 15360
rect 27939 15320 27988 15348
rect 27939 15317 27951 15320
rect 27893 15311 27951 15317
rect 27982 15308 27988 15320
rect 28040 15308 28046 15360
rect 28166 15308 28172 15360
rect 28224 15308 28230 15360
rect 2760 15258 32200 15280
rect 2760 15206 6286 15258
rect 6338 15206 6350 15258
rect 6402 15206 6414 15258
rect 6466 15206 6478 15258
rect 6530 15206 6542 15258
rect 6594 15206 13646 15258
rect 13698 15206 13710 15258
rect 13762 15206 13774 15258
rect 13826 15206 13838 15258
rect 13890 15206 13902 15258
rect 13954 15206 21006 15258
rect 21058 15206 21070 15258
rect 21122 15206 21134 15258
rect 21186 15206 21198 15258
rect 21250 15206 21262 15258
rect 21314 15206 28366 15258
rect 28418 15206 28430 15258
rect 28482 15206 28494 15258
rect 28546 15206 28558 15258
rect 28610 15206 28622 15258
rect 28674 15206 32200 15258
rect 2760 15184 32200 15206
rect 5902 15104 5908 15156
rect 5960 15144 5966 15156
rect 6181 15147 6239 15153
rect 6181 15144 6193 15147
rect 5960 15116 6193 15144
rect 5960 15104 5966 15116
rect 6181 15113 6193 15116
rect 6227 15113 6239 15147
rect 7374 15144 7380 15156
rect 6181 15107 6239 15113
rect 7116 15116 7380 15144
rect 7116 15076 7144 15116
rect 7374 15104 7380 15116
rect 7432 15104 7438 15156
rect 8757 15147 8815 15153
rect 8757 15113 8769 15147
rect 8803 15144 8815 15147
rect 9030 15144 9036 15156
rect 8803 15116 9036 15144
rect 8803 15113 8815 15116
rect 8757 15107 8815 15113
rect 9030 15104 9036 15116
rect 9088 15104 9094 15156
rect 9214 15104 9220 15156
rect 9272 15144 9278 15156
rect 9950 15144 9956 15156
rect 9272 15116 9956 15144
rect 9272 15104 9278 15116
rect 9950 15104 9956 15116
rect 10008 15144 10014 15156
rect 11057 15147 11115 15153
rect 11057 15144 11069 15147
rect 10008 15116 11069 15144
rect 10008 15104 10014 15116
rect 11057 15113 11069 15116
rect 11103 15113 11115 15147
rect 11057 15107 11115 15113
rect 11974 15104 11980 15156
rect 12032 15144 12038 15156
rect 12253 15147 12311 15153
rect 12253 15144 12265 15147
rect 12032 15116 12265 15144
rect 12032 15104 12038 15116
rect 12253 15113 12265 15116
rect 12299 15144 12311 15147
rect 12802 15144 12808 15156
rect 12299 15116 12808 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 13446 15144 13452 15156
rect 12952 15116 13452 15144
rect 12952 15104 12958 15116
rect 13446 15104 13452 15116
rect 13504 15104 13510 15156
rect 15378 15104 15384 15156
rect 15436 15104 15442 15156
rect 16850 15104 16856 15156
rect 16908 15104 16914 15156
rect 17034 15104 17040 15156
rect 17092 15104 17098 15156
rect 17954 15104 17960 15156
rect 18012 15104 18018 15156
rect 19242 15104 19248 15156
rect 19300 15144 19306 15156
rect 19300 15116 22094 15144
rect 19300 15104 19306 15116
rect 4908 15048 7144 15076
rect 4908 15017 4936 15048
rect 10870 15036 10876 15088
rect 10928 15076 10934 15088
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 10928 15048 11897 15076
rect 10928 15036 10934 15048
rect 11885 15045 11897 15048
rect 11931 15045 11943 15079
rect 11885 15039 11943 15045
rect 12621 15079 12679 15085
rect 12621 15045 12633 15079
rect 12667 15076 12679 15079
rect 12986 15076 12992 15088
rect 12667 15048 12992 15076
rect 12667 15045 12679 15048
rect 12621 15039 12679 15045
rect 12986 15036 12992 15048
rect 13044 15036 13050 15088
rect 17972 15076 18000 15104
rect 15580 15048 18000 15076
rect 22066 15076 22094 15116
rect 22554 15104 22560 15156
rect 22612 15144 22618 15156
rect 23753 15147 23811 15153
rect 23753 15144 23765 15147
rect 22612 15116 23765 15144
rect 22612 15104 22618 15116
rect 23753 15113 23765 15116
rect 23799 15113 23811 15147
rect 23753 15107 23811 15113
rect 26878 15104 26884 15156
rect 26936 15144 26942 15156
rect 27893 15147 27951 15153
rect 27893 15144 27905 15147
rect 26936 15116 27905 15144
rect 26936 15104 26942 15116
rect 27893 15113 27905 15116
rect 27939 15113 27951 15147
rect 27893 15107 27951 15113
rect 31294 15104 31300 15156
rect 31352 15104 31358 15156
rect 29549 15079 29607 15085
rect 22066 15048 25636 15076
rect 4893 15011 4951 15017
rect 4893 14977 4905 15011
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5626 15008 5632 15020
rect 5123 14980 5632 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 6273 15011 6331 15017
rect 6273 15008 6285 15011
rect 5776 14980 6285 15008
rect 5776 14968 5782 14980
rect 6273 14977 6285 14980
rect 6319 14977 6331 15011
rect 6273 14971 6331 14977
rect 7009 15011 7067 15017
rect 7009 14977 7021 15011
rect 7055 15008 7067 15011
rect 7282 15008 7288 15020
rect 7055 14980 7288 15008
rect 7055 14977 7067 14980
rect 7009 14971 7067 14977
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 10686 14968 10692 15020
rect 10744 15008 10750 15020
rect 10965 15011 11023 15017
rect 10965 15008 10977 15011
rect 10744 14980 10977 15008
rect 10744 14968 10750 14980
rect 10965 14977 10977 14980
rect 11011 15008 11023 15011
rect 11011 14980 11560 15008
rect 11011 14977 11023 14980
rect 10965 14971 11023 14977
rect 11532 14952 11560 14980
rect 12526 14968 12532 15020
rect 12584 15008 12590 15020
rect 12584 14980 14044 15008
rect 12584 14968 12590 14980
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14940 3847 14943
rect 3835 14912 4292 14940
rect 3835 14909 3847 14912
rect 3789 14903 3847 14909
rect 4264 14816 4292 14912
rect 5810 14900 5816 14952
rect 5868 14900 5874 14952
rect 6086 14900 6092 14952
rect 6144 14900 6150 14952
rect 11241 14943 11299 14949
rect 11241 14909 11253 14943
rect 11287 14940 11299 14943
rect 11330 14940 11336 14952
rect 11287 14912 11336 14940
rect 11287 14909 11299 14912
rect 11241 14903 11299 14909
rect 11330 14900 11336 14912
rect 11388 14900 11394 14952
rect 11514 14900 11520 14952
rect 11572 14900 11578 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 11790 14940 11796 14952
rect 11655 14912 11796 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 11790 14900 11796 14912
rect 11848 14900 11854 14952
rect 11977 14943 12035 14949
rect 11977 14940 11989 14943
rect 11900 14912 11989 14940
rect 4341 14875 4399 14881
rect 4341 14841 4353 14875
rect 4387 14872 4399 14875
rect 4801 14875 4859 14881
rect 4801 14872 4813 14875
rect 4387 14844 4813 14872
rect 4387 14841 4399 14844
rect 4341 14835 4399 14841
rect 4801 14841 4813 14844
rect 4847 14841 4859 14875
rect 6104 14872 6132 14900
rect 11900 14884 11928 14912
rect 11977 14909 11989 14912
rect 12023 14909 12035 14943
rect 11977 14903 12035 14909
rect 13078 14900 13084 14952
rect 13136 14949 13142 14952
rect 13136 14943 13185 14949
rect 13136 14909 13139 14943
rect 13173 14909 13185 14943
rect 13136 14903 13185 14909
rect 13136 14900 13142 14903
rect 13354 14900 13360 14952
rect 13412 14900 13418 14952
rect 14016 14949 14044 14980
rect 14108 14980 14964 15008
rect 14001 14943 14059 14949
rect 14001 14909 14013 14943
rect 14047 14909 14059 14943
rect 14001 14903 14059 14909
rect 7285 14875 7343 14881
rect 6104 14844 7236 14872
rect 4801 14835 4859 14841
rect 4246 14764 4252 14816
rect 4304 14764 4310 14816
rect 4430 14764 4436 14816
rect 4488 14764 4494 14816
rect 5721 14807 5779 14813
rect 5721 14773 5733 14807
rect 5767 14804 5779 14807
rect 6546 14804 6552 14816
rect 5767 14776 6552 14804
rect 5767 14773 5779 14776
rect 5721 14767 5779 14773
rect 6546 14764 6552 14776
rect 6604 14804 6610 14816
rect 6917 14807 6975 14813
rect 6917 14804 6929 14807
rect 6604 14776 6929 14804
rect 6604 14764 6610 14776
rect 6917 14773 6929 14776
rect 6963 14773 6975 14807
rect 7208 14804 7236 14844
rect 7285 14841 7297 14875
rect 7331 14872 7343 14875
rect 7558 14872 7564 14884
rect 7331 14844 7564 14872
rect 7331 14841 7343 14844
rect 7285 14835 7343 14841
rect 7558 14832 7564 14844
rect 7616 14832 7622 14884
rect 8018 14832 8024 14884
rect 8076 14832 8082 14884
rect 11882 14872 11888 14884
rect 11256 14844 11888 14872
rect 11256 14816 11284 14844
rect 11882 14832 11888 14844
rect 11940 14832 11946 14884
rect 12253 14875 12311 14881
rect 12253 14841 12265 14875
rect 12299 14872 12311 14875
rect 13372 14872 13400 14900
rect 14108 14872 14136 14980
rect 14936 14952 14964 14980
rect 14642 14900 14648 14952
rect 14700 14900 14706 14952
rect 14826 14900 14832 14952
rect 14884 14900 14890 14952
rect 14918 14900 14924 14952
rect 14976 14900 14982 14952
rect 15105 14943 15163 14949
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15470 14940 15476 14952
rect 15151 14912 15476 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15470 14900 15476 14912
rect 15528 14900 15534 14952
rect 15580 14949 15608 15048
rect 15838 14968 15844 15020
rect 15896 15008 15902 15020
rect 17405 15011 17463 15017
rect 15896 14980 16344 15008
rect 15896 14968 15902 14980
rect 15565 14943 15623 14949
rect 15565 14909 15577 14943
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 15933 14943 15991 14949
rect 15933 14909 15945 14943
rect 15979 14909 15991 14943
rect 15933 14903 15991 14909
rect 12299 14844 12848 14872
rect 13372 14844 14136 14872
rect 14844 14872 14872 14900
rect 15948 14872 15976 14903
rect 16114 14900 16120 14952
rect 16172 14900 16178 14952
rect 16316 14949 16344 14980
rect 17405 14977 17417 15011
rect 17451 15008 17463 15011
rect 17586 15008 17592 15020
rect 17451 14980 17592 15008
rect 17451 14977 17463 14980
rect 17405 14971 17463 14977
rect 17586 14968 17592 14980
rect 17644 15008 17650 15020
rect 17644 14980 18000 15008
rect 17644 14968 17650 14980
rect 16301 14943 16359 14949
rect 16301 14909 16313 14943
rect 16347 14909 16359 14943
rect 16761 14943 16819 14949
rect 16761 14940 16773 14943
rect 16301 14903 16359 14909
rect 16500 14912 16773 14940
rect 14844 14844 16160 14872
rect 12299 14841 12311 14844
rect 12253 14835 12311 14841
rect 12820 14816 12848 14844
rect 16132 14816 16160 14844
rect 9030 14804 9036 14816
rect 7208 14776 9036 14804
rect 6917 14767 6975 14773
rect 9030 14764 9036 14776
rect 9088 14804 9094 14816
rect 9309 14807 9367 14813
rect 9309 14804 9321 14807
rect 9088 14776 9321 14804
rect 9088 14764 9094 14776
rect 9309 14773 9321 14776
rect 9355 14804 9367 14807
rect 10778 14804 10784 14816
rect 9355 14776 10784 14804
rect 9355 14773 9367 14776
rect 9309 14767 9367 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 11238 14764 11244 14816
rect 11296 14764 11302 14816
rect 11330 14764 11336 14816
rect 11388 14764 11394 14816
rect 12069 14807 12127 14813
rect 12069 14773 12081 14807
rect 12115 14804 12127 14807
rect 12342 14804 12348 14816
rect 12115 14776 12348 14804
rect 12115 14773 12127 14776
rect 12069 14767 12127 14773
rect 12342 14764 12348 14776
rect 12400 14764 12406 14816
rect 12802 14764 12808 14816
rect 12860 14764 12866 14816
rect 12989 14807 13047 14813
rect 12989 14773 13001 14807
rect 13035 14804 13047 14807
rect 13078 14804 13084 14816
rect 13035 14776 13084 14804
rect 13035 14773 13047 14776
rect 12989 14767 13047 14773
rect 13078 14764 13084 14776
rect 13136 14804 13142 14816
rect 13538 14804 13544 14816
rect 13136 14776 13544 14804
rect 13136 14764 13142 14776
rect 13538 14764 13544 14776
rect 13596 14804 13602 14816
rect 15746 14804 15752 14816
rect 13596 14776 15752 14804
rect 13596 14764 13602 14776
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 16114 14764 16120 14816
rect 16172 14764 16178 14816
rect 16206 14764 16212 14816
rect 16264 14804 16270 14816
rect 16500 14804 16528 14912
rect 16761 14909 16773 14912
rect 16807 14940 16819 14943
rect 17494 14940 17500 14952
rect 16807 14912 17500 14940
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 17494 14900 17500 14912
rect 17552 14900 17558 14952
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17604 14912 17877 14940
rect 16574 14832 16580 14884
rect 16632 14872 16638 14884
rect 17604 14872 17632 14912
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17972 14940 18000 14980
rect 18138 14968 18144 15020
rect 18196 15008 18202 15020
rect 18969 15011 19027 15017
rect 18969 15008 18981 15011
rect 18196 14980 18981 15008
rect 18196 14968 18202 14980
rect 18969 14977 18981 14980
rect 19015 14977 19027 15011
rect 18969 14971 19027 14977
rect 19245 15011 19303 15017
rect 19245 14977 19257 15011
rect 19291 15008 19303 15011
rect 19886 15008 19892 15020
rect 19291 14980 19892 15008
rect 19291 14977 19303 14980
rect 19245 14971 19303 14977
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 20717 15011 20775 15017
rect 20717 14977 20729 15011
rect 20763 15008 20775 15011
rect 20993 15011 21051 15017
rect 20993 15008 21005 15011
rect 20763 14980 21005 15008
rect 20763 14977 20775 14980
rect 20717 14971 20775 14977
rect 20993 14977 21005 14980
rect 21039 14977 21051 15011
rect 20993 14971 21051 14977
rect 22186 14968 22192 15020
rect 22244 15008 22250 15020
rect 22373 15011 22431 15017
rect 22373 15008 22385 15011
rect 22244 14980 22385 15008
rect 22244 14968 22250 14980
rect 22373 14977 22385 14980
rect 22419 15008 22431 15011
rect 22922 15008 22928 15020
rect 22419 14980 22928 15008
rect 22419 14977 22431 14980
rect 22373 14971 22431 14977
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 23569 15011 23627 15017
rect 23569 14977 23581 15011
rect 23615 14977 23627 15011
rect 23569 14971 23627 14977
rect 17972 14912 18276 14940
rect 17865 14903 17923 14909
rect 16632 14844 17080 14872
rect 16632 14832 16638 14844
rect 17052 14813 17080 14844
rect 17236 14844 17632 14872
rect 17236 14816 17264 14844
rect 17678 14832 17684 14884
rect 17736 14832 17742 14884
rect 16264 14776 16528 14804
rect 17037 14807 17095 14813
rect 16264 14764 16270 14776
rect 17037 14773 17049 14807
rect 17083 14773 17095 14807
rect 17037 14767 17095 14773
rect 17218 14764 17224 14816
rect 17276 14764 17282 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 17589 14807 17647 14813
rect 17589 14804 17601 14807
rect 17460 14776 17601 14804
rect 17460 14764 17466 14776
rect 17589 14773 17601 14776
rect 17635 14773 17647 14807
rect 17589 14767 17647 14773
rect 17954 14764 17960 14816
rect 18012 14764 18018 14816
rect 18046 14764 18052 14816
rect 18104 14804 18110 14816
rect 18141 14807 18199 14813
rect 18141 14804 18153 14807
rect 18104 14776 18153 14804
rect 18104 14764 18110 14776
rect 18141 14773 18153 14776
rect 18187 14773 18199 14807
rect 18248 14804 18276 14912
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 20346 14900 20352 14952
rect 20404 14900 20410 14952
rect 20622 14900 20628 14952
rect 20680 14940 20686 14952
rect 21913 14943 21971 14949
rect 21913 14940 21925 14943
rect 20680 14912 21925 14940
rect 20680 14900 20686 14912
rect 21913 14909 21925 14912
rect 21959 14940 21971 14943
rect 21959 14912 22416 14940
rect 21959 14909 21971 14912
rect 21913 14903 21971 14909
rect 18322 14832 18328 14884
rect 18380 14872 18386 14884
rect 19518 14872 19524 14884
rect 18380 14844 19524 14872
rect 18380 14832 18386 14844
rect 19518 14832 19524 14844
rect 19576 14832 19582 14884
rect 21821 14875 21879 14881
rect 21821 14872 21833 14875
rect 21468 14844 21833 14872
rect 21468 14816 21496 14844
rect 21821 14841 21833 14844
rect 21867 14841 21879 14875
rect 21821 14835 21879 14841
rect 20990 14804 20996 14816
rect 18248 14776 20996 14804
rect 18141 14767 18199 14773
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 21450 14764 21456 14816
rect 21508 14764 21514 14816
rect 21542 14764 21548 14816
rect 21600 14804 21606 14816
rect 21637 14807 21695 14813
rect 21637 14804 21649 14807
rect 21600 14776 21649 14804
rect 21600 14764 21606 14776
rect 21637 14773 21649 14776
rect 21683 14804 21695 14807
rect 22002 14804 22008 14816
rect 21683 14776 22008 14804
rect 21683 14773 21695 14776
rect 21637 14767 21695 14773
rect 22002 14764 22008 14776
rect 22060 14764 22066 14816
rect 22388 14804 22416 14912
rect 22462 14900 22468 14952
rect 22520 14900 22526 14952
rect 22554 14900 22560 14952
rect 22612 14900 22618 14952
rect 23584 14872 23612 14971
rect 24302 14900 24308 14952
rect 24360 14900 24366 14952
rect 22940 14844 23612 14872
rect 22830 14804 22836 14816
rect 22388 14776 22836 14804
rect 22830 14764 22836 14776
rect 22888 14764 22894 14816
rect 22940 14813 22968 14844
rect 22925 14807 22983 14813
rect 22925 14773 22937 14807
rect 22971 14773 22983 14807
rect 22925 14767 22983 14773
rect 23014 14764 23020 14816
rect 23072 14764 23078 14816
rect 23198 14764 23204 14816
rect 23256 14804 23262 14816
rect 24762 14804 24768 14816
rect 23256 14776 24768 14804
rect 23256 14764 23262 14776
rect 24762 14764 24768 14776
rect 24820 14764 24826 14816
rect 25608 14804 25636 15048
rect 29549 15045 29561 15079
rect 29595 15076 29607 15079
rect 30926 15076 30932 15088
rect 29595 15048 30932 15076
rect 29595 15045 29607 15048
rect 29549 15039 29607 15045
rect 30926 15036 30932 15048
rect 30984 15036 30990 15088
rect 26326 14968 26332 15020
rect 26384 14968 26390 15020
rect 27801 15011 27859 15017
rect 27801 14977 27813 15011
rect 27847 15008 27859 15011
rect 28074 15008 28080 15020
rect 27847 14980 28080 15008
rect 27847 14977 27859 14980
rect 27801 14971 27859 14977
rect 28074 14968 28080 14980
rect 28132 15008 28138 15020
rect 29181 15011 29239 15017
rect 29181 15008 29193 15011
rect 28132 14980 29193 15008
rect 28132 14968 28138 14980
rect 29181 14977 29193 14980
rect 29227 14977 29239 15011
rect 30469 15011 30527 15017
rect 30469 15008 30481 15011
rect 29181 14971 29239 14977
rect 29656 14980 30481 15008
rect 25685 14943 25743 14949
rect 25685 14909 25697 14943
rect 25731 14940 25743 14943
rect 25866 14940 25872 14952
rect 25731 14912 25872 14940
rect 25731 14909 25743 14912
rect 25685 14903 25743 14909
rect 25866 14900 25872 14912
rect 25924 14900 25930 14952
rect 26050 14900 26056 14952
rect 26108 14900 26114 14952
rect 28442 14900 28448 14952
rect 28500 14900 28506 14952
rect 28626 14900 28632 14952
rect 28684 14940 28690 14952
rect 29656 14940 29684 14980
rect 30469 14977 30481 14980
rect 30515 15008 30527 15011
rect 30515 14980 31708 15008
rect 30515 14977 30527 14980
rect 30469 14971 30527 14977
rect 28684 14912 29684 14940
rect 28684 14900 28690 14912
rect 29730 14900 29736 14952
rect 29788 14940 29794 14952
rect 29825 14943 29883 14949
rect 29825 14940 29837 14943
rect 29788 14912 29837 14940
rect 29788 14900 29794 14912
rect 29825 14909 29837 14912
rect 29871 14909 29883 14943
rect 29825 14903 29883 14909
rect 30653 14943 30711 14949
rect 30653 14909 30665 14943
rect 30699 14909 30711 14943
rect 30653 14903 30711 14909
rect 25777 14875 25835 14881
rect 25777 14841 25789 14875
rect 25823 14872 25835 14875
rect 28534 14872 28540 14884
rect 25823 14844 26818 14872
rect 27816 14844 28540 14872
rect 25823 14841 25835 14844
rect 25777 14835 25835 14841
rect 27816 14804 27844 14844
rect 28534 14832 28540 14844
rect 28592 14832 28598 14884
rect 30101 14875 30159 14881
rect 30101 14841 30113 14875
rect 30147 14841 30159 14875
rect 30668 14872 30696 14903
rect 30742 14900 30748 14952
rect 30800 14940 30806 14952
rect 31205 14943 31263 14949
rect 31205 14940 31217 14943
rect 30800 14912 31217 14940
rect 30800 14900 30806 14912
rect 31205 14909 31217 14912
rect 31251 14909 31263 14943
rect 31205 14903 31263 14909
rect 31680 14884 31708 14980
rect 30834 14872 30840 14884
rect 30668 14844 30840 14872
rect 30101 14835 30159 14841
rect 25608 14776 27844 14804
rect 27890 14764 27896 14816
rect 27948 14804 27954 14816
rect 28629 14807 28687 14813
rect 28629 14804 28641 14807
rect 27948 14776 28641 14804
rect 27948 14764 27954 14776
rect 28629 14773 28641 14776
rect 28675 14773 28687 14807
rect 28629 14767 28687 14773
rect 29454 14764 29460 14816
rect 29512 14804 29518 14816
rect 29733 14807 29791 14813
rect 29733 14804 29745 14807
rect 29512 14776 29745 14804
rect 29512 14764 29518 14776
rect 29733 14773 29745 14776
rect 29779 14773 29791 14807
rect 29733 14767 29791 14773
rect 29914 14764 29920 14816
rect 29972 14764 29978 14816
rect 30116 14804 30144 14835
rect 30834 14832 30840 14844
rect 30892 14832 30898 14884
rect 31662 14832 31668 14884
rect 31720 14832 31726 14884
rect 30650 14804 30656 14816
rect 30116 14776 30656 14804
rect 30650 14764 30656 14776
rect 30708 14764 30714 14816
rect 2760 14714 32200 14736
rect 2760 14662 6946 14714
rect 6998 14662 7010 14714
rect 7062 14662 7074 14714
rect 7126 14662 7138 14714
rect 7190 14662 7202 14714
rect 7254 14662 14306 14714
rect 14358 14662 14370 14714
rect 14422 14662 14434 14714
rect 14486 14662 14498 14714
rect 14550 14662 14562 14714
rect 14614 14662 21666 14714
rect 21718 14662 21730 14714
rect 21782 14662 21794 14714
rect 21846 14662 21858 14714
rect 21910 14662 21922 14714
rect 21974 14662 29026 14714
rect 29078 14662 29090 14714
rect 29142 14662 29154 14714
rect 29206 14662 29218 14714
rect 29270 14662 29282 14714
rect 29334 14662 32200 14714
rect 2760 14640 32200 14662
rect 6089 14603 6147 14609
rect 6089 14569 6101 14603
rect 6135 14600 6147 14603
rect 6135 14572 6500 14600
rect 6135 14569 6147 14572
rect 6089 14563 6147 14569
rect 5445 14535 5503 14541
rect 5445 14532 5457 14535
rect 4554 14504 5457 14532
rect 5445 14501 5457 14504
rect 5491 14501 5503 14535
rect 6178 14532 6184 14544
rect 5445 14495 5503 14501
rect 5552 14504 6184 14532
rect 5552 14473 5580 14504
rect 6178 14492 6184 14504
rect 6236 14492 6242 14544
rect 6472 14473 6500 14572
rect 6546 14560 6552 14612
rect 6604 14560 6610 14612
rect 6825 14603 6883 14609
rect 6825 14569 6837 14603
rect 6871 14600 6883 14603
rect 7650 14600 7656 14612
rect 6871 14572 7656 14600
rect 6871 14569 6883 14572
rect 6825 14563 6883 14569
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 8018 14560 8024 14612
rect 8076 14600 8082 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 8076 14572 8125 14600
rect 8076 14560 8082 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 8478 14560 8484 14612
rect 8536 14560 8542 14612
rect 8938 14560 8944 14612
rect 8996 14560 9002 14612
rect 9858 14560 9864 14612
rect 9916 14600 9922 14612
rect 10318 14600 10324 14612
rect 9916 14572 10324 14600
rect 9916 14560 9922 14572
rect 10318 14560 10324 14572
rect 10376 14600 10382 14612
rect 10689 14603 10747 14609
rect 10689 14600 10701 14603
rect 10376 14572 10701 14600
rect 10376 14560 10382 14572
rect 10689 14569 10701 14572
rect 10735 14569 10747 14603
rect 10689 14563 10747 14569
rect 11146 14560 11152 14612
rect 11204 14600 11210 14612
rect 11701 14603 11759 14609
rect 11701 14600 11713 14603
rect 11204 14572 11713 14600
rect 11204 14560 11210 14572
rect 11701 14569 11713 14572
rect 11747 14569 11759 14603
rect 12894 14600 12900 14612
rect 11701 14563 11759 14569
rect 11900 14572 12900 14600
rect 6564 14473 6592 14560
rect 7374 14532 7380 14544
rect 6656 14504 7380 14532
rect 6656 14473 6684 14504
rect 7374 14492 7380 14504
rect 7432 14532 7438 14544
rect 8496 14532 8524 14560
rect 7432 14504 8524 14532
rect 10520 14504 11284 14532
rect 7432 14492 7438 14504
rect 5537 14467 5595 14473
rect 5537 14433 5549 14467
rect 5583 14433 5595 14467
rect 5537 14427 5595 14433
rect 6273 14467 6331 14473
rect 6273 14433 6285 14467
rect 6319 14433 6331 14467
rect 6273 14427 6331 14433
rect 6457 14467 6515 14473
rect 6457 14433 6469 14467
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 6641 14467 6699 14473
rect 6641 14433 6653 14467
rect 6687 14433 6699 14467
rect 6641 14427 6699 14433
rect 4430 14356 4436 14408
rect 4488 14396 4494 14408
rect 4985 14399 5043 14405
rect 4985 14396 4997 14399
rect 4488 14368 4997 14396
rect 4488 14356 4494 14368
rect 4985 14365 4997 14368
rect 5031 14365 5043 14399
rect 4985 14359 5043 14365
rect 5261 14399 5319 14405
rect 5261 14365 5273 14399
rect 5307 14396 5319 14399
rect 5442 14396 5448 14408
rect 5307 14368 5448 14396
rect 5307 14365 5319 14368
rect 5261 14359 5319 14365
rect 5442 14356 5448 14368
rect 5500 14356 5506 14408
rect 6288 14328 6316 14427
rect 6472 14396 6500 14427
rect 8018 14424 8024 14476
rect 8076 14424 8082 14476
rect 8849 14467 8907 14473
rect 8849 14433 8861 14467
rect 8895 14464 8907 14467
rect 9309 14467 9367 14473
rect 9309 14464 9321 14467
rect 8895 14436 9321 14464
rect 8895 14433 8907 14436
rect 8849 14427 8907 14433
rect 9309 14433 9321 14436
rect 9355 14433 9367 14467
rect 9309 14427 9367 14433
rect 6472 14368 7880 14396
rect 7742 14328 7748 14340
rect 6288 14300 7748 14328
rect 7742 14288 7748 14300
rect 7800 14288 7806 14340
rect 7852 14328 7880 14368
rect 9030 14356 9036 14408
rect 9088 14356 9094 14408
rect 9122 14356 9128 14408
rect 9180 14396 9186 14408
rect 9861 14399 9919 14405
rect 9861 14396 9873 14399
rect 9180 14368 9873 14396
rect 9180 14356 9186 14368
rect 9861 14365 9873 14368
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 9674 14328 9680 14340
rect 7852 14300 9680 14328
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 3513 14263 3571 14269
rect 3513 14229 3525 14263
rect 3559 14260 3571 14263
rect 4246 14260 4252 14272
rect 3559 14232 4252 14260
rect 3559 14229 3571 14232
rect 3513 14223 3571 14229
rect 4246 14220 4252 14232
rect 4304 14220 4310 14272
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 10226 14220 10232 14272
rect 10284 14260 10290 14272
rect 10520 14269 10548 14504
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14464 11023 14467
rect 11146 14464 11152 14476
rect 11011 14436 11152 14464
rect 11011 14433 11023 14436
rect 10965 14427 11023 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 11256 14473 11284 14504
rect 11330 14492 11336 14544
rect 11388 14532 11394 14544
rect 11900 14532 11928 14572
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13262 14560 13268 14612
rect 13320 14560 13326 14612
rect 13354 14560 13360 14612
rect 13412 14600 13418 14612
rect 13998 14600 14004 14612
rect 13412 14572 14004 14600
rect 13412 14560 13418 14572
rect 13998 14560 14004 14572
rect 14056 14560 14062 14612
rect 14642 14560 14648 14612
rect 14700 14560 14706 14612
rect 15381 14603 15439 14609
rect 15381 14569 15393 14603
rect 15427 14600 15439 14603
rect 17034 14600 17040 14612
rect 15427 14572 17040 14600
rect 15427 14569 15439 14572
rect 15381 14563 15439 14569
rect 17034 14560 17040 14572
rect 17092 14560 17098 14612
rect 17405 14603 17463 14609
rect 17405 14569 17417 14603
rect 17451 14600 17463 14603
rect 17451 14572 17632 14600
rect 17451 14569 17463 14572
rect 17405 14563 17463 14569
rect 13280 14532 13308 14560
rect 11388 14504 11928 14532
rect 11388 14492 11394 14504
rect 11241 14467 11299 14473
rect 11241 14433 11253 14467
rect 11287 14433 11299 14467
rect 11241 14427 11299 14433
rect 11422 14424 11428 14476
rect 11480 14464 11486 14476
rect 11900 14473 11928 14504
rect 13188 14504 13308 14532
rect 11517 14467 11575 14473
rect 11517 14464 11529 14467
rect 11480 14436 11529 14464
rect 11480 14424 11486 14436
rect 11517 14433 11529 14436
rect 11563 14433 11575 14467
rect 11517 14427 11575 14433
rect 11607 14467 11665 14473
rect 11607 14433 11619 14467
rect 11653 14464 11665 14467
rect 11885 14467 11943 14473
rect 11653 14436 11836 14464
rect 11653 14433 11665 14436
rect 11607 14427 11665 14433
rect 11808 14408 11836 14436
rect 11885 14433 11897 14467
rect 11931 14433 11943 14467
rect 11885 14427 11943 14433
rect 11974 14424 11980 14476
rect 12032 14424 12038 14476
rect 12345 14467 12403 14473
rect 12345 14464 12357 14467
rect 12084 14436 12357 14464
rect 10870 14356 10876 14408
rect 10928 14356 10934 14408
rect 11790 14356 11796 14408
rect 11848 14396 11854 14408
rect 12084 14405 12112 14436
rect 12345 14433 12357 14436
rect 12391 14464 12403 14467
rect 12618 14464 12624 14476
rect 12391 14436 12624 14464
rect 12391 14433 12403 14436
rect 12345 14427 12403 14433
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 12713 14467 12771 14473
rect 12713 14433 12725 14467
rect 12759 14464 12771 14467
rect 13078 14464 13084 14476
rect 12759 14436 13084 14464
rect 12759 14433 12771 14436
rect 12713 14427 12771 14433
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13188 14473 13216 14504
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14433 13231 14467
rect 13173 14427 13231 14433
rect 13265 14467 13323 14473
rect 13265 14433 13277 14467
rect 13311 14464 13323 14467
rect 13372 14464 13400 14560
rect 14660 14532 14688 14560
rect 13832 14504 14780 14532
rect 13311 14436 13400 14464
rect 13311 14433 13323 14436
rect 13265 14427 13323 14433
rect 13446 14424 13452 14476
rect 13504 14424 13510 14476
rect 12069 14399 12127 14405
rect 12069 14396 12081 14399
rect 11848 14368 12081 14396
rect 11848 14356 11854 14368
rect 12069 14365 12081 14368
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12636 14396 12664 14424
rect 13832 14396 13860 14504
rect 14642 14424 14648 14476
rect 14700 14424 14706 14476
rect 14752 14473 14780 14504
rect 15028 14504 15332 14532
rect 14737 14467 14795 14473
rect 14737 14433 14749 14467
rect 14783 14433 14795 14467
rect 14737 14427 14795 14433
rect 12636 14368 13860 14396
rect 13909 14399 13967 14405
rect 12161 14359 12219 14365
rect 13909 14365 13921 14399
rect 13955 14396 13967 14399
rect 14090 14396 14096 14408
rect 13955 14368 14096 14396
rect 13955 14365 13967 14368
rect 13909 14359 13967 14365
rect 10888 14328 10916 14356
rect 12176 14328 12204 14359
rect 14090 14356 14096 14368
rect 14148 14396 14154 14408
rect 14550 14396 14556 14408
rect 14148 14368 14556 14396
rect 14148 14356 14154 14368
rect 14550 14356 14556 14368
rect 14608 14396 14614 14408
rect 15028 14405 15056 14504
rect 15197 14467 15255 14473
rect 15197 14464 15209 14467
rect 15120 14436 15209 14464
rect 15013 14399 15071 14405
rect 15013 14396 15025 14399
rect 14608 14368 15025 14396
rect 14608 14356 14614 14368
rect 15013 14365 15025 14368
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15120 14328 15148 14436
rect 15197 14433 15209 14436
rect 15243 14433 15255 14467
rect 15197 14427 15255 14433
rect 15304 14396 15332 14504
rect 15470 14492 15476 14544
rect 15528 14532 15534 14544
rect 15838 14532 15844 14544
rect 15528 14504 15844 14532
rect 15528 14492 15534 14504
rect 15838 14492 15844 14504
rect 15896 14532 15902 14544
rect 17604 14532 17632 14572
rect 17678 14560 17684 14612
rect 17736 14600 17742 14612
rect 18141 14603 18199 14609
rect 18141 14600 18153 14603
rect 17736 14572 18153 14600
rect 17736 14560 17742 14572
rect 18141 14569 18153 14572
rect 18187 14569 18199 14603
rect 18141 14563 18199 14569
rect 18690 14560 18696 14612
rect 18748 14560 18754 14612
rect 20346 14560 20352 14612
rect 20404 14600 20410 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 20404 14572 20453 14600
rect 20404 14560 20410 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 23014 14600 23020 14612
rect 20441 14563 20499 14569
rect 21652 14572 23020 14600
rect 18708 14532 18736 14560
rect 15896 14504 17448 14532
rect 17604 14504 18736 14532
rect 20165 14535 20223 14541
rect 15896 14492 15902 14504
rect 15562 14424 15568 14476
rect 15620 14464 15626 14476
rect 15657 14467 15715 14473
rect 15657 14464 15669 14467
rect 15620 14436 15669 14464
rect 15620 14424 15626 14436
rect 15657 14433 15669 14436
rect 15703 14433 15715 14467
rect 15657 14427 15715 14433
rect 16666 14424 16672 14476
rect 16724 14464 16730 14476
rect 16853 14467 16911 14473
rect 16853 14464 16865 14467
rect 16724 14436 16865 14464
rect 16724 14424 16730 14436
rect 16853 14433 16865 14436
rect 16899 14433 16911 14467
rect 16853 14427 16911 14433
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 17037 14467 17095 14473
rect 17037 14464 17049 14467
rect 17000 14436 17049 14464
rect 17000 14424 17006 14436
rect 17037 14433 17049 14436
rect 17083 14433 17095 14467
rect 17037 14427 17095 14433
rect 17129 14467 17187 14473
rect 17129 14433 17141 14467
rect 17175 14433 17187 14467
rect 17129 14427 17187 14433
rect 17221 14467 17279 14473
rect 17221 14433 17233 14467
rect 17267 14464 17279 14467
rect 17310 14464 17316 14476
rect 17267 14436 17316 14464
rect 17267 14433 17279 14436
rect 17221 14427 17279 14433
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15304 14368 15853 14396
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15930 14356 15936 14408
rect 15988 14356 15994 14408
rect 10888 14300 12204 14328
rect 12268 14300 15148 14328
rect 15473 14331 15531 14337
rect 10505 14263 10563 14269
rect 10505 14260 10517 14263
rect 10284 14232 10517 14260
rect 10284 14220 10290 14232
rect 10505 14229 10517 14232
rect 10551 14229 10563 14263
rect 10505 14223 10563 14229
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 10873 14263 10931 14269
rect 10873 14260 10885 14263
rect 10744 14232 10885 14260
rect 10744 14220 10750 14232
rect 10873 14229 10885 14232
rect 10919 14229 10931 14263
rect 10873 14223 10931 14229
rect 11606 14220 11612 14272
rect 11664 14220 11670 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 12268 14260 12296 14300
rect 15473 14297 15485 14331
rect 15519 14297 15531 14331
rect 17144 14328 17172 14427
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17420 14464 17448 14504
rect 20165 14501 20177 14535
rect 20211 14532 20223 14535
rect 20898 14532 20904 14544
rect 20211 14504 20904 14532
rect 20211 14501 20223 14504
rect 20165 14495 20223 14501
rect 20898 14492 20904 14504
rect 20956 14492 20962 14544
rect 20990 14492 20996 14544
rect 21048 14492 21054 14544
rect 21652 14541 21680 14572
rect 23014 14560 23020 14572
rect 23072 14560 23078 14612
rect 23566 14560 23572 14612
rect 23624 14560 23630 14612
rect 25866 14560 25872 14612
rect 25924 14600 25930 14612
rect 25924 14572 27108 14600
rect 25924 14560 25930 14572
rect 21637 14535 21695 14541
rect 21637 14501 21649 14535
rect 21683 14501 21695 14535
rect 23845 14535 23903 14541
rect 23845 14532 23857 14535
rect 22862 14504 23857 14532
rect 21637 14495 21695 14501
rect 23845 14501 23857 14504
rect 23891 14501 23903 14535
rect 26050 14532 26056 14544
rect 23845 14495 23903 14501
rect 25516 14504 26056 14532
rect 18322 14464 18328 14476
rect 17420 14436 18328 14464
rect 18322 14424 18328 14436
rect 18380 14424 18386 14476
rect 18601 14467 18659 14473
rect 18601 14433 18613 14467
rect 18647 14464 18659 14467
rect 19150 14464 19156 14476
rect 18647 14436 19156 14464
rect 18647 14433 18659 14436
rect 18601 14427 18659 14433
rect 19150 14424 19156 14436
rect 19208 14464 19214 14476
rect 20533 14467 20591 14473
rect 20533 14464 20545 14467
rect 19208 14436 20545 14464
rect 19208 14424 19214 14436
rect 20533 14433 20545 14436
rect 20579 14464 20591 14467
rect 20622 14464 20628 14476
rect 20579 14436 20628 14464
rect 20579 14433 20591 14436
rect 20533 14427 20591 14433
rect 20622 14424 20628 14436
rect 20680 14424 20686 14476
rect 20717 14467 20775 14473
rect 20717 14433 20729 14467
rect 20763 14433 20775 14467
rect 21177 14467 21235 14473
rect 21177 14464 21189 14467
rect 20717 14427 20775 14433
rect 20824 14436 21189 14464
rect 17494 14356 17500 14408
rect 17552 14356 17558 14408
rect 19426 14356 19432 14408
rect 19484 14356 19490 14408
rect 18874 14328 18880 14340
rect 17144 14300 18880 14328
rect 15473 14291 15531 14297
rect 11940 14232 12296 14260
rect 13633 14263 13691 14269
rect 11940 14220 11946 14232
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 14090 14260 14096 14272
rect 13679 14232 14096 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 14090 14220 14096 14232
rect 14148 14220 14154 14272
rect 14826 14220 14832 14272
rect 14884 14220 14890 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15488 14260 15516 14291
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 20732 14328 20760 14427
rect 20824 14408 20852 14436
rect 21177 14433 21189 14436
rect 21223 14433 21235 14467
rect 21177 14427 21235 14433
rect 22922 14424 22928 14476
rect 22980 14464 22986 14476
rect 23658 14464 23664 14476
rect 22980 14436 23664 14464
rect 22980 14424 22986 14436
rect 23658 14424 23664 14436
rect 23716 14464 23722 14476
rect 23937 14467 23995 14473
rect 23937 14464 23949 14467
rect 23716 14436 23949 14464
rect 23716 14424 23722 14436
rect 23937 14433 23949 14436
rect 23983 14433 23995 14467
rect 23937 14427 23995 14433
rect 24026 14424 24032 14476
rect 24084 14424 24090 14476
rect 25516 14473 25544 14504
rect 26050 14492 26056 14504
rect 26108 14492 26114 14544
rect 27080 14532 27108 14572
rect 27154 14560 27160 14612
rect 27212 14600 27218 14612
rect 27617 14603 27675 14609
rect 27617 14600 27629 14603
rect 27212 14572 27629 14600
rect 27212 14560 27218 14572
rect 27617 14569 27629 14572
rect 27663 14569 27675 14603
rect 27617 14563 27675 14569
rect 27798 14560 27804 14612
rect 27856 14600 27862 14612
rect 28077 14603 28135 14609
rect 27856 14572 27936 14600
rect 27856 14560 27862 14572
rect 27908 14532 27936 14572
rect 28077 14569 28089 14603
rect 28123 14600 28135 14603
rect 28442 14600 28448 14612
rect 28123 14572 28448 14600
rect 28123 14569 28135 14572
rect 28077 14563 28135 14569
rect 28442 14560 28448 14572
rect 28500 14560 28506 14612
rect 28534 14560 28540 14612
rect 28592 14600 28598 14612
rect 31665 14603 31723 14609
rect 31665 14600 31677 14603
rect 28592 14572 31677 14600
rect 28592 14560 28598 14572
rect 31665 14569 31677 14572
rect 31711 14569 31723 14603
rect 31665 14563 31723 14569
rect 28810 14541 28816 14544
rect 28261 14535 28319 14541
rect 28261 14532 28273 14535
rect 27080 14504 27844 14532
rect 27908 14504 28273 14532
rect 25501 14467 25559 14473
rect 25501 14433 25513 14467
rect 25547 14433 25559 14467
rect 27522 14464 27528 14476
rect 26910 14436 27528 14464
rect 25501 14427 25559 14433
rect 27522 14424 27528 14436
rect 27580 14424 27586 14476
rect 27706 14424 27712 14476
rect 27764 14424 27770 14476
rect 27816 14464 27844 14504
rect 28261 14501 28273 14504
rect 28307 14501 28319 14535
rect 28261 14495 28319 14501
rect 28797 14535 28816 14541
rect 28797 14501 28809 14535
rect 28797 14495 28816 14501
rect 28810 14492 28816 14495
rect 28868 14492 28874 14544
rect 28997 14535 29055 14541
rect 28997 14501 29009 14535
rect 29043 14501 29055 14535
rect 28997 14495 29055 14501
rect 28353 14467 28411 14473
rect 28353 14464 28365 14467
rect 27816 14436 28365 14464
rect 28353 14433 28365 14436
rect 28399 14464 28411 14467
rect 28626 14464 28632 14476
rect 28399 14436 28632 14464
rect 28399 14433 28411 14436
rect 28353 14427 28411 14433
rect 28626 14424 28632 14436
rect 28684 14424 28690 14476
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 21358 14356 21364 14408
rect 21416 14356 21422 14408
rect 25406 14396 25412 14408
rect 21468 14368 25412 14396
rect 20898 14328 20904 14340
rect 20732 14300 20904 14328
rect 20898 14288 20904 14300
rect 20956 14288 20962 14340
rect 21468 14328 21496 14368
rect 25406 14356 25412 14368
rect 25464 14356 25470 14408
rect 25774 14356 25780 14408
rect 25832 14356 25838 14408
rect 27433 14399 27491 14405
rect 27433 14365 27445 14399
rect 27479 14396 27491 14399
rect 27614 14396 27620 14408
rect 27479 14368 27620 14396
rect 27479 14365 27491 14368
rect 27433 14359 27491 14365
rect 27614 14356 27620 14368
rect 27672 14396 27678 14408
rect 27982 14396 27988 14408
rect 27672 14368 27988 14396
rect 27672 14356 27678 14368
rect 27982 14356 27988 14368
rect 28040 14396 28046 14408
rect 29012 14396 29040 14495
rect 30282 14492 30288 14544
rect 30340 14532 30346 14544
rect 30340 14504 30880 14532
rect 30340 14492 30346 14504
rect 30852 14476 30880 14504
rect 30650 14424 30656 14476
rect 30708 14424 30714 14476
rect 30834 14424 30840 14476
rect 30892 14424 30898 14476
rect 31849 14467 31907 14473
rect 31849 14433 31861 14467
rect 31895 14464 31907 14467
rect 31895 14436 33180 14464
rect 31895 14433 31907 14436
rect 31849 14427 31907 14433
rect 33152 14408 33180 14436
rect 28040 14368 29040 14396
rect 28040 14356 28046 14368
rect 29270 14356 29276 14408
rect 29328 14356 29334 14408
rect 29914 14356 29920 14408
rect 29972 14396 29978 14408
rect 31018 14396 31024 14408
rect 29972 14368 31024 14396
rect 29972 14356 29978 14368
rect 31018 14356 31024 14368
rect 31076 14356 31082 14408
rect 31294 14356 31300 14408
rect 31352 14356 31358 14408
rect 33134 14356 33140 14408
rect 33192 14356 33198 14408
rect 21008 14300 21496 14328
rect 23109 14331 23167 14337
rect 14976 14232 15516 14260
rect 14976 14220 14982 14232
rect 16574 14220 16580 14272
rect 16632 14220 16638 14272
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 18598 14260 18604 14272
rect 17460 14232 18604 14260
rect 17460 14220 17466 14232
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 18690 14220 18696 14272
rect 18748 14220 18754 14272
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 21008 14260 21036 14300
rect 23109 14297 23121 14331
rect 23155 14328 23167 14331
rect 24302 14328 24308 14340
rect 23155 14300 24308 14328
rect 23155 14297 23167 14300
rect 23109 14291 23167 14297
rect 24302 14288 24308 14300
rect 24360 14288 24366 14340
rect 27249 14331 27307 14337
rect 27249 14297 27261 14331
rect 27295 14328 27307 14331
rect 27798 14328 27804 14340
rect 27295 14300 27804 14328
rect 27295 14297 27307 14300
rect 27249 14291 27307 14297
rect 27798 14288 27804 14300
rect 27856 14328 27862 14340
rect 27856 14300 28856 14328
rect 27856 14288 27862 14300
rect 20128 14232 21036 14260
rect 20128 14220 20134 14232
rect 22646 14220 22652 14272
rect 22704 14260 22710 14272
rect 24213 14263 24271 14269
rect 24213 14260 24225 14263
rect 22704 14232 24225 14260
rect 22704 14220 22710 14232
rect 24213 14229 24225 14232
rect 24259 14229 24271 14263
rect 24213 14223 24271 14229
rect 24762 14220 24768 14272
rect 24820 14260 24826 14272
rect 25409 14263 25467 14269
rect 25409 14260 25421 14263
rect 24820 14232 25421 14260
rect 24820 14220 24826 14232
rect 25409 14229 25421 14232
rect 25455 14260 25467 14263
rect 26142 14260 26148 14272
rect 25455 14232 26148 14260
rect 25455 14229 25467 14232
rect 25409 14223 25467 14229
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 27338 14220 27344 14272
rect 27396 14260 27402 14272
rect 28828 14269 28856 14300
rect 28902 14288 28908 14340
rect 28960 14328 28966 14340
rect 30469 14331 30527 14337
rect 30469 14328 30481 14331
rect 28960 14300 30481 14328
rect 28960 14288 28966 14300
rect 30469 14297 30481 14300
rect 30515 14297 30527 14331
rect 30469 14291 30527 14297
rect 28629 14263 28687 14269
rect 28629 14260 28641 14263
rect 27396 14232 28641 14260
rect 27396 14220 27402 14232
rect 28629 14229 28641 14232
rect 28675 14229 28687 14263
rect 28629 14223 28687 14229
rect 28813 14263 28871 14269
rect 28813 14229 28825 14263
rect 28859 14229 28871 14263
rect 28813 14223 28871 14229
rect 29638 14220 29644 14272
rect 29696 14260 29702 14272
rect 29917 14263 29975 14269
rect 29917 14260 29929 14263
rect 29696 14232 29929 14260
rect 29696 14220 29702 14232
rect 29917 14229 29929 14232
rect 29963 14229 29975 14263
rect 29917 14223 29975 14229
rect 30742 14220 30748 14272
rect 30800 14220 30806 14272
rect 2760 14170 32200 14192
rect 2760 14118 6286 14170
rect 6338 14118 6350 14170
rect 6402 14118 6414 14170
rect 6466 14118 6478 14170
rect 6530 14118 6542 14170
rect 6594 14118 13646 14170
rect 13698 14118 13710 14170
rect 13762 14118 13774 14170
rect 13826 14118 13838 14170
rect 13890 14118 13902 14170
rect 13954 14118 21006 14170
rect 21058 14118 21070 14170
rect 21122 14118 21134 14170
rect 21186 14118 21198 14170
rect 21250 14118 21262 14170
rect 21314 14118 28366 14170
rect 28418 14118 28430 14170
rect 28482 14118 28494 14170
rect 28546 14118 28558 14170
rect 28610 14118 28622 14170
rect 28674 14118 32200 14170
rect 2760 14096 32200 14118
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 6273 14059 6331 14065
rect 6273 14056 6285 14059
rect 5684 14028 6285 14056
rect 5684 14016 5690 14028
rect 6273 14025 6285 14028
rect 6319 14056 6331 14059
rect 6638 14056 6644 14068
rect 6319 14028 6644 14056
rect 6319 14025 6331 14028
rect 6273 14019 6331 14025
rect 6638 14016 6644 14028
rect 6696 14016 6702 14068
rect 6904 14059 6962 14065
rect 6904 14025 6916 14059
rect 6950 14056 6962 14059
rect 8478 14056 8484 14068
rect 6950 14028 8484 14056
rect 6950 14025 6962 14028
rect 6904 14019 6962 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 9122 14016 9128 14068
rect 9180 14016 9186 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11149 14059 11207 14065
rect 11149 14056 11161 14059
rect 11112 14028 11161 14056
rect 11112 14016 11118 14028
rect 11149 14025 11161 14028
rect 11195 14025 11207 14059
rect 11149 14019 11207 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12492 14028 12940 14056
rect 12492 14016 12498 14028
rect 8389 13991 8447 13997
rect 8389 13957 8401 13991
rect 8435 13988 8447 13991
rect 9140 13988 9168 14016
rect 8435 13960 9168 13988
rect 10689 13991 10747 13997
rect 8435 13957 8447 13960
rect 8389 13951 8447 13957
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 11330 13988 11336 14000
rect 10735 13960 11336 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 11330 13948 11336 13960
rect 11388 13948 11394 14000
rect 12912 13988 12940 14028
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 13136 14028 13369 14056
rect 13136 14016 13142 14028
rect 13357 14025 13369 14028
rect 13403 14025 13415 14059
rect 13357 14019 13415 14025
rect 14185 14059 14243 14065
rect 14185 14025 14197 14059
rect 14231 14056 14243 14059
rect 14642 14056 14648 14068
rect 14231 14028 14648 14056
rect 14231 14025 14243 14028
rect 14185 14019 14243 14025
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 14737 14059 14795 14065
rect 14737 14025 14749 14059
rect 14783 14056 14795 14059
rect 14826 14056 14832 14068
rect 14783 14028 14832 14056
rect 14783 14025 14795 14028
rect 14737 14019 14795 14025
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 15102 14016 15108 14068
rect 15160 14056 15166 14068
rect 15197 14059 15255 14065
rect 15197 14056 15209 14059
rect 15160 14028 15209 14056
rect 15160 14016 15166 14028
rect 15197 14025 15209 14028
rect 15243 14025 15255 14059
rect 15197 14019 15255 14025
rect 17494 14016 17500 14068
rect 17552 14016 17558 14068
rect 18138 14056 18144 14068
rect 17696 14028 18144 14056
rect 13449 13991 13507 13997
rect 13449 13988 13461 13991
rect 12912 13960 13461 13988
rect 13449 13957 13461 13960
rect 13495 13957 13507 13991
rect 13449 13951 13507 13957
rect 14274 13948 14280 14000
rect 14332 13988 14338 14000
rect 15013 13991 15071 13997
rect 15013 13988 15025 13991
rect 14332 13960 15025 13988
rect 14332 13948 14338 13960
rect 15013 13957 15025 13960
rect 15059 13957 15071 13991
rect 15013 13951 15071 13957
rect 1302 13880 1308 13932
rect 1360 13920 1366 13932
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 1360 13892 3249 13920
rect 1360 13880 1366 13892
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 3237 13883 3295 13889
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 6641 13923 6699 13929
rect 6641 13920 6653 13923
rect 5500 13892 6653 13920
rect 5500 13880 5506 13892
rect 6641 13889 6653 13892
rect 6687 13920 6699 13923
rect 7282 13920 7288 13932
rect 6687 13892 7288 13920
rect 6687 13889 6699 13892
rect 6641 13883 6699 13889
rect 7282 13880 7288 13892
rect 7340 13920 7346 13932
rect 8202 13920 8208 13932
rect 7340 13892 8208 13920
rect 7340 13880 7346 13892
rect 8202 13880 8208 13892
rect 8260 13920 8266 13932
rect 8849 13923 8907 13929
rect 8849 13920 8861 13923
rect 8260 13892 8861 13920
rect 8260 13880 8266 13892
rect 8849 13889 8861 13892
rect 8895 13920 8907 13923
rect 10042 13920 10048 13932
rect 8895 13892 10048 13920
rect 8895 13889 8907 13892
rect 8849 13883 8907 13889
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10152 13892 10732 13920
rect 4246 13812 4252 13864
rect 4304 13812 4310 13864
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13852 9643 13855
rect 9861 13855 9919 13861
rect 9631 13824 9812 13852
rect 9631 13821 9643 13824
rect 9585 13815 9643 13821
rect 7650 13744 7656 13796
rect 7708 13744 7714 13796
rect 9784 13784 9812 13824
rect 9861 13821 9873 13855
rect 9907 13852 9919 13855
rect 10152 13852 10180 13892
rect 9907 13824 10180 13852
rect 10321 13855 10379 13861
rect 9907 13821 9919 13824
rect 9861 13815 9919 13821
rect 10321 13821 10333 13855
rect 10367 13852 10379 13855
rect 10594 13852 10600 13864
rect 10367 13824 10600 13852
rect 10367 13821 10379 13824
rect 10321 13815 10379 13821
rect 10594 13812 10600 13824
rect 10652 13812 10658 13864
rect 10704 13852 10732 13892
rect 10870 13880 10876 13932
rect 10928 13880 10934 13932
rect 11609 13923 11667 13929
rect 11609 13920 11621 13923
rect 11164 13892 11621 13920
rect 11164 13864 11192 13892
rect 11609 13889 11621 13892
rect 11655 13920 11667 13923
rect 14182 13920 14188 13932
rect 11655 13892 14188 13920
rect 11655 13889 11667 13892
rect 11609 13883 11667 13889
rect 14182 13880 14188 13892
rect 14240 13920 14246 13932
rect 15749 13923 15807 13929
rect 15749 13920 15761 13923
rect 14240 13892 15761 13920
rect 14240 13880 14246 13892
rect 15749 13889 15761 13892
rect 15795 13889 15807 13923
rect 15749 13883 15807 13889
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16574 13920 16580 13932
rect 16071 13892 16580 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16574 13880 16580 13892
rect 16632 13880 16638 13932
rect 17696 13929 17724 14028
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 18598 14016 18604 14068
rect 18656 14056 18662 14068
rect 18656 14028 19380 14056
rect 18656 14016 18662 14028
rect 19352 13988 19380 14028
rect 19426 14016 19432 14068
rect 19484 14016 19490 14068
rect 20806 14056 20812 14068
rect 20456 14028 20812 14056
rect 20456 13988 20484 14028
rect 20806 14016 20812 14028
rect 20864 14056 20870 14068
rect 25225 14059 25283 14065
rect 20864 14028 22876 14056
rect 20864 14016 20870 14028
rect 19352 13960 20484 13988
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 17957 13923 18015 13929
rect 17957 13889 17969 13923
rect 18003 13920 18015 13923
rect 18046 13920 18052 13932
rect 18003 13892 18052 13920
rect 18003 13889 18015 13892
rect 17957 13883 18015 13889
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 11054 13852 11060 13864
rect 10704 13824 11060 13852
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11146 13812 11152 13864
rect 11204 13812 11210 13864
rect 11238 13812 11244 13864
rect 11296 13812 11302 13864
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 14001 13855 14059 13861
rect 14001 13852 14013 13855
rect 13596 13824 14013 13852
rect 13596 13812 13602 13824
rect 14001 13821 14013 13824
rect 14047 13821 14059 13855
rect 14001 13815 14059 13821
rect 14274 13812 14280 13864
rect 14332 13861 14338 13864
rect 14332 13855 14368 13861
rect 14356 13821 14368 13855
rect 14332 13815 14368 13821
rect 14829 13855 14887 13861
rect 14829 13821 14841 13855
rect 14875 13852 14887 13855
rect 14918 13852 14924 13864
rect 14875 13824 14924 13852
rect 14875 13821 14887 13824
rect 14829 13815 14887 13821
rect 14332 13812 14338 13815
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13852 15623 13855
rect 15654 13852 15660 13864
rect 15611 13824 15660 13852
rect 15611 13821 15623 13824
rect 15565 13815 15623 13821
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 20070 13812 20076 13864
rect 20128 13812 20134 13864
rect 20456 13861 20484 13960
rect 20625 13991 20683 13997
rect 20625 13957 20637 13991
rect 20671 13988 20683 13991
rect 20671 13960 22784 13988
rect 20671 13957 20683 13960
rect 20625 13951 20683 13957
rect 20898 13920 20904 13932
rect 20732 13892 20904 13920
rect 20732 13861 20760 13892
rect 20898 13880 20904 13892
rect 20956 13920 20962 13932
rect 22278 13920 22284 13932
rect 20956 13892 22284 13920
rect 20956 13880 20962 13892
rect 22278 13880 22284 13892
rect 22336 13920 22342 13932
rect 22646 13920 22652 13932
rect 22336 13892 22652 13920
rect 22336 13880 22342 13892
rect 22646 13880 22652 13892
rect 22704 13880 22710 13932
rect 20441 13855 20499 13861
rect 20441 13821 20453 13855
rect 20487 13821 20499 13855
rect 20441 13815 20499 13821
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13821 20775 13855
rect 20717 13815 20775 13821
rect 20806 13812 20812 13864
rect 20864 13852 20870 13864
rect 21453 13855 21511 13861
rect 21453 13852 21465 13855
rect 20864 13824 21465 13852
rect 20864 13812 20870 13824
rect 21453 13821 21465 13824
rect 21499 13821 21511 13855
rect 21453 13815 21511 13821
rect 22094 13812 22100 13864
rect 22152 13852 22158 13864
rect 22189 13855 22247 13861
rect 22189 13852 22201 13855
rect 22152 13824 22201 13852
rect 22152 13812 22158 13824
rect 22189 13821 22201 13824
rect 22235 13821 22247 13855
rect 22189 13815 22247 13821
rect 10410 13784 10416 13796
rect 9784 13756 10416 13784
rect 10410 13744 10416 13756
rect 10468 13744 10474 13796
rect 11790 13784 11796 13796
rect 11072 13756 11796 13784
rect 9766 13676 9772 13728
rect 9824 13676 9830 13728
rect 11072 13725 11100 13756
rect 11790 13744 11796 13756
rect 11848 13744 11854 13796
rect 11882 13744 11888 13796
rect 11940 13744 11946 13796
rect 12618 13744 12624 13796
rect 12676 13744 12682 13796
rect 14090 13744 14096 13796
rect 14148 13784 14154 13796
rect 14148 13756 14412 13784
rect 14148 13744 14154 13756
rect 11057 13719 11115 13725
rect 11057 13685 11069 13719
rect 11103 13685 11115 13719
rect 11057 13679 11115 13685
rect 11149 13719 11207 13725
rect 11149 13685 11161 13719
rect 11195 13716 11207 13719
rect 11422 13716 11428 13728
rect 11195 13688 11428 13716
rect 11195 13685 11207 13688
rect 11149 13679 11207 13685
rect 11422 13676 11428 13688
rect 11480 13716 11486 13728
rect 11974 13716 11980 13728
rect 11480 13688 11980 13716
rect 11480 13676 11486 13688
rect 11974 13676 11980 13688
rect 12032 13716 12038 13728
rect 13906 13716 13912 13728
rect 12032 13688 13912 13716
rect 12032 13676 12038 13688
rect 13906 13676 13912 13688
rect 13964 13716 13970 13728
rect 14274 13716 14280 13728
rect 13964 13688 14280 13716
rect 13964 13676 13970 13688
rect 14274 13676 14280 13688
rect 14332 13676 14338 13728
rect 14384 13725 14412 13756
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 15151 13787 15209 13793
rect 15151 13784 15163 13787
rect 15068 13756 15163 13784
rect 15068 13744 15074 13756
rect 15151 13753 15163 13756
rect 15197 13753 15209 13787
rect 17954 13784 17960 13796
rect 17250 13756 17960 13784
rect 15151 13747 15209 13753
rect 17954 13744 17960 13756
rect 18012 13744 18018 13796
rect 18690 13744 18696 13796
rect 18748 13744 18754 13796
rect 22756 13784 22784 13960
rect 22848 13861 22876 14028
rect 25225 14025 25237 14059
rect 25271 14056 25283 14059
rect 25774 14056 25780 14068
rect 25271 14028 25780 14056
rect 25271 14025 25283 14028
rect 25225 14019 25283 14025
rect 25774 14016 25780 14028
rect 25832 14016 25838 14068
rect 26329 14059 26387 14065
rect 26329 14025 26341 14059
rect 26375 14056 26387 14059
rect 26602 14056 26608 14068
rect 26375 14028 26608 14056
rect 26375 14025 26387 14028
rect 26329 14019 26387 14025
rect 26602 14016 26608 14028
rect 26660 14016 26666 14068
rect 27154 14056 27160 14068
rect 26804 14028 27160 14056
rect 26237 13991 26295 13997
rect 26237 13957 26249 13991
rect 26283 13988 26295 13991
rect 26804 13988 26832 14028
rect 27154 14016 27160 14028
rect 27212 14016 27218 14068
rect 27706 14016 27712 14068
rect 27764 14056 27770 14068
rect 27893 14059 27951 14065
rect 27893 14056 27905 14059
rect 27764 14028 27905 14056
rect 27764 14016 27770 14028
rect 27893 14025 27905 14028
rect 27939 14025 27951 14059
rect 27893 14019 27951 14025
rect 29181 14059 29239 14065
rect 29181 14025 29193 14059
rect 29227 14056 29239 14059
rect 29270 14056 29276 14068
rect 29227 14028 29276 14056
rect 29227 14025 29239 14028
rect 29181 14019 29239 14025
rect 29270 14016 29276 14028
rect 29328 14016 29334 14068
rect 29362 14016 29368 14068
rect 29420 14016 29426 14068
rect 29546 14016 29552 14068
rect 29604 14056 29610 14068
rect 30190 14056 30196 14068
rect 29604 14028 30196 14056
rect 29604 14016 29610 14028
rect 30190 14016 30196 14028
rect 30248 14016 30254 14068
rect 30742 14016 30748 14068
rect 30800 14016 30806 14068
rect 31018 14016 31024 14068
rect 31076 14016 31082 14068
rect 26283 13960 26832 13988
rect 26283 13957 26295 13960
rect 26237 13951 26295 13957
rect 26804 13929 26832 13960
rect 27522 13948 27528 14000
rect 27580 13988 27586 14000
rect 28445 13991 28503 13997
rect 28445 13988 28457 13991
rect 27580 13960 28457 13988
rect 27580 13948 27586 13960
rect 28445 13957 28457 13960
rect 28491 13957 28503 13991
rect 28810 13988 28816 14000
rect 28445 13951 28503 13957
rect 28552 13960 28816 13988
rect 26789 13923 26847 13929
rect 26789 13889 26801 13923
rect 26835 13889 26847 13923
rect 26789 13883 26847 13889
rect 26973 13923 27031 13929
rect 26973 13889 26985 13923
rect 27019 13920 27031 13923
rect 27019 13892 27752 13920
rect 27019 13889 27031 13892
rect 26973 13883 27031 13889
rect 22833 13855 22891 13861
rect 22833 13821 22845 13855
rect 22879 13821 22891 13855
rect 23474 13852 23480 13864
rect 22833 13815 22891 13821
rect 22940 13824 23480 13852
rect 22940 13784 22968 13824
rect 23474 13812 23480 13824
rect 23532 13812 23538 13864
rect 23569 13855 23627 13861
rect 23569 13821 23581 13855
rect 23615 13821 23627 13855
rect 23569 13815 23627 13821
rect 22756 13756 22968 13784
rect 23584 13784 23612 13815
rect 25866 13812 25872 13864
rect 25924 13812 25930 13864
rect 26053 13855 26111 13861
rect 26053 13821 26065 13855
rect 26099 13852 26111 13855
rect 26142 13852 26148 13864
rect 26099 13824 26148 13852
rect 26099 13821 26111 13824
rect 26053 13815 26111 13821
rect 26142 13812 26148 13824
rect 26200 13812 26206 13864
rect 26237 13855 26295 13861
rect 26237 13821 26249 13855
rect 26283 13852 26295 13855
rect 26697 13855 26755 13861
rect 26697 13852 26709 13855
rect 26283 13824 26709 13852
rect 26283 13821 26295 13824
rect 26237 13815 26295 13821
rect 26697 13821 26709 13824
rect 26743 13852 26755 13855
rect 27338 13852 27344 13864
rect 26743 13824 27344 13852
rect 26743 13821 26755 13824
rect 26697 13815 26755 13821
rect 27338 13812 27344 13824
rect 27396 13812 27402 13864
rect 27724 13852 27752 13892
rect 27798 13880 27804 13932
rect 27856 13920 27862 13932
rect 28261 13923 28319 13929
rect 28261 13920 28273 13923
rect 27856 13892 28273 13920
rect 27856 13880 27862 13892
rect 28261 13889 28273 13892
rect 28307 13889 28319 13923
rect 28552 13920 28580 13960
rect 28810 13948 28816 13960
rect 28868 13948 28874 14000
rect 28261 13883 28319 13889
rect 28368 13892 28580 13920
rect 29273 13923 29331 13929
rect 27890 13852 27896 13864
rect 27724 13824 27896 13852
rect 27890 13812 27896 13824
rect 27948 13812 27954 13864
rect 28077 13855 28135 13861
rect 28077 13821 28089 13855
rect 28123 13852 28135 13855
rect 28368 13852 28396 13892
rect 29273 13889 29285 13923
rect 29319 13920 29331 13923
rect 29380 13920 29408 14016
rect 29319 13892 29408 13920
rect 29549 13923 29607 13929
rect 29319 13889 29331 13892
rect 29273 13883 29331 13889
rect 29549 13889 29561 13923
rect 29595 13920 29607 13923
rect 30760 13920 30788 14016
rect 29595 13892 30788 13920
rect 29595 13889 29607 13892
rect 29549 13883 29607 13889
rect 28123 13824 28396 13852
rect 28537 13855 28595 13861
rect 28123 13821 28135 13824
rect 28077 13815 28135 13821
rect 28537 13821 28549 13855
rect 28583 13852 28595 13855
rect 28626 13852 28632 13864
rect 28583 13824 28632 13852
rect 28583 13821 28595 13824
rect 28537 13815 28595 13821
rect 24118 13784 24124 13796
rect 23584 13756 24124 13784
rect 24118 13744 24124 13756
rect 24176 13744 24182 13796
rect 24854 13744 24860 13796
rect 24912 13744 24918 13796
rect 26970 13744 26976 13796
rect 27028 13784 27034 13796
rect 28092 13784 28120 13815
rect 28626 13812 28632 13824
rect 28684 13812 28690 13864
rect 28718 13812 28724 13864
rect 28776 13812 28782 13864
rect 28813 13855 28871 13861
rect 28813 13821 28825 13855
rect 28859 13852 28871 13855
rect 28859 13824 28948 13852
rect 28859 13821 28871 13824
rect 28813 13815 28871 13821
rect 27028 13756 28120 13784
rect 27028 13744 27034 13756
rect 14369 13719 14427 13725
rect 14369 13685 14381 13719
rect 14415 13685 14427 13719
rect 14369 13679 14427 13685
rect 16666 13676 16672 13728
rect 16724 13716 16730 13728
rect 17678 13716 17684 13728
rect 16724 13688 17684 13716
rect 16724 13676 16730 13688
rect 17678 13676 17684 13688
rect 17736 13676 17742 13728
rect 19518 13676 19524 13728
rect 19576 13676 19582 13728
rect 20898 13676 20904 13728
rect 20956 13676 20962 13728
rect 21542 13676 21548 13728
rect 21600 13716 21606 13728
rect 21637 13719 21695 13725
rect 21637 13716 21649 13719
rect 21600 13688 21649 13716
rect 21600 13676 21606 13688
rect 21637 13685 21649 13688
rect 21683 13685 21695 13719
rect 21637 13679 21695 13685
rect 23382 13676 23388 13728
rect 23440 13716 23446 13728
rect 23477 13719 23535 13725
rect 23477 13716 23489 13719
rect 23440 13688 23489 13716
rect 23440 13676 23446 13688
rect 23477 13685 23489 13688
rect 23523 13685 23535 13719
rect 23477 13679 23535 13685
rect 27157 13719 27215 13725
rect 27157 13685 27169 13719
rect 27203 13716 27215 13719
rect 27982 13716 27988 13728
rect 27203 13688 27988 13716
rect 27203 13685 27215 13688
rect 27157 13679 27215 13685
rect 27982 13676 27988 13688
rect 28040 13676 28046 13728
rect 28920 13716 28948 13824
rect 28994 13812 29000 13864
rect 29052 13812 29058 13864
rect 30682 13824 31340 13852
rect 30834 13744 30840 13796
rect 30892 13784 30898 13796
rect 31205 13787 31263 13793
rect 31205 13784 31217 13787
rect 30892 13756 31217 13784
rect 30892 13744 30898 13756
rect 31205 13753 31217 13756
rect 31251 13753 31263 13787
rect 31312 13784 31340 13824
rect 31754 13812 31760 13864
rect 31812 13812 31818 13864
rect 31570 13784 31576 13796
rect 31312 13756 31576 13784
rect 31205 13747 31263 13753
rect 31570 13744 31576 13756
rect 31628 13744 31634 13796
rect 30282 13716 30288 13728
rect 28920 13688 30288 13716
rect 30282 13676 30288 13688
rect 30340 13676 30346 13728
rect 2760 13626 32200 13648
rect 2760 13574 6946 13626
rect 6998 13574 7010 13626
rect 7062 13574 7074 13626
rect 7126 13574 7138 13626
rect 7190 13574 7202 13626
rect 7254 13574 14306 13626
rect 14358 13574 14370 13626
rect 14422 13574 14434 13626
rect 14486 13574 14498 13626
rect 14550 13574 14562 13626
rect 14614 13574 21666 13626
rect 21718 13574 21730 13626
rect 21782 13574 21794 13626
rect 21846 13574 21858 13626
rect 21910 13574 21922 13626
rect 21974 13574 29026 13626
rect 29078 13574 29090 13626
rect 29142 13574 29154 13626
rect 29206 13574 29218 13626
rect 29270 13574 29282 13626
rect 29334 13574 32200 13626
rect 2760 13552 32200 13574
rect 7650 13472 7656 13524
rect 7708 13472 7714 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10468 13484 13492 13512
rect 10468 13472 10474 13484
rect 9766 13444 9772 13456
rect 9338 13416 9772 13444
rect 9766 13404 9772 13416
rect 9824 13404 9830 13456
rect 11146 13444 11152 13456
rect 10612 13416 11152 13444
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13376 4491 13379
rect 5994 13376 6000 13388
rect 4479 13348 6000 13376
rect 4479 13345 4491 13348
rect 4433 13339 4491 13345
rect 5994 13336 6000 13348
rect 6052 13336 6058 13388
rect 7561 13379 7619 13385
rect 7561 13345 7573 13379
rect 7607 13345 7619 13379
rect 7561 13339 7619 13345
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 1360 13280 3249 13308
rect 1360 13268 1366 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 7576 13308 7604 13339
rect 10042 13336 10048 13388
rect 10100 13336 10106 13388
rect 10612 13385 10640 13416
rect 11146 13404 11152 13416
rect 11204 13404 11210 13456
rect 11330 13404 11336 13456
rect 11388 13404 11394 13456
rect 12618 13404 12624 13456
rect 12676 13444 12682 13456
rect 12805 13447 12863 13453
rect 12805 13444 12817 13447
rect 12676 13416 12817 13444
rect 12676 13404 12682 13416
rect 12805 13413 12817 13416
rect 12851 13413 12863 13447
rect 12805 13407 12863 13413
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 10597 13339 10655 13345
rect 12894 13336 12900 13388
rect 12952 13336 12958 13388
rect 13464 13385 13492 13484
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14553 13515 14611 13521
rect 13964 13484 14504 13512
rect 13964 13472 13970 13484
rect 14182 13404 14188 13456
rect 14240 13404 14246 13456
rect 13449 13379 13507 13385
rect 13449 13345 13461 13379
rect 13495 13376 13507 13379
rect 14090 13376 14096 13388
rect 13495 13348 14096 13376
rect 13495 13345 13507 13348
rect 13449 13339 13507 13345
rect 14090 13336 14096 13348
rect 14148 13336 14154 13388
rect 14476 13385 14504 13484
rect 14553 13481 14565 13515
rect 14599 13512 14611 13515
rect 15102 13512 15108 13524
rect 14599 13484 15108 13512
rect 14599 13481 14611 13484
rect 14553 13475 14611 13481
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15841 13515 15899 13521
rect 15841 13481 15853 13515
rect 15887 13512 15899 13515
rect 15930 13512 15936 13524
rect 15887 13484 15936 13512
rect 15887 13481 15899 13484
rect 15841 13475 15899 13481
rect 15930 13472 15936 13484
rect 15988 13472 15994 13524
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 16669 13515 16727 13521
rect 16669 13512 16681 13515
rect 16632 13484 16681 13512
rect 16632 13472 16638 13484
rect 16669 13481 16681 13484
rect 16715 13481 16727 13515
rect 16669 13475 16727 13481
rect 16850 13472 16856 13524
rect 16908 13472 16914 13524
rect 17954 13472 17960 13524
rect 18012 13512 18018 13524
rect 18506 13512 18512 13524
rect 18012 13484 18512 13512
rect 18012 13472 18018 13484
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 18874 13472 18880 13524
rect 18932 13472 18938 13524
rect 18969 13515 19027 13521
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19518 13512 19524 13524
rect 19015 13484 19524 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19518 13472 19524 13484
rect 19576 13472 19582 13524
rect 20898 13512 20904 13524
rect 19904 13484 20904 13512
rect 14918 13404 14924 13456
rect 14976 13444 14982 13456
rect 15013 13447 15071 13453
rect 15013 13444 15025 13447
rect 14976 13416 15025 13444
rect 14976 13404 14982 13416
rect 15013 13413 15025 13416
rect 15059 13413 15071 13447
rect 16868 13444 16896 13472
rect 15013 13407 15071 13413
rect 16316 13416 16896 13444
rect 18892 13444 18920 13472
rect 19904 13453 19932 13484
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 21361 13515 21419 13521
rect 21361 13481 21373 13515
rect 21407 13512 21419 13515
rect 22094 13512 22100 13524
rect 21407 13484 22100 13512
rect 21407 13481 21419 13484
rect 21361 13475 21419 13481
rect 22094 13472 22100 13484
rect 22152 13472 22158 13524
rect 23247 13515 23305 13521
rect 23247 13481 23259 13515
rect 23293 13512 23305 13515
rect 24026 13512 24032 13524
rect 23293 13484 24032 13512
rect 23293 13481 23305 13484
rect 23247 13475 23305 13481
rect 24026 13472 24032 13484
rect 24084 13472 24090 13524
rect 24762 13472 24768 13524
rect 24820 13472 24826 13524
rect 24854 13472 24860 13524
rect 24912 13512 24918 13524
rect 24949 13515 25007 13521
rect 24949 13512 24961 13515
rect 24912 13484 24961 13512
rect 24912 13472 24918 13484
rect 24949 13481 24961 13484
rect 24995 13481 25007 13515
rect 24949 13475 25007 13481
rect 25866 13472 25872 13524
rect 25924 13512 25930 13524
rect 25961 13515 26019 13521
rect 25961 13512 25973 13515
rect 25924 13484 25973 13512
rect 25924 13472 25930 13484
rect 25961 13481 25973 13484
rect 26007 13481 26019 13515
rect 25961 13475 26019 13481
rect 26329 13515 26387 13521
rect 26329 13481 26341 13515
rect 26375 13512 26387 13515
rect 26375 13484 28120 13512
rect 26375 13481 26387 13484
rect 26329 13475 26387 13481
rect 19061 13447 19119 13453
rect 19061 13444 19073 13447
rect 18892 13416 19073 13444
rect 14461 13379 14519 13385
rect 14461 13345 14473 13379
rect 14507 13345 14519 13379
rect 14461 13339 14519 13345
rect 14550 13336 14556 13388
rect 14608 13376 14614 13388
rect 14734 13376 14740 13388
rect 14608 13348 14740 13376
rect 14608 13336 14614 13348
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 16022 13336 16028 13388
rect 16080 13336 16086 13388
rect 16114 13336 16120 13388
rect 16172 13336 16178 13388
rect 16316 13385 16344 13416
rect 19061 13413 19073 13416
rect 19107 13413 19119 13447
rect 19061 13407 19119 13413
rect 19889 13447 19947 13453
rect 19889 13413 19901 13447
rect 19935 13413 19947 13447
rect 21450 13444 21456 13456
rect 21114 13416 21456 13444
rect 19889 13407 19947 13413
rect 21450 13404 21456 13416
rect 21508 13404 21514 13456
rect 22646 13404 22652 13456
rect 22704 13404 22710 13456
rect 24118 13404 24124 13456
rect 24176 13444 24182 13456
rect 26344 13444 26372 13475
rect 26970 13444 26976 13456
rect 24176 13416 26372 13444
rect 26528 13416 26976 13444
rect 24176 13404 24182 13416
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13345 16359 13379
rect 16301 13339 16359 13345
rect 16850 13336 16856 13388
rect 16908 13336 16914 13388
rect 17402 13376 17408 13388
rect 17144 13348 17408 13376
rect 8018 13308 8024 13320
rect 7576 13280 8024 13308
rect 3237 13271 3295 13277
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 9766 13268 9772 13320
rect 9824 13268 9830 13320
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13308 10931 13311
rect 10962 13308 10968 13320
rect 10919 13280 10968 13308
rect 10919 13277 10931 13280
rect 10873 13271 10931 13277
rect 10962 13268 10968 13280
rect 11020 13268 11026 13320
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 12621 13311 12679 13317
rect 12621 13308 12633 13311
rect 12584 13280 12633 13308
rect 12584 13268 12590 13280
rect 12621 13277 12633 13280
rect 12667 13277 12679 13311
rect 12621 13271 12679 13277
rect 16209 13311 16267 13317
rect 16209 13277 16221 13311
rect 16255 13308 16267 13311
rect 17144 13308 17172 13348
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 18966 13376 18972 13388
rect 18156 13348 18972 13376
rect 16255 13280 17172 13308
rect 16255 13277 16267 13280
rect 16209 13271 16267 13277
rect 17218 13268 17224 13320
rect 17276 13268 17282 13320
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 7340 13212 8432 13240
rect 7340 13200 7346 13212
rect 8294 13132 8300 13184
rect 8352 13132 8358 13184
rect 8404 13172 8432 13212
rect 13998 13200 14004 13252
rect 14056 13240 14062 13252
rect 14734 13240 14740 13252
rect 14056 13212 14740 13240
rect 14056 13200 14062 13212
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 14921 13243 14979 13249
rect 14921 13209 14933 13243
rect 14967 13240 14979 13243
rect 15289 13243 15347 13249
rect 15289 13240 15301 13243
rect 14967 13212 15301 13240
rect 14967 13209 14979 13212
rect 14921 13203 14979 13209
rect 15289 13209 15301 13212
rect 15335 13209 15347 13243
rect 15289 13203 15347 13209
rect 15396 13212 16528 13240
rect 15396 13172 15424 13212
rect 8404 13144 15424 13172
rect 15473 13175 15531 13181
rect 15473 13141 15485 13175
rect 15519 13172 15531 13175
rect 15746 13172 15752 13184
rect 15519 13144 15752 13172
rect 15519 13141 15531 13144
rect 15473 13135 15531 13141
rect 15746 13132 15752 13144
rect 15804 13132 15810 13184
rect 16500 13172 16528 13212
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 18156 13240 18184 13348
rect 18966 13336 18972 13348
rect 19024 13376 19030 13388
rect 19024 13348 19196 13376
rect 19024 13336 19030 13348
rect 18690 13268 18696 13320
rect 18748 13308 18754 13320
rect 19168 13317 19196 13348
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 24780 13385 24808 13416
rect 23661 13379 23719 13385
rect 23661 13376 23673 13379
rect 23532 13348 23673 13376
rect 23532 13336 23538 13348
rect 23661 13345 23673 13348
rect 23707 13345 23719 13379
rect 23661 13339 23719 13345
rect 24765 13379 24823 13385
rect 24765 13345 24777 13379
rect 24811 13345 24823 13379
rect 24765 13339 24823 13345
rect 25590 13336 25596 13388
rect 25648 13376 25654 13388
rect 26528 13376 26556 13416
rect 26970 13404 26976 13416
rect 27028 13404 27034 13456
rect 27893 13379 27951 13385
rect 27893 13376 27905 13379
rect 25648 13348 26556 13376
rect 26620 13348 27905 13376
rect 25648 13336 25654 13348
rect 19153 13311 19211 13317
rect 18748 13280 19104 13308
rect 18748 13268 18754 13280
rect 19076 13240 19104 13280
rect 19153 13277 19165 13311
rect 19199 13277 19211 13311
rect 19153 13271 19211 13277
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 21358 13308 21364 13320
rect 19659 13280 21364 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 19628 13240 19656 13271
rect 21358 13268 21364 13280
rect 21416 13308 21422 13320
rect 21453 13311 21511 13317
rect 21453 13308 21465 13311
rect 21416 13280 21465 13308
rect 21416 13268 21422 13280
rect 21453 13277 21465 13280
rect 21499 13277 21511 13311
rect 21453 13271 21511 13277
rect 21818 13268 21824 13320
rect 21876 13268 21882 13320
rect 26418 13268 26424 13320
rect 26476 13268 26482 13320
rect 26620 13317 26648 13348
rect 27893 13345 27905 13348
rect 27939 13376 27951 13379
rect 27939 13348 28028 13376
rect 27939 13345 27951 13348
rect 27893 13339 27951 13345
rect 26605 13311 26663 13317
rect 26605 13277 26617 13311
rect 26651 13277 26663 13311
rect 26605 13271 26663 13277
rect 26694 13268 26700 13320
rect 26752 13308 26758 13320
rect 27341 13311 27399 13317
rect 27341 13308 27353 13311
rect 26752 13280 27353 13308
rect 26752 13268 26758 13280
rect 27341 13277 27353 13280
rect 27387 13277 27399 13311
rect 27341 13271 27399 13277
rect 27614 13268 27620 13320
rect 27672 13308 27678 13320
rect 27801 13311 27859 13317
rect 27801 13308 27813 13311
rect 27672 13280 27813 13308
rect 27672 13268 27678 13280
rect 27801 13277 27813 13280
rect 27847 13277 27859 13311
rect 27801 13271 27859 13277
rect 28000 13252 28028 13348
rect 28092 13308 28120 13484
rect 28276 13484 30788 13512
rect 28276 13385 28304 13484
rect 28626 13404 28632 13456
rect 28684 13444 28690 13456
rect 29362 13444 29368 13456
rect 28684 13416 28764 13444
rect 28684 13404 28690 13416
rect 28736 13385 28764 13416
rect 29012 13416 29368 13444
rect 29012 13388 29040 13416
rect 29362 13404 29368 13416
rect 29420 13404 29426 13456
rect 30558 13444 30564 13456
rect 30498 13416 30564 13444
rect 30558 13404 30564 13416
rect 30616 13404 30622 13456
rect 28261 13379 28319 13385
rect 28261 13345 28273 13379
rect 28307 13345 28319 13379
rect 28261 13339 28319 13345
rect 28721 13379 28779 13385
rect 28721 13345 28733 13379
rect 28767 13345 28779 13379
rect 28721 13339 28779 13345
rect 28994 13336 29000 13388
rect 29052 13336 29058 13388
rect 30760 13376 30788 13484
rect 30926 13472 30932 13524
rect 30984 13512 30990 13524
rect 31205 13515 31263 13521
rect 31205 13512 31217 13515
rect 30984 13484 31217 13512
rect 30984 13472 30990 13484
rect 31205 13481 31217 13484
rect 31251 13481 31263 13515
rect 31205 13475 31263 13481
rect 31573 13515 31631 13521
rect 31573 13481 31585 13515
rect 31619 13512 31631 13515
rect 31754 13512 31760 13524
rect 31619 13484 31760 13512
rect 31619 13481 31631 13484
rect 31573 13475 31631 13481
rect 31754 13472 31760 13484
rect 31812 13472 31818 13524
rect 31018 13404 31024 13456
rect 31076 13444 31082 13456
rect 31113 13447 31171 13453
rect 31113 13444 31125 13447
rect 31076 13416 31125 13444
rect 31076 13404 31082 13416
rect 31113 13413 31125 13416
rect 31159 13413 31171 13447
rect 31113 13407 31171 13413
rect 30760 13348 30972 13376
rect 30944 13320 30972 13348
rect 31662 13336 31668 13388
rect 31720 13336 31726 13388
rect 29273 13311 29331 13317
rect 28092 13280 28994 13308
rect 28966 13252 28994 13280
rect 29273 13277 29285 13311
rect 29319 13308 29331 13311
rect 30834 13308 30840 13320
rect 29319 13280 30840 13308
rect 29319 13277 29331 13280
rect 29273 13271 29331 13277
rect 30834 13268 30840 13280
rect 30892 13268 30898 13320
rect 30926 13268 30932 13320
rect 30984 13268 30990 13320
rect 31754 13268 31760 13320
rect 31812 13268 31818 13320
rect 16632 13212 18184 13240
rect 18524 13212 18736 13240
rect 19076 13212 19656 13240
rect 16632 13200 16638 13212
rect 18524 13172 18552 13212
rect 16500 13144 18552 13172
rect 18598 13132 18604 13184
rect 18656 13132 18662 13184
rect 18708 13172 18736 13212
rect 27982 13200 27988 13252
rect 28040 13200 28046 13252
rect 28276 13212 28764 13240
rect 28966 13212 29000 13252
rect 19518 13172 19524 13184
rect 18708 13144 19524 13172
rect 19518 13132 19524 13144
rect 19576 13132 19582 13184
rect 26786 13132 26792 13184
rect 26844 13132 26850 13184
rect 28276 13181 28304 13212
rect 28736 13184 28764 13212
rect 28994 13200 29000 13212
rect 29052 13200 29058 13252
rect 30760 13212 31754 13240
rect 28261 13175 28319 13181
rect 28261 13141 28273 13175
rect 28307 13141 28319 13175
rect 28261 13135 28319 13141
rect 28442 13132 28448 13184
rect 28500 13132 28506 13184
rect 28718 13132 28724 13184
rect 28776 13132 28782 13184
rect 28813 13175 28871 13181
rect 28813 13141 28825 13175
rect 28859 13172 28871 13175
rect 29822 13172 29828 13184
rect 28859 13144 29828 13172
rect 28859 13141 28871 13144
rect 28813 13135 28871 13141
rect 29822 13132 29828 13144
rect 29880 13132 29886 13184
rect 30760 13181 30788 13212
rect 31726 13184 31754 13212
rect 30745 13175 30803 13181
rect 30745 13141 30757 13175
rect 30791 13141 30803 13175
rect 31726 13144 31760 13184
rect 30745 13135 30803 13141
rect 31754 13132 31760 13144
rect 31812 13132 31818 13184
rect 2760 13082 32200 13104
rect 2760 13030 6286 13082
rect 6338 13030 6350 13082
rect 6402 13030 6414 13082
rect 6466 13030 6478 13082
rect 6530 13030 6542 13082
rect 6594 13030 13646 13082
rect 13698 13030 13710 13082
rect 13762 13030 13774 13082
rect 13826 13030 13838 13082
rect 13890 13030 13902 13082
rect 13954 13030 21006 13082
rect 21058 13030 21070 13082
rect 21122 13030 21134 13082
rect 21186 13030 21198 13082
rect 21250 13030 21262 13082
rect 21314 13030 28366 13082
rect 28418 13030 28430 13082
rect 28482 13030 28494 13082
rect 28546 13030 28558 13082
rect 28610 13030 28622 13082
rect 28674 13030 32200 13082
rect 2760 13008 32200 13030
rect 6638 12928 6644 12980
rect 6696 12928 6702 12980
rect 7374 12928 7380 12980
rect 7432 12928 7438 12980
rect 8294 12928 8300 12980
rect 8352 12928 8358 12980
rect 10229 12971 10287 12977
rect 10229 12937 10241 12971
rect 10275 12968 10287 12971
rect 10410 12968 10416 12980
rect 10275 12940 10416 12968
rect 10275 12937 10287 12940
rect 10229 12931 10287 12937
rect 8312 12832 8340 12928
rect 8665 12835 8723 12841
rect 8665 12832 8677 12835
rect 8312 12804 8677 12832
rect 8665 12801 8677 12804
rect 8711 12801 8723 12835
rect 8665 12795 8723 12801
rect 5718 12724 5724 12776
rect 5776 12764 5782 12776
rect 6181 12767 6239 12773
rect 6181 12764 6193 12767
rect 5776 12736 6193 12764
rect 5776 12724 5782 12736
rect 6181 12733 6193 12736
rect 6227 12733 6239 12767
rect 6181 12727 6239 12733
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 8754 12764 8760 12776
rect 7975 12736 8760 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 7852 12696 7880 12727
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9861 12767 9919 12773
rect 9861 12733 9873 12767
rect 9907 12764 9919 12767
rect 10244 12764 10272 12931
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 11606 12928 11612 12980
rect 11664 12928 11670 12980
rect 11882 12928 11888 12980
rect 11940 12968 11946 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11940 12940 11989 12968
rect 11940 12928 11946 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 11977 12931 12035 12937
rect 12161 12971 12219 12977
rect 12161 12937 12173 12971
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 11624 12900 11652 12928
rect 12176 12900 12204 12931
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 14550 12968 14556 12980
rect 13228 12940 14556 12968
rect 13228 12928 13234 12940
rect 14550 12928 14556 12940
rect 14608 12968 14614 12980
rect 15289 12971 15347 12977
rect 15289 12968 15301 12971
rect 14608 12940 15301 12968
rect 14608 12928 14614 12940
rect 15289 12937 15301 12940
rect 15335 12937 15347 12971
rect 15289 12931 15347 12937
rect 16761 12971 16819 12977
rect 16761 12937 16773 12971
rect 16807 12968 16819 12971
rect 16850 12968 16856 12980
rect 16807 12940 16856 12968
rect 16807 12937 16819 12940
rect 16761 12931 16819 12937
rect 16850 12928 16856 12940
rect 16908 12928 16914 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17310 12968 17316 12980
rect 17092 12940 17316 12968
rect 17092 12928 17098 12940
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 17678 12928 17684 12980
rect 17736 12928 17742 12980
rect 18138 12928 18144 12980
rect 18196 12928 18202 12980
rect 20806 12928 20812 12980
rect 20864 12968 20870 12980
rect 20901 12971 20959 12977
rect 20901 12968 20913 12971
rect 20864 12940 20913 12968
rect 20864 12928 20870 12940
rect 20901 12937 20913 12940
rect 20947 12937 20959 12971
rect 21542 12968 21548 12980
rect 20901 12931 20959 12937
rect 21284 12940 21548 12968
rect 11624 12872 12204 12900
rect 12342 12860 12348 12912
rect 12400 12900 12406 12912
rect 12529 12903 12587 12909
rect 12529 12900 12541 12903
rect 12400 12872 12541 12900
rect 12400 12860 12406 12872
rect 12529 12869 12541 12872
rect 12575 12869 12587 12903
rect 13538 12900 13544 12912
rect 12529 12863 12587 12869
rect 13004 12872 13544 12900
rect 13004 12844 13032 12872
rect 13538 12860 13544 12872
rect 13596 12860 13602 12912
rect 17126 12860 17132 12912
rect 17184 12900 17190 12912
rect 17494 12900 17500 12912
rect 17184 12872 17500 12900
rect 17184 12860 17190 12872
rect 17494 12860 17500 12872
rect 17552 12900 17558 12912
rect 17957 12903 18015 12909
rect 17957 12900 17969 12903
rect 17552 12872 17969 12900
rect 17552 12860 17558 12872
rect 17957 12869 17969 12872
rect 18003 12869 18015 12903
rect 17957 12863 18015 12869
rect 10870 12792 10876 12844
rect 10928 12832 10934 12844
rect 12066 12832 12072 12844
rect 10928 12804 12072 12832
rect 10928 12792 10934 12804
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 12986 12792 12992 12844
rect 13044 12792 13050 12844
rect 14182 12792 14188 12844
rect 14240 12832 14246 12844
rect 15010 12832 15016 12844
rect 14240 12804 15016 12832
rect 14240 12792 14246 12804
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 16942 12832 16948 12844
rect 16408 12804 16948 12832
rect 9907 12736 10272 12764
rect 9907 12733 9919 12736
rect 9861 12727 9919 12733
rect 10778 12724 10784 12776
rect 10836 12764 10842 12776
rect 11606 12764 11612 12776
rect 10836 12736 11612 12764
rect 10836 12724 10842 12736
rect 11606 12724 11612 12736
rect 11664 12724 11670 12776
rect 8018 12696 8024 12708
rect 7852 12668 8024 12696
rect 8018 12656 8024 12668
rect 8076 12656 8082 12708
rect 8478 12656 8484 12708
rect 8536 12696 8542 12708
rect 9033 12699 9091 12705
rect 9033 12696 9045 12699
rect 8536 12668 9045 12696
rect 8536 12656 8542 12668
rect 9033 12665 9045 12668
rect 9079 12665 9091 12699
rect 9033 12659 9091 12665
rect 12158 12656 12164 12708
rect 12216 12656 12222 12708
rect 12897 12699 12955 12705
rect 12897 12665 12909 12699
rect 12943 12696 12955 12699
rect 13170 12696 13176 12708
rect 12943 12668 13176 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 13170 12656 13176 12668
rect 13228 12656 13234 12708
rect 13998 12656 14004 12708
rect 14056 12656 14062 12708
rect 14642 12656 14648 12708
rect 14700 12696 14706 12708
rect 14737 12699 14795 12705
rect 14737 12696 14749 12699
rect 14700 12668 14749 12696
rect 14700 12656 14706 12668
rect 14737 12665 14749 12668
rect 14783 12665 14795 12699
rect 14737 12659 14795 12665
rect 5626 12588 5632 12640
rect 5684 12588 5690 12640
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7009 12631 7067 12637
rect 7009 12628 7021 12631
rect 6972 12600 7021 12628
rect 6972 12588 6978 12600
rect 7009 12597 7021 12600
rect 7055 12597 7067 12631
rect 7009 12591 7067 12597
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 8113 12631 8171 12637
rect 8113 12628 8125 12631
rect 7984 12600 8125 12628
rect 7984 12588 7990 12600
rect 8113 12597 8125 12600
rect 8159 12628 8171 12631
rect 8570 12628 8576 12640
rect 8159 12600 8576 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8570 12588 8576 12600
rect 8628 12588 8634 12640
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11698 12628 11704 12640
rect 11204 12600 11704 12628
rect 11204 12588 11210 12600
rect 11698 12588 11704 12600
rect 11756 12628 11762 12640
rect 16408 12637 16436 12804
rect 16942 12792 16948 12804
rect 17000 12832 17006 12844
rect 18156 12832 18184 12928
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 17000 12804 17264 12832
rect 18156 12804 18245 12832
rect 17000 12792 17006 12804
rect 16666 12724 16672 12776
rect 16724 12764 16730 12776
rect 17034 12764 17040 12776
rect 16724 12736 17040 12764
rect 16724 12724 16730 12736
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17236 12773 17264 12804
rect 18233 12801 18245 12804
rect 18279 12832 18291 12835
rect 18598 12832 18604 12844
rect 18279 12804 18604 12832
rect 18279 12801 18291 12804
rect 18233 12795 18291 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12733 17279 12767
rect 17221 12727 17279 12733
rect 17405 12767 17463 12773
rect 17405 12733 17417 12767
rect 17451 12764 17463 12767
rect 17954 12764 17960 12776
rect 17451 12736 17960 12764
rect 17451 12733 17463 12736
rect 17405 12727 17463 12733
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 21284 12773 21312 12940
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 21818 12928 21824 12980
rect 21876 12928 21882 12980
rect 24305 12971 24363 12977
rect 24305 12937 24317 12971
rect 24351 12968 24363 12971
rect 25590 12968 25596 12980
rect 24351 12940 25596 12968
rect 24351 12937 24363 12940
rect 24305 12931 24363 12937
rect 25590 12928 25596 12940
rect 25648 12928 25654 12980
rect 26316 12971 26374 12977
rect 26316 12937 26328 12971
rect 26362 12968 26374 12971
rect 26786 12968 26792 12980
rect 26362 12940 26792 12968
rect 26362 12937 26374 12940
rect 26316 12931 26374 12937
rect 26786 12928 26792 12940
rect 26844 12928 26850 12980
rect 26878 12928 26884 12980
rect 26936 12968 26942 12980
rect 27893 12971 27951 12977
rect 27893 12968 27905 12971
rect 26936 12940 27905 12968
rect 26936 12928 26942 12940
rect 27893 12937 27905 12940
rect 27939 12937 27951 12971
rect 27893 12931 27951 12937
rect 28997 12971 29055 12977
rect 28997 12937 29009 12971
rect 29043 12968 29055 12971
rect 29454 12968 29460 12980
rect 29043 12940 29460 12968
rect 29043 12937 29055 12940
rect 28997 12931 29055 12937
rect 29454 12928 29460 12940
rect 29512 12928 29518 12980
rect 30650 12928 30656 12980
rect 30708 12968 30714 12980
rect 30837 12971 30895 12977
rect 30837 12968 30849 12971
rect 30708 12940 30849 12968
rect 30708 12928 30714 12940
rect 30837 12937 30849 12940
rect 30883 12937 30895 12971
rect 30837 12931 30895 12937
rect 21358 12860 21364 12912
rect 21416 12900 21422 12912
rect 21416 12872 22600 12900
rect 21416 12860 21422 12872
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 22002 12832 22008 12844
rect 21560 12804 22008 12832
rect 18141 12767 18199 12773
rect 18141 12733 18153 12767
rect 18187 12764 18199 12767
rect 21269 12767 21327 12773
rect 18187 12736 18276 12764
rect 18187 12733 18199 12736
rect 18141 12727 18199 12733
rect 18248 12708 18276 12736
rect 21269 12733 21281 12767
rect 21315 12733 21327 12767
rect 21269 12727 21327 12733
rect 17129 12699 17187 12705
rect 17129 12665 17141 12699
rect 17175 12665 17187 12699
rect 18046 12696 18052 12708
rect 17129 12659 17187 12665
rect 17604 12668 18052 12696
rect 16025 12631 16083 12637
rect 16025 12628 16037 12631
rect 11756 12600 16037 12628
rect 11756 12588 11762 12600
rect 16025 12597 16037 12600
rect 16071 12628 16083 12631
rect 16393 12631 16451 12637
rect 16393 12628 16405 12631
rect 16071 12600 16405 12628
rect 16071 12597 16083 12600
rect 16025 12591 16083 12597
rect 16393 12597 16405 12600
rect 16439 12597 16451 12631
rect 16393 12591 16451 12597
rect 16850 12588 16856 12640
rect 16908 12588 16914 12640
rect 17144 12628 17172 12659
rect 17604 12628 17632 12668
rect 18046 12656 18052 12668
rect 18104 12656 18110 12708
rect 18230 12656 18236 12708
rect 18288 12656 18294 12708
rect 18414 12656 18420 12708
rect 18472 12696 18478 12708
rect 18509 12699 18567 12705
rect 18509 12696 18521 12699
rect 18472 12668 18521 12696
rect 18472 12656 18478 12668
rect 18509 12665 18521 12668
rect 18555 12665 18567 12699
rect 20162 12696 20168 12708
rect 19734 12668 20168 12696
rect 18509 12659 18567 12665
rect 20162 12656 20168 12668
rect 20220 12656 20226 12708
rect 21361 12699 21419 12705
rect 21361 12665 21373 12699
rect 21407 12696 21419 12699
rect 21560 12696 21588 12804
rect 22002 12792 22008 12804
rect 22060 12792 22066 12844
rect 22572 12841 22600 12872
rect 27540 12872 29132 12900
rect 22557 12835 22615 12841
rect 22557 12801 22569 12835
rect 22603 12801 22615 12835
rect 22557 12795 22615 12801
rect 26050 12792 26056 12844
rect 26108 12832 26114 12844
rect 26326 12832 26332 12844
rect 26108 12804 26332 12832
rect 26108 12792 26114 12804
rect 26326 12792 26332 12804
rect 26384 12832 26390 12844
rect 27540 12832 27568 12872
rect 29104 12844 29132 12872
rect 26384 12804 27568 12832
rect 26384 12792 26390 12804
rect 27798 12792 27804 12844
rect 27856 12832 27862 12844
rect 28077 12835 28135 12841
rect 28077 12832 28089 12835
rect 27856 12804 28089 12832
rect 27856 12792 27862 12804
rect 28077 12801 28089 12804
rect 28123 12801 28135 12835
rect 28077 12795 28135 12801
rect 28166 12792 28172 12844
rect 28224 12792 28230 12844
rect 29086 12792 29092 12844
rect 29144 12792 29150 12844
rect 30098 12792 30104 12844
rect 30156 12832 30162 12844
rect 31757 12835 31815 12841
rect 31757 12832 31769 12835
rect 30156 12804 31769 12832
rect 30156 12792 30162 12804
rect 31757 12801 31769 12804
rect 31803 12801 31815 12835
rect 31757 12795 31815 12801
rect 22370 12724 22376 12776
rect 22428 12724 22434 12776
rect 23934 12724 23940 12776
rect 23992 12724 23998 12776
rect 25685 12767 25743 12773
rect 25685 12733 25697 12767
rect 25731 12764 25743 12767
rect 25774 12764 25780 12776
rect 25731 12736 25780 12764
rect 25731 12733 25743 12736
rect 25685 12727 25743 12733
rect 25774 12724 25780 12736
rect 25832 12724 25838 12776
rect 28261 12767 28319 12773
rect 28261 12733 28273 12767
rect 28307 12733 28319 12767
rect 28261 12727 28319 12733
rect 21407 12668 21588 12696
rect 21407 12665 21419 12668
rect 21361 12659 21419 12665
rect 22830 12656 22836 12708
rect 22888 12656 22894 12708
rect 26234 12696 26240 12708
rect 24136 12668 26240 12696
rect 17144 12600 17632 12628
rect 19981 12631 20039 12637
rect 19981 12597 19993 12631
rect 20027 12628 20039 12631
rect 20070 12628 20076 12640
rect 20027 12600 20076 12628
rect 20027 12597 20039 12600
rect 19981 12591 20039 12597
rect 20070 12588 20076 12600
rect 20128 12628 20134 12640
rect 24136 12628 24164 12668
rect 26234 12656 26240 12668
rect 26292 12656 26298 12708
rect 26436 12668 26818 12696
rect 20128 12600 24164 12628
rect 25777 12631 25835 12637
rect 20128 12588 20134 12600
rect 25777 12597 25789 12631
rect 25823 12628 25835 12631
rect 26436 12628 26464 12668
rect 27614 12656 27620 12708
rect 27672 12696 27678 12708
rect 27672 12668 27936 12696
rect 27672 12656 27678 12668
rect 25823 12600 26464 12628
rect 25823 12597 25835 12600
rect 25777 12591 25835 12597
rect 27798 12588 27804 12640
rect 27856 12588 27862 12640
rect 27908 12628 27936 12668
rect 28074 12656 28080 12708
rect 28132 12696 28138 12708
rect 28276 12696 28304 12727
rect 28350 12724 28356 12776
rect 28408 12724 28414 12776
rect 28624 12767 28682 12773
rect 28624 12733 28636 12767
rect 28670 12764 28682 12767
rect 28670 12736 29132 12764
rect 28670 12733 28682 12736
rect 28624 12727 28682 12733
rect 28132 12668 28304 12696
rect 28721 12699 28779 12705
rect 28132 12656 28138 12668
rect 28721 12665 28733 12699
rect 28767 12665 28779 12699
rect 28721 12659 28779 12665
rect 28166 12628 28172 12640
rect 27908 12600 28172 12628
rect 28166 12588 28172 12600
rect 28224 12588 28230 12640
rect 28626 12588 28632 12640
rect 28684 12628 28690 12640
rect 28736 12628 28764 12659
rect 28810 12656 28816 12708
rect 28868 12656 28874 12708
rect 28997 12699 29055 12705
rect 28997 12665 29009 12699
rect 29043 12665 29055 12699
rect 29104 12696 29132 12736
rect 29270 12696 29276 12708
rect 29104 12668 29276 12696
rect 28997 12659 29055 12665
rect 28684 12600 28764 12628
rect 29012 12628 29040 12659
rect 29270 12656 29276 12668
rect 29328 12656 29334 12708
rect 29365 12699 29423 12705
rect 29365 12665 29377 12699
rect 29411 12696 29423 12699
rect 29638 12696 29644 12708
rect 29411 12668 29644 12696
rect 29411 12665 29423 12668
rect 29365 12659 29423 12665
rect 29638 12656 29644 12668
rect 29696 12656 29702 12708
rect 29822 12656 29828 12708
rect 29880 12656 29886 12708
rect 30650 12628 30656 12640
rect 29012 12600 30656 12628
rect 28684 12588 28690 12600
rect 30650 12588 30656 12600
rect 30708 12628 30714 12640
rect 31205 12631 31263 12637
rect 31205 12628 31217 12631
rect 30708 12600 31217 12628
rect 30708 12588 30714 12600
rect 31205 12597 31217 12600
rect 31251 12597 31263 12631
rect 31205 12591 31263 12597
rect 2760 12538 32200 12560
rect 2760 12486 6946 12538
rect 6998 12486 7010 12538
rect 7062 12486 7074 12538
rect 7126 12486 7138 12538
rect 7190 12486 7202 12538
rect 7254 12486 14306 12538
rect 14358 12486 14370 12538
rect 14422 12486 14434 12538
rect 14486 12486 14498 12538
rect 14550 12486 14562 12538
rect 14614 12486 21666 12538
rect 21718 12486 21730 12538
rect 21782 12486 21794 12538
rect 21846 12486 21858 12538
rect 21910 12486 21922 12538
rect 21974 12486 29026 12538
rect 29078 12486 29090 12538
rect 29142 12486 29154 12538
rect 29206 12486 29218 12538
rect 29270 12486 29282 12538
rect 29334 12486 32200 12538
rect 2760 12464 32200 12486
rect 5718 12384 5724 12436
rect 5776 12384 5782 12436
rect 6181 12427 6239 12433
rect 6181 12393 6193 12427
rect 6227 12424 6239 12427
rect 7926 12424 7932 12436
rect 6227 12396 7932 12424
rect 6227 12393 6239 12396
rect 6181 12387 6239 12393
rect 7926 12384 7932 12396
rect 7984 12384 7990 12436
rect 8110 12384 8116 12436
rect 8168 12384 8174 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 8628 12396 9628 12424
rect 8628 12384 8634 12396
rect 4338 12316 4344 12368
rect 4396 12316 4402 12368
rect 5353 12359 5411 12365
rect 5353 12325 5365 12359
rect 5399 12356 5411 12359
rect 5626 12356 5632 12368
rect 5399 12328 5632 12356
rect 5399 12325 5411 12328
rect 5353 12319 5411 12325
rect 5626 12316 5632 12328
rect 5684 12316 5690 12368
rect 6914 12316 6920 12368
rect 6972 12316 6978 12368
rect 7834 12316 7840 12368
rect 7892 12356 7898 12368
rect 8128 12356 8156 12384
rect 7892 12328 8156 12356
rect 7892 12316 7898 12328
rect 8754 12316 8760 12368
rect 8812 12316 8818 12368
rect 9600 12356 9628 12396
rect 9766 12384 9772 12436
rect 9824 12424 9830 12436
rect 9861 12427 9919 12433
rect 9861 12424 9873 12427
rect 9824 12396 9873 12424
rect 9824 12384 9830 12396
rect 9861 12393 9873 12396
rect 9907 12393 9919 12427
rect 9861 12387 9919 12393
rect 11606 12384 11612 12436
rect 11664 12424 11670 12436
rect 12434 12424 12440 12436
rect 11664 12396 12440 12424
rect 11664 12384 11670 12396
rect 12434 12384 12440 12396
rect 12492 12424 12498 12436
rect 12492 12396 12940 12424
rect 12492 12384 12498 12396
rect 10413 12359 10471 12365
rect 10413 12356 10425 12359
rect 9600 12328 10425 12356
rect 10413 12325 10425 12328
rect 10459 12325 10471 12359
rect 10413 12319 10471 12325
rect 11146 12316 11152 12368
rect 11204 12356 11210 12368
rect 11698 12356 11704 12368
rect 11204 12328 11704 12356
rect 11204 12316 11210 12328
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 12250 12316 12256 12368
rect 12308 12316 12314 12368
rect 12912 12356 12940 12396
rect 12986 12384 12992 12436
rect 13044 12384 13050 12436
rect 13096 12396 16160 12424
rect 13096 12356 13124 12396
rect 12912 12328 13124 12356
rect 14090 12316 14096 12368
rect 14148 12316 14154 12368
rect 14277 12359 14335 12365
rect 14277 12325 14289 12359
rect 14323 12356 14335 12359
rect 14642 12356 14648 12368
rect 14323 12328 14648 12356
rect 14323 12325 14335 12328
rect 14277 12319 14335 12325
rect 14642 12316 14648 12328
rect 14700 12316 14706 12368
rect 15378 12316 15384 12368
rect 15436 12316 15442 12368
rect 15746 12316 15752 12368
rect 15804 12356 15810 12368
rect 16025 12359 16083 12365
rect 16025 12356 16037 12359
rect 15804 12328 16037 12356
rect 15804 12316 15810 12328
rect 16025 12325 16037 12328
rect 16071 12325 16083 12359
rect 16132 12356 16160 12396
rect 18414 12384 18420 12436
rect 18472 12424 18478 12436
rect 18601 12427 18659 12433
rect 18601 12424 18613 12427
rect 18472 12396 18613 12424
rect 18472 12384 18478 12396
rect 18601 12393 18613 12396
rect 18647 12393 18659 12427
rect 18601 12387 18659 12393
rect 18966 12384 18972 12436
rect 19024 12384 19030 12436
rect 20162 12384 20168 12436
rect 20220 12384 20226 12436
rect 20622 12384 20628 12436
rect 20680 12384 20686 12436
rect 22005 12427 22063 12433
rect 22005 12393 22017 12427
rect 22051 12424 22063 12427
rect 22370 12424 22376 12436
rect 22051 12396 22376 12424
rect 22051 12393 22063 12396
rect 22005 12387 22063 12393
rect 22370 12384 22376 12396
rect 22428 12384 22434 12436
rect 22646 12384 22652 12436
rect 22704 12384 22710 12436
rect 22738 12384 22744 12436
rect 22796 12384 22802 12436
rect 22922 12384 22928 12436
rect 22980 12384 22986 12436
rect 23750 12424 23756 12436
rect 23400 12396 23756 12424
rect 18984 12356 19012 12384
rect 16132 12328 19012 12356
rect 16025 12319 16083 12325
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 6089 12291 6147 12297
rect 6089 12288 6101 12291
rect 5776 12260 6101 12288
rect 5776 12248 5782 12260
rect 6089 12257 6101 12260
rect 6135 12257 6147 12291
rect 6089 12251 6147 12257
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12257 6791 12291
rect 6733 12251 6791 12257
rect 3881 12223 3939 12229
rect 3881 12189 3893 12223
rect 3927 12220 3939 12223
rect 3927 12192 5580 12220
rect 3927 12189 3939 12192
rect 3881 12183 3939 12189
rect 5552 12152 5580 12192
rect 5626 12180 5632 12232
rect 5684 12180 5690 12232
rect 5736 12152 5764 12248
rect 6365 12223 6423 12229
rect 6365 12189 6377 12223
rect 6411 12220 6423 12223
rect 6638 12220 6644 12232
rect 6411 12192 6644 12220
rect 6411 12189 6423 12192
rect 6365 12183 6423 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6748 12220 6776 12251
rect 6822 12248 6828 12300
rect 6880 12248 6886 12300
rect 7098 12248 7104 12300
rect 7156 12248 7162 12300
rect 7374 12288 7380 12300
rect 7208 12260 7380 12288
rect 7208 12220 7236 12260
rect 7374 12248 7380 12260
rect 7432 12288 7438 12300
rect 7926 12288 7932 12300
rect 7432 12260 7932 12288
rect 7432 12248 7438 12260
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 8018 12248 8024 12300
rect 8076 12248 8082 12300
rect 10134 12248 10140 12300
rect 10192 12248 10198 12300
rect 10870 12288 10876 12300
rect 10428 12260 10876 12288
rect 6748 12192 7236 12220
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12220 7895 12223
rect 8297 12223 8355 12229
rect 8297 12220 8309 12223
rect 7883 12192 8309 12220
rect 7883 12189 7895 12192
rect 7837 12183 7895 12189
rect 8297 12189 8309 12192
rect 8343 12189 8355 12223
rect 8297 12183 8355 12189
rect 5552 12124 5764 12152
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 6549 12087 6607 12093
rect 6549 12084 6561 12087
rect 4764 12056 6561 12084
rect 4764 12044 4770 12056
rect 6549 12053 6561 12056
rect 6595 12053 6607 12087
rect 7300 12084 7328 12183
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10428 12220 10456 12260
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 16850 12248 16856 12300
rect 16908 12248 16914 12300
rect 18598 12248 18604 12300
rect 18656 12288 18662 12300
rect 19153 12291 19211 12297
rect 19153 12288 19165 12291
rect 18656 12260 19165 12288
rect 18656 12248 18662 12260
rect 19153 12257 19165 12260
rect 19199 12257 19211 12291
rect 19153 12251 19211 12257
rect 19242 12248 19248 12300
rect 19300 12288 19306 12300
rect 20257 12291 20315 12297
rect 20257 12288 20269 12291
rect 19300 12260 20269 12288
rect 19300 12248 19306 12260
rect 20257 12257 20269 12260
rect 20303 12288 20315 12291
rect 20640 12288 20668 12384
rect 21450 12316 21456 12368
rect 21508 12356 21514 12368
rect 21821 12359 21879 12365
rect 21821 12356 21833 12359
rect 21508 12328 21833 12356
rect 21508 12316 21514 12328
rect 21821 12325 21833 12328
rect 21867 12356 21879 12359
rect 22094 12356 22100 12368
rect 21867 12328 22100 12356
rect 21867 12325 21879 12328
rect 21821 12319 21879 12325
rect 22094 12316 22100 12328
rect 22152 12316 22158 12368
rect 22278 12316 22284 12368
rect 22336 12316 22342 12368
rect 22756 12356 22784 12384
rect 23400 12356 23428 12396
rect 23750 12384 23756 12396
rect 23808 12384 23814 12436
rect 23934 12384 23940 12436
rect 23992 12424 23998 12436
rect 24029 12427 24087 12433
rect 24029 12424 24041 12427
rect 23992 12396 24041 12424
rect 23992 12384 23998 12396
rect 24029 12393 24041 12396
rect 24075 12393 24087 12427
rect 24029 12387 24087 12393
rect 24118 12384 24124 12436
rect 24176 12384 24182 12436
rect 24854 12384 24860 12436
rect 24912 12424 24918 12436
rect 25682 12424 25688 12436
rect 24912 12396 25688 12424
rect 24912 12384 24918 12396
rect 25682 12384 25688 12396
rect 25740 12384 25746 12436
rect 26053 12427 26111 12433
rect 26053 12393 26065 12427
rect 26099 12424 26111 12427
rect 26694 12424 26700 12436
rect 26099 12396 26700 12424
rect 26099 12393 26111 12396
rect 26053 12387 26111 12393
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 27617 12427 27675 12433
rect 27617 12424 27629 12427
rect 26804 12396 27108 12424
rect 22756 12328 23428 12356
rect 20303 12260 20668 12288
rect 22189 12291 22247 12297
rect 20303 12257 20315 12260
rect 20257 12251 20315 12257
rect 22189 12257 22201 12291
rect 22235 12257 22247 12291
rect 22296 12288 22324 12316
rect 22756 12297 22784 12328
rect 23474 12316 23480 12368
rect 23532 12356 23538 12368
rect 23845 12359 23903 12365
rect 23845 12356 23857 12359
rect 23532 12328 23857 12356
rect 23532 12316 23538 12328
rect 23845 12325 23857 12328
rect 23891 12325 23903 12359
rect 24136 12356 24164 12384
rect 23845 12319 23903 12325
rect 24044 12328 24164 12356
rect 25225 12359 25283 12365
rect 22373 12291 22431 12297
rect 22373 12288 22385 12291
rect 22296 12260 22385 12288
rect 22189 12251 22247 12257
rect 22373 12257 22385 12260
rect 22419 12257 22431 12291
rect 22373 12251 22431 12257
rect 22465 12291 22523 12297
rect 22465 12257 22477 12291
rect 22511 12288 22523 12291
rect 22741 12291 22799 12297
rect 22511 12260 22692 12288
rect 22511 12257 22523 12260
rect 22465 12251 22523 12257
rect 10100 12192 10456 12220
rect 10100 12180 10106 12192
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 10781 12223 10839 12229
rect 10781 12220 10793 12223
rect 10560 12192 10793 12220
rect 10560 12180 10566 12192
rect 10781 12189 10793 12192
rect 10827 12220 10839 12223
rect 12618 12220 12624 12232
rect 10827 12192 12624 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 12618 12180 12624 12192
rect 12676 12180 12682 12232
rect 13078 12180 13084 12232
rect 13136 12220 13142 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 13136 12192 13277 12220
rect 13136 12180 13142 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 15286 12220 15292 12232
rect 13265 12183 13323 12189
rect 13832 12192 15292 12220
rect 9674 12112 9680 12164
rect 9732 12152 9738 12164
rect 13832 12152 13860 12192
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 16298 12180 16304 12232
rect 16356 12180 16362 12232
rect 16942 12180 16948 12232
rect 17000 12220 17006 12232
rect 17497 12223 17555 12229
rect 17497 12220 17509 12223
rect 17000 12192 17509 12220
rect 17000 12180 17006 12192
rect 17497 12189 17509 12192
rect 17543 12189 17555 12223
rect 17497 12183 17555 12189
rect 19426 12180 19432 12232
rect 19484 12180 19490 12232
rect 9732 12124 13860 12152
rect 9732 12112 9738 12124
rect 8846 12084 8852 12096
rect 7300 12056 8852 12084
rect 6549 12047 6607 12053
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 9766 12044 9772 12096
rect 9824 12044 9830 12096
rect 12618 12044 12624 12096
rect 12676 12044 12682 12096
rect 16666 12044 16672 12096
rect 16724 12084 16730 12096
rect 16850 12084 16856 12096
rect 16724 12056 16856 12084
rect 16724 12044 16730 12056
rect 16850 12044 16856 12056
rect 16908 12044 16914 12096
rect 17402 12044 17408 12096
rect 17460 12044 17466 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 19058 12084 19064 12096
rect 18196 12056 19064 12084
rect 18196 12044 18202 12056
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19978 12044 19984 12096
rect 20036 12044 20042 12096
rect 22204 12084 22232 12251
rect 22664 12152 22692 12260
rect 22741 12257 22753 12291
rect 22787 12257 22799 12291
rect 22741 12251 22799 12257
rect 22830 12248 22836 12300
rect 22888 12248 22894 12300
rect 23017 12291 23075 12297
rect 23017 12257 23029 12291
rect 23063 12288 23075 12291
rect 23382 12288 23388 12300
rect 23063 12260 23388 12288
rect 23063 12257 23075 12260
rect 23017 12251 23075 12257
rect 23382 12248 23388 12260
rect 23440 12248 23446 12300
rect 23661 12291 23719 12297
rect 23661 12257 23673 12291
rect 23707 12288 23719 12291
rect 24044 12288 24072 12328
rect 25225 12325 25237 12359
rect 25271 12356 25283 12359
rect 25777 12359 25835 12365
rect 25777 12356 25789 12359
rect 25271 12328 25789 12356
rect 25271 12325 25283 12328
rect 25225 12319 25283 12325
rect 25777 12325 25789 12328
rect 25823 12325 25835 12359
rect 25777 12319 25835 12325
rect 26326 12316 26332 12368
rect 26384 12316 26390 12368
rect 26602 12316 26608 12368
rect 26660 12356 26666 12368
rect 26804 12356 26832 12396
rect 26660 12328 26832 12356
rect 26660 12316 26666 12328
rect 26878 12316 26884 12368
rect 26936 12316 26942 12368
rect 23707 12260 24072 12288
rect 24121 12291 24179 12297
rect 23707 12257 23719 12260
rect 23661 12251 23719 12257
rect 24121 12257 24133 12291
rect 24167 12257 24179 12291
rect 24121 12251 24179 12257
rect 23400 12220 23428 12248
rect 23400 12192 23704 12220
rect 23676 12152 23704 12192
rect 23750 12180 23756 12232
rect 23808 12220 23814 12232
rect 24136 12220 24164 12251
rect 24946 12248 24952 12300
rect 25004 12288 25010 12300
rect 25133 12291 25191 12297
rect 25133 12288 25145 12291
rect 25004 12260 25145 12288
rect 25004 12248 25010 12260
rect 25133 12257 25145 12260
rect 25179 12257 25191 12291
rect 25547 12291 25605 12297
rect 25547 12288 25559 12291
rect 25133 12251 25191 12257
rect 25332 12260 25559 12288
rect 23808 12192 24164 12220
rect 23808 12180 23814 12192
rect 25332 12152 25360 12260
rect 25547 12257 25559 12260
rect 25593 12257 25605 12291
rect 25547 12251 25605 12257
rect 25682 12248 25688 12300
rect 25740 12248 25746 12300
rect 25869 12291 25927 12297
rect 25869 12257 25881 12291
rect 25915 12288 25927 12291
rect 26896 12288 26924 12316
rect 25915 12260 26924 12288
rect 25915 12257 25927 12260
rect 25869 12251 25927 12257
rect 26970 12248 26976 12300
rect 27028 12288 27034 12300
rect 27080 12297 27108 12396
rect 27448 12396 27629 12424
rect 27448 12356 27476 12396
rect 27617 12393 27629 12396
rect 27663 12393 27675 12427
rect 27617 12387 27675 12393
rect 28626 12384 28632 12436
rect 28684 12424 28690 12436
rect 29730 12424 29736 12436
rect 28684 12396 29736 12424
rect 28684 12384 28690 12396
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 28350 12356 28356 12368
rect 27448 12328 28356 12356
rect 27065 12291 27123 12297
rect 27065 12288 27077 12291
rect 27028 12260 27077 12288
rect 27028 12248 27034 12260
rect 27065 12257 27077 12260
rect 27111 12288 27123 12291
rect 27341 12291 27399 12297
rect 27341 12288 27353 12291
rect 27111 12260 27353 12288
rect 27111 12257 27123 12260
rect 27065 12251 27123 12257
rect 27341 12257 27353 12260
rect 27387 12257 27399 12291
rect 27341 12251 27399 12257
rect 27448 12232 27476 12328
rect 28350 12316 28356 12328
rect 28408 12316 28414 12368
rect 28718 12316 28724 12368
rect 28776 12356 28782 12368
rect 28776 12328 29500 12356
rect 28776 12316 28782 12328
rect 27798 12248 27804 12300
rect 27856 12248 27862 12300
rect 29178 12248 29184 12300
rect 29236 12248 29242 12300
rect 29472 12297 29500 12328
rect 29546 12316 29552 12368
rect 29604 12316 29610 12368
rect 30098 12356 30104 12368
rect 29656 12328 30104 12356
rect 29457 12291 29515 12297
rect 29457 12257 29469 12291
rect 29503 12257 29515 12291
rect 29457 12251 29515 12257
rect 25409 12223 25467 12229
rect 25409 12189 25421 12223
rect 25455 12220 25467 12223
rect 27430 12220 27436 12232
rect 25455 12192 27436 12220
rect 25455 12189 25467 12192
rect 25409 12183 25467 12189
rect 27430 12180 27436 12192
rect 27488 12180 27494 12232
rect 29089 12223 29147 12229
rect 29089 12189 29101 12223
rect 29135 12220 29147 12223
rect 29564 12220 29592 12316
rect 29656 12297 29684 12328
rect 30098 12316 30104 12328
rect 30156 12316 30162 12368
rect 29641 12291 29699 12297
rect 29641 12257 29653 12291
rect 29687 12257 29699 12291
rect 29641 12251 29699 12257
rect 29730 12248 29736 12300
rect 29788 12288 29794 12300
rect 29825 12291 29883 12297
rect 29825 12288 29837 12291
rect 29788 12260 29837 12288
rect 29788 12248 29794 12260
rect 29825 12257 29837 12260
rect 29871 12257 29883 12291
rect 29825 12251 29883 12257
rect 30190 12248 30196 12300
rect 30248 12248 30254 12300
rect 30469 12291 30527 12297
rect 30469 12257 30481 12291
rect 30515 12257 30527 12291
rect 30469 12251 30527 12257
rect 31665 12291 31723 12297
rect 31665 12257 31677 12291
rect 31711 12288 31723 12291
rect 33134 12288 33140 12300
rect 31711 12260 33140 12288
rect 31711 12257 31723 12260
rect 31665 12251 31723 12257
rect 29135 12192 29592 12220
rect 29135 12189 29147 12192
rect 29089 12183 29147 12189
rect 26142 12152 26148 12164
rect 22664 12124 23520 12152
rect 23676 12124 26148 12152
rect 23492 12096 23520 12124
rect 26142 12112 26148 12124
rect 26200 12112 26206 12164
rect 26234 12112 26240 12164
rect 26292 12152 26298 12164
rect 30484 12152 30512 12251
rect 33134 12248 33140 12260
rect 33192 12248 33198 12300
rect 26292 12124 30512 12152
rect 26292 12112 26298 12124
rect 22830 12084 22836 12096
rect 22204 12056 22836 12084
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 23474 12044 23480 12096
rect 23532 12044 23538 12096
rect 25130 12044 25136 12096
rect 25188 12084 25194 12096
rect 25866 12084 25872 12096
rect 25188 12056 25872 12084
rect 25188 12044 25194 12056
rect 25866 12044 25872 12056
rect 25924 12044 25930 12096
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 28810 12084 28816 12096
rect 26660 12056 28816 12084
rect 26660 12044 26666 12056
rect 28810 12044 28816 12056
rect 28868 12044 28874 12096
rect 28997 12087 29055 12093
rect 28997 12053 29009 12087
rect 29043 12084 29055 12087
rect 29178 12084 29184 12096
rect 29043 12056 29184 12084
rect 29043 12053 29055 12056
rect 28997 12047 29055 12053
rect 29178 12044 29184 12056
rect 29236 12084 29242 12096
rect 29822 12084 29828 12096
rect 29236 12056 29828 12084
rect 29236 12044 29242 12056
rect 29822 12044 29828 12056
rect 29880 12044 29886 12096
rect 2760 11994 32200 12016
rect 2760 11942 6286 11994
rect 6338 11942 6350 11994
rect 6402 11942 6414 11994
rect 6466 11942 6478 11994
rect 6530 11942 6542 11994
rect 6594 11942 13646 11994
rect 13698 11942 13710 11994
rect 13762 11942 13774 11994
rect 13826 11942 13838 11994
rect 13890 11942 13902 11994
rect 13954 11942 21006 11994
rect 21058 11942 21070 11994
rect 21122 11942 21134 11994
rect 21186 11942 21198 11994
rect 21250 11942 21262 11994
rect 21314 11942 28366 11994
rect 28418 11942 28430 11994
rect 28482 11942 28494 11994
rect 28546 11942 28558 11994
rect 28610 11942 28622 11994
rect 28674 11942 32200 11994
rect 2760 11920 32200 11942
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4396 11852 4445 11880
rect 4396 11840 4402 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4433 11843 4491 11849
rect 4706 11840 4712 11892
rect 4764 11840 4770 11892
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6822 11880 6828 11892
rect 6052 11852 6828 11880
rect 6052 11840 6058 11852
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7834 11880 7840 11892
rect 6932 11852 7840 11880
rect 4724 11753 4752 11840
rect 6932 11812 6960 11852
rect 7834 11840 7840 11852
rect 7892 11840 7898 11892
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 8076 11852 8953 11880
rect 8076 11840 8082 11852
rect 8941 11849 8953 11852
rect 8987 11880 8999 11883
rect 8987 11852 9674 11880
rect 8987 11849 8999 11852
rect 8941 11843 8999 11849
rect 5736 11784 6960 11812
rect 4709 11747 4767 11753
rect 4709 11713 4721 11747
rect 4755 11713 4767 11747
rect 4709 11707 4767 11713
rect 5736 11685 5764 11784
rect 8478 11744 8484 11756
rect 6104 11716 8484 11744
rect 6104 11688 6132 11716
rect 8478 11704 8484 11716
rect 8536 11744 8542 11756
rect 8662 11744 8668 11756
rect 8536 11716 8668 11744
rect 8536 11704 8542 11716
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11676 4583 11679
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 4571 11648 5641 11676
rect 4571 11645 4583 11648
rect 4525 11639 4583 11645
rect 5629 11645 5641 11648
rect 5675 11676 5687 11679
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 5675 11648 5733 11676
rect 5675 11645 5687 11648
rect 5629 11639 5687 11645
rect 5721 11645 5733 11648
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 6086 11636 6092 11688
rect 6144 11636 6150 11688
rect 6638 11636 6644 11688
rect 6696 11636 6702 11688
rect 9490 11636 9496 11688
rect 9548 11676 9554 11688
rect 9646 11676 9674 11852
rect 9766 11840 9772 11892
rect 9824 11840 9830 11892
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 10652 11852 12434 11880
rect 10652 11840 10658 11852
rect 9784 11753 9812 11840
rect 11333 11815 11391 11821
rect 11333 11781 11345 11815
rect 11379 11781 11391 11815
rect 12406 11812 12434 11852
rect 14090 11840 14096 11892
rect 14148 11880 14154 11892
rect 14461 11883 14519 11889
rect 14461 11880 14473 11883
rect 14148 11852 14473 11880
rect 14148 11840 14154 11852
rect 14461 11849 14473 11852
rect 14507 11880 14519 11883
rect 14829 11883 14887 11889
rect 14829 11880 14841 11883
rect 14507 11852 14841 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 14829 11849 14841 11852
rect 14875 11880 14887 11883
rect 19702 11880 19708 11892
rect 14875 11852 19708 11880
rect 14875 11849 14887 11852
rect 14829 11843 14887 11849
rect 19702 11840 19708 11852
rect 19760 11880 19766 11892
rect 20625 11883 20683 11889
rect 20625 11880 20637 11883
rect 19760 11852 20637 11880
rect 19760 11840 19766 11852
rect 20625 11849 20637 11852
rect 20671 11849 20683 11883
rect 20625 11843 20683 11849
rect 12406 11784 14964 11812
rect 11333 11775 11391 11781
rect 9769 11747 9827 11753
rect 9769 11713 9781 11747
rect 9815 11713 9827 11747
rect 9769 11707 9827 11713
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11241 11747 11299 11753
rect 11241 11713 11253 11747
rect 11287 11744 11299 11747
rect 11348 11744 11376 11775
rect 14936 11756 14964 11784
rect 15378 11772 15384 11824
rect 15436 11772 15442 11824
rect 16942 11772 16948 11824
rect 17000 11772 17006 11824
rect 17218 11772 17224 11824
rect 17276 11772 17282 11824
rect 17402 11772 17408 11824
rect 17460 11772 17466 11824
rect 19426 11772 19432 11824
rect 19484 11812 19490 11824
rect 19521 11815 19579 11821
rect 19521 11812 19533 11815
rect 19484 11784 19533 11812
rect 19484 11772 19490 11784
rect 19521 11781 19533 11784
rect 19567 11781 19579 11815
rect 19521 11775 19579 11781
rect 12894 11744 12900 11756
rect 11287 11716 11376 11744
rect 11440 11716 12900 11744
rect 11287 11713 11299 11716
rect 11241 11707 11299 11713
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 9548 11648 10333 11676
rect 9548 11636 9554 11648
rect 10321 11645 10333 11648
rect 10367 11676 10379 11679
rect 10502 11676 10508 11688
rect 10367 11648 10508 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 11072 11676 11100 11704
rect 11440 11676 11468 11716
rect 11072 11648 11468 11676
rect 11517 11679 11575 11685
rect 11517 11645 11529 11679
rect 11563 11645 11575 11679
rect 11517 11639 11575 11645
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11676 11667 11679
rect 11885 11679 11943 11685
rect 11655 11648 11836 11676
rect 11655 11645 11667 11648
rect 11609 11639 11667 11645
rect 4448 11580 6776 11608
rect 4448 11552 4476 11580
rect 4430 11500 4436 11552
rect 4488 11500 4494 11552
rect 5258 11500 5264 11552
rect 5316 11500 5322 11552
rect 5534 11500 5540 11552
rect 5592 11500 5598 11552
rect 5810 11500 5816 11552
rect 5868 11500 5874 11552
rect 6748 11549 6776 11580
rect 7742 11568 7748 11620
rect 7800 11568 7806 11620
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 8570 11608 8576 11620
rect 8251 11580 8576 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8570 11568 8576 11580
rect 8628 11568 8634 11620
rect 10520 11608 10548 11636
rect 11532 11608 11560 11639
rect 10520 11580 11560 11608
rect 11698 11568 11704 11620
rect 11756 11568 11762 11620
rect 11808 11608 11836 11648
rect 11885 11645 11897 11679
rect 11931 11676 11943 11679
rect 12066 11676 12072 11688
rect 11931 11648 12072 11676
rect 11931 11645 11943 11648
rect 11885 11639 11943 11645
rect 12066 11636 12072 11648
rect 12124 11636 12130 11688
rect 12176 11685 12204 11716
rect 12894 11704 12900 11716
rect 12952 11744 12958 11756
rect 12952 11716 14228 11744
rect 12952 11704 12958 11716
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11645 12219 11679
rect 12161 11639 12219 11645
rect 12250 11636 12256 11688
rect 12308 11636 12314 11688
rect 13538 11636 13544 11688
rect 13596 11636 13602 11688
rect 13998 11636 14004 11688
rect 14056 11676 14062 11688
rect 14200 11685 14228 11716
rect 14918 11704 14924 11756
rect 14976 11704 14982 11756
rect 17236 11744 17264 11772
rect 15488 11716 17264 11744
rect 17420 11744 17448 11772
rect 18417 11747 18475 11753
rect 18417 11744 18429 11747
rect 17420 11716 18429 11744
rect 15488 11685 15516 11716
rect 18417 11713 18429 11716
rect 18463 11713 18475 11747
rect 18417 11707 18475 11713
rect 18966 11704 18972 11756
rect 19024 11704 19030 11756
rect 19058 11704 19064 11756
rect 19116 11704 19122 11756
rect 14093 11679 14151 11685
rect 14093 11676 14105 11679
rect 14056 11648 14105 11676
rect 14056 11636 14062 11648
rect 14093 11645 14105 11648
rect 14139 11645 14151 11679
rect 14093 11639 14151 11645
rect 14185 11679 14243 11685
rect 14185 11645 14197 11679
rect 14231 11676 14243 11679
rect 15473 11679 15531 11685
rect 15473 11676 15485 11679
rect 14231 11648 15485 11676
rect 14231 11645 14243 11648
rect 14185 11639 14243 11645
rect 15473 11645 15485 11648
rect 15519 11645 15531 11679
rect 15473 11639 15531 11645
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11676 15807 11679
rect 15838 11676 15844 11688
rect 15795 11648 15844 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 11808 11580 12434 11608
rect 12406 11552 12434 11580
rect 6733 11543 6791 11549
rect 6733 11509 6745 11543
rect 6779 11540 6791 11543
rect 8386 11540 8392 11552
rect 6779 11512 8392 11540
rect 6779 11509 6791 11512
rect 6733 11503 6791 11509
rect 8386 11500 8392 11512
rect 8444 11500 8450 11552
rect 9122 11500 9128 11552
rect 9180 11500 9186 11552
rect 10594 11500 10600 11552
rect 10652 11500 10658 11552
rect 12066 11500 12072 11552
rect 12124 11500 12130 11552
rect 12342 11500 12348 11552
rect 12400 11540 12434 11552
rect 12897 11543 12955 11549
rect 12897 11540 12909 11543
rect 12400 11512 12909 11540
rect 12400 11500 12406 11512
rect 12897 11509 12909 11512
rect 12943 11509 12955 11543
rect 12897 11503 12955 11509
rect 12986 11500 12992 11552
rect 13044 11500 13050 11552
rect 15470 11500 15476 11552
rect 15528 11540 15534 11552
rect 15764 11540 15792 11639
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 18690 11636 18696 11688
rect 18748 11676 18754 11688
rect 20162 11676 20168 11688
rect 18748 11648 20168 11676
rect 18748 11636 18754 11648
rect 20162 11636 20168 11648
rect 20220 11636 20226 11688
rect 20349 11679 20407 11685
rect 20349 11645 20361 11679
rect 20395 11676 20407 11679
rect 20530 11676 20536 11688
rect 20395 11648 20536 11676
rect 20395 11645 20407 11648
rect 20349 11639 20407 11645
rect 17954 11568 17960 11620
rect 18012 11568 18018 11620
rect 18414 11568 18420 11620
rect 18472 11608 18478 11620
rect 20364 11608 20392 11639
rect 20530 11636 20536 11648
rect 20588 11636 20594 11688
rect 20640 11676 20668 11843
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 26602 11880 26608 11892
rect 23532 11852 26608 11880
rect 23532 11840 23538 11852
rect 26602 11840 26608 11852
rect 26660 11840 26666 11892
rect 27430 11840 27436 11892
rect 27488 11880 27494 11892
rect 27617 11883 27675 11889
rect 27617 11880 27629 11883
rect 27488 11852 27629 11880
rect 27488 11840 27494 11852
rect 27617 11849 27629 11852
rect 27663 11849 27675 11883
rect 27617 11843 27675 11849
rect 29730 11840 29736 11892
rect 29788 11880 29794 11892
rect 30653 11883 30711 11889
rect 30653 11880 30665 11883
rect 29788 11852 30665 11880
rect 29788 11840 29794 11852
rect 30653 11849 30665 11852
rect 30699 11849 30711 11883
rect 30653 11843 30711 11849
rect 30926 11840 30932 11892
rect 30984 11880 30990 11892
rect 31205 11883 31263 11889
rect 31205 11880 31217 11883
rect 30984 11852 31217 11880
rect 30984 11840 30990 11852
rect 31205 11849 31217 11852
rect 31251 11849 31263 11883
rect 31205 11843 31263 11849
rect 24210 11772 24216 11824
rect 24268 11812 24274 11824
rect 24486 11812 24492 11824
rect 24268 11784 24492 11812
rect 24268 11772 24274 11784
rect 24486 11772 24492 11784
rect 24544 11772 24550 11824
rect 24946 11772 24952 11824
rect 25004 11812 25010 11824
rect 27246 11812 27252 11824
rect 25004 11784 27252 11812
rect 25004 11772 25010 11784
rect 27246 11772 27252 11784
rect 27304 11812 27310 11824
rect 27304 11784 28488 11812
rect 27304 11772 27310 11784
rect 21358 11704 21364 11756
rect 21416 11744 21422 11756
rect 28460 11753 28488 11784
rect 30282 11772 30288 11824
rect 30340 11812 30346 11824
rect 30834 11812 30840 11824
rect 30340 11784 30840 11812
rect 30340 11772 30346 11784
rect 30834 11772 30840 11784
rect 30892 11772 30898 11824
rect 21637 11747 21695 11753
rect 21637 11744 21649 11747
rect 21416 11716 21649 11744
rect 21416 11704 21422 11716
rect 21637 11713 21649 11716
rect 21683 11713 21695 11747
rect 21637 11707 21695 11713
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11744 27215 11747
rect 28445 11747 28503 11753
rect 27203 11716 28120 11744
rect 27203 11713 27215 11716
rect 27157 11707 27215 11713
rect 27816 11688 27844 11716
rect 20714 11676 20720 11688
rect 20640 11648 20720 11676
rect 20714 11636 20720 11648
rect 20772 11676 20778 11688
rect 20901 11679 20959 11685
rect 20901 11676 20913 11679
rect 20772 11648 20913 11676
rect 20772 11636 20778 11648
rect 20901 11645 20913 11648
rect 20947 11676 20959 11679
rect 24213 11679 24271 11685
rect 24213 11676 24225 11679
rect 20947 11648 24225 11676
rect 20947 11645 20959 11648
rect 20901 11639 20959 11645
rect 24213 11645 24225 11648
rect 24259 11676 24271 11679
rect 24578 11676 24584 11688
rect 24259 11648 24584 11676
rect 24259 11645 24271 11648
rect 24213 11639 24271 11645
rect 24578 11636 24584 11648
rect 24636 11636 24642 11688
rect 24673 11679 24731 11685
rect 24673 11645 24685 11679
rect 24719 11676 24731 11679
rect 24854 11676 24860 11688
rect 24719 11648 24860 11676
rect 24719 11645 24731 11648
rect 24673 11639 24731 11645
rect 24854 11636 24860 11648
rect 24912 11636 24918 11688
rect 24946 11636 24952 11688
rect 25004 11636 25010 11688
rect 25130 11636 25136 11688
rect 25188 11636 25194 11688
rect 25407 11636 25413 11688
rect 25465 11636 25471 11688
rect 25866 11636 25872 11688
rect 25924 11676 25930 11688
rect 25924 11648 26924 11676
rect 25924 11636 25930 11648
rect 26896 11620 26924 11648
rect 26970 11636 26976 11688
rect 27028 11676 27034 11688
rect 27249 11679 27307 11685
rect 27028 11648 27070 11676
rect 27028 11636 27034 11648
rect 27249 11645 27261 11679
rect 27295 11645 27307 11679
rect 27249 11639 27307 11645
rect 18472 11580 20392 11608
rect 18472 11568 18478 11580
rect 25498 11568 25504 11620
rect 25556 11568 25562 11620
rect 25590 11568 25596 11620
rect 25648 11568 25654 11620
rect 25731 11611 25789 11617
rect 25731 11577 25743 11611
rect 25777 11608 25789 11611
rect 26142 11608 26148 11620
rect 25777 11580 26148 11608
rect 25777 11577 25789 11580
rect 25731 11571 25789 11577
rect 26142 11568 26148 11580
rect 26200 11568 26206 11620
rect 26237 11611 26295 11617
rect 26237 11577 26249 11611
rect 26283 11608 26295 11611
rect 26418 11608 26424 11620
rect 26283 11580 26424 11608
rect 26283 11577 26295 11580
rect 26237 11571 26295 11577
rect 26418 11568 26424 11580
rect 26476 11568 26482 11620
rect 26878 11568 26884 11620
rect 26936 11608 26942 11620
rect 27264 11608 27292 11639
rect 27430 11636 27436 11688
rect 27488 11636 27494 11688
rect 27617 11679 27675 11685
rect 27617 11645 27629 11679
rect 27663 11676 27675 11679
rect 27706 11676 27712 11688
rect 27663 11648 27712 11676
rect 27663 11645 27675 11648
rect 27617 11639 27675 11645
rect 27706 11636 27712 11648
rect 27764 11636 27770 11688
rect 27798 11636 27804 11688
rect 27856 11636 27862 11688
rect 27982 11636 27988 11688
rect 28040 11636 28046 11688
rect 28092 11685 28120 11716
rect 28445 11713 28457 11747
rect 28491 11744 28503 11747
rect 29362 11744 29368 11756
rect 28491 11716 29368 11744
rect 28491 11713 28503 11716
rect 28445 11707 28503 11713
rect 29362 11704 29368 11716
rect 29420 11704 29426 11756
rect 29454 11704 29460 11756
rect 29512 11744 29518 11756
rect 29733 11747 29791 11753
rect 29733 11744 29745 11747
rect 29512 11716 29745 11744
rect 29512 11704 29518 11716
rect 29733 11713 29745 11716
rect 29779 11713 29791 11747
rect 29733 11707 29791 11713
rect 31754 11704 31760 11756
rect 31812 11704 31818 11756
rect 28077 11679 28135 11685
rect 28077 11645 28089 11679
rect 28123 11645 28135 11679
rect 28077 11639 28135 11645
rect 28166 11636 28172 11688
rect 28224 11636 28230 11688
rect 28629 11679 28687 11685
rect 28629 11645 28641 11679
rect 28675 11645 28687 11679
rect 28629 11639 28687 11645
rect 30208 11648 30604 11676
rect 26936 11580 27292 11608
rect 27448 11608 27476 11636
rect 27893 11611 27951 11617
rect 27893 11608 27905 11611
rect 27448 11580 27905 11608
rect 26936 11568 26942 11580
rect 27893 11577 27905 11580
rect 27939 11577 27951 11611
rect 28000 11608 28028 11636
rect 28261 11611 28319 11617
rect 28261 11608 28273 11611
rect 28000 11580 28273 11608
rect 27893 11571 27951 11577
rect 28261 11577 28273 11580
rect 28307 11577 28319 11611
rect 28644 11608 28672 11639
rect 28261 11571 28319 11577
rect 28368 11580 28672 11608
rect 15528 11512 15792 11540
rect 15528 11500 15534 11512
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 16264 11512 16405 11540
rect 16264 11500 16270 11512
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 16758 11500 16764 11552
rect 16816 11540 16822 11552
rect 18782 11540 18788 11552
rect 16816 11512 18788 11540
rect 16816 11500 16822 11512
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 19153 11543 19211 11549
rect 19153 11509 19165 11543
rect 19199 11540 19211 11543
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 19199 11512 19717 11540
rect 19199 11509 19211 11512
rect 19153 11503 19211 11509
rect 19705 11509 19717 11512
rect 19751 11509 19763 11543
rect 19705 11503 19763 11509
rect 25130 11500 25136 11552
rect 25188 11500 25194 11552
rect 25222 11500 25228 11552
rect 25280 11500 25286 11552
rect 25608 11540 25636 11568
rect 26326 11540 26332 11552
rect 25608 11512 26332 11540
rect 26326 11500 26332 11512
rect 26384 11500 26390 11552
rect 27798 11500 27804 11552
rect 27856 11500 27862 11552
rect 28074 11500 28080 11552
rect 28132 11540 28138 11552
rect 28368 11540 28396 11580
rect 30208 11552 30236 11648
rect 30466 11568 30472 11620
rect 30524 11568 30530 11620
rect 30576 11608 30604 11648
rect 30669 11611 30727 11617
rect 30669 11608 30681 11611
rect 30576 11580 30681 11608
rect 30669 11577 30681 11580
rect 30715 11577 30727 11611
rect 30669 11571 30727 11577
rect 28132 11512 28396 11540
rect 28132 11500 28138 11512
rect 28902 11500 28908 11552
rect 28960 11540 28966 11552
rect 29273 11543 29331 11549
rect 29273 11540 29285 11543
rect 28960 11512 29285 11540
rect 28960 11500 28966 11512
rect 29273 11509 29285 11512
rect 29319 11509 29331 11543
rect 29273 11503 29331 11509
rect 30190 11500 30196 11552
rect 30248 11500 30254 11552
rect 30374 11500 30380 11552
rect 30432 11500 30438 11552
rect 2760 11450 32200 11472
rect 2760 11398 6946 11450
rect 6998 11398 7010 11450
rect 7062 11398 7074 11450
rect 7126 11398 7138 11450
rect 7190 11398 7202 11450
rect 7254 11398 14306 11450
rect 14358 11398 14370 11450
rect 14422 11398 14434 11450
rect 14486 11398 14498 11450
rect 14550 11398 14562 11450
rect 14614 11398 21666 11450
rect 21718 11398 21730 11450
rect 21782 11398 21794 11450
rect 21846 11398 21858 11450
rect 21910 11398 21922 11450
rect 21974 11398 29026 11450
rect 29078 11398 29090 11450
rect 29142 11398 29154 11450
rect 29206 11398 29218 11450
rect 29270 11398 29282 11450
rect 29334 11398 32200 11450
rect 2760 11376 32200 11398
rect 5626 11336 5632 11348
rect 5000 11308 5632 11336
rect 4430 11160 4436 11212
rect 4488 11160 4494 11212
rect 5000 11209 5028 11308
rect 5626 11296 5632 11308
rect 5684 11336 5690 11348
rect 6086 11336 6092 11348
rect 5684 11308 6092 11336
rect 5684 11296 5690 11308
rect 6086 11296 6092 11308
rect 6144 11296 6150 11348
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6696 11308 6745 11336
rect 6696 11296 6702 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 7742 11296 7748 11348
rect 7800 11296 7806 11348
rect 7834 11296 7840 11348
rect 7892 11296 7898 11348
rect 8386 11296 8392 11348
rect 8444 11296 8450 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 9122 11336 9128 11348
rect 8527 11308 9128 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 11977 11339 12035 11345
rect 11977 11305 11989 11339
rect 12023 11336 12035 11339
rect 12250 11336 12256 11348
rect 12023 11308 12256 11336
rect 12023 11305 12035 11308
rect 11977 11299 12035 11305
rect 12250 11296 12256 11308
rect 12308 11296 12314 11348
rect 12342 11296 12348 11348
rect 12400 11296 12406 11348
rect 12805 11339 12863 11345
rect 12805 11305 12817 11339
rect 12851 11336 12863 11339
rect 13538 11336 13544 11348
rect 12851 11308 13544 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 17954 11296 17960 11348
rect 18012 11296 18018 11348
rect 18966 11336 18972 11348
rect 18064 11308 18972 11336
rect 5258 11228 5264 11280
rect 5316 11228 5322 11280
rect 5810 11228 5816 11280
rect 5868 11228 5874 11280
rect 4985 11203 5043 11209
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 6730 11160 6736 11212
rect 6788 11200 6794 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 6788 11172 7481 11200
rect 6788 11160 6794 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 7469 11163 7527 11169
rect 7653 11203 7711 11209
rect 7653 11169 7665 11203
rect 7699 11200 7711 11203
rect 7852 11200 7880 11296
rect 8662 11228 8668 11280
rect 8720 11268 8726 11280
rect 10410 11268 10416 11280
rect 8720 11240 10416 11268
rect 8720 11228 8726 11240
rect 7699 11172 7880 11200
rect 9033 11203 9091 11209
rect 7699 11169 7711 11172
rect 7653 11163 7711 11169
rect 9033 11169 9045 11203
rect 9079 11169 9091 11203
rect 9033 11163 9091 11169
rect 3234 11092 3240 11144
rect 3292 11092 3298 11144
rect 7484 11064 7512 11163
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11101 8631 11135
rect 8573 11095 8631 11101
rect 8588 11064 8616 11095
rect 8846 11092 8852 11144
rect 8904 11092 8910 11144
rect 9048 11132 9076 11163
rect 9122 11160 9128 11212
rect 9180 11160 9186 11212
rect 9217 11203 9275 11209
rect 9217 11169 9229 11203
rect 9263 11200 9275 11203
rect 9306 11200 9312 11212
rect 9263 11172 9312 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11200 9459 11203
rect 9674 11200 9680 11212
rect 9447 11172 9680 11200
rect 9447 11169 9459 11172
rect 9401 11163 9459 11169
rect 9674 11160 9680 11172
rect 9732 11160 9738 11212
rect 9858 11160 9864 11212
rect 9916 11160 9922 11212
rect 10244 11209 10272 11240
rect 10410 11228 10416 11240
rect 10468 11228 10474 11280
rect 10505 11271 10563 11277
rect 10505 11237 10517 11271
rect 10551 11268 10563 11271
rect 10594 11268 10600 11280
rect 10551 11240 10600 11268
rect 10551 11237 10563 11240
rect 10505 11231 10563 11237
rect 10594 11228 10600 11240
rect 10652 11228 10658 11280
rect 12066 11268 12072 11280
rect 11730 11240 12072 11268
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 13633 11271 13691 11277
rect 13633 11268 13645 11271
rect 12176 11240 13645 11268
rect 10229 11203 10287 11209
rect 10229 11169 10241 11203
rect 10275 11169 10287 11203
rect 10229 11163 10287 11169
rect 9048 11104 9168 11132
rect 7484 11036 8616 11064
rect 8018 10956 8024 11008
rect 8076 10956 8082 11008
rect 8864 11005 8892 11092
rect 9140 11064 9168 11104
rect 9490 11092 9496 11144
rect 9548 11092 9554 11144
rect 9582 11092 9588 11144
rect 9640 11092 9646 11144
rect 9953 11135 10011 11141
rect 9953 11101 9965 11135
rect 9999 11132 10011 11135
rect 10042 11132 10048 11144
rect 9999 11104 10048 11132
rect 9999 11101 10011 11104
rect 9953 11095 10011 11101
rect 10042 11092 10048 11104
rect 10100 11132 10106 11144
rect 10502 11132 10508 11144
rect 10100 11104 10508 11132
rect 10100 11092 10106 11104
rect 10502 11092 10508 11104
rect 10560 11132 10566 11144
rect 12176 11132 12204 11240
rect 13633 11237 13645 11240
rect 13679 11268 13691 11271
rect 17773 11271 17831 11277
rect 13679 11240 13952 11268
rect 13679 11237 13691 11240
rect 13633 11231 13691 11237
rect 13924 11209 13952 11240
rect 17773 11237 17785 11271
rect 17819 11268 17831 11271
rect 18064 11268 18092 11308
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 21729 11339 21787 11345
rect 21729 11305 21741 11339
rect 21775 11336 21787 11339
rect 22554 11336 22560 11348
rect 21775 11308 22560 11336
rect 21775 11305 21787 11308
rect 21729 11299 21787 11305
rect 22554 11296 22560 11308
rect 22612 11296 22618 11348
rect 26418 11336 26424 11348
rect 24964 11308 26424 11336
rect 17819 11240 18092 11268
rect 17819 11237 17831 11240
rect 17773 11231 17831 11237
rect 18874 11228 18880 11280
rect 18932 11228 18938 11280
rect 19889 11271 19947 11277
rect 19889 11237 19901 11271
rect 19935 11268 19947 11271
rect 19978 11268 19984 11280
rect 19935 11240 19984 11268
rect 19935 11237 19947 11240
rect 19889 11231 19947 11237
rect 19978 11228 19984 11240
rect 20036 11228 20042 11280
rect 24964 11268 24992 11308
rect 26418 11296 26424 11308
rect 26476 11336 26482 11348
rect 28797 11339 28855 11345
rect 26476 11308 27200 11336
rect 26476 11296 26482 11308
rect 27172 11280 27200 11308
rect 28797 11305 28809 11339
rect 28843 11336 28855 11339
rect 28902 11336 28908 11348
rect 28843 11308 28908 11336
rect 28843 11305 28855 11308
rect 28797 11299 28855 11305
rect 28902 11296 28908 11308
rect 28960 11296 28966 11348
rect 29362 11336 29368 11348
rect 29104 11308 29368 11336
rect 24872 11240 24992 11268
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11200 12495 11203
rect 13909 11203 13967 11209
rect 12483 11172 12572 11200
rect 12483 11169 12495 11172
rect 12437 11163 12495 11169
rect 10560 11104 12204 11132
rect 12253 11135 12311 11141
rect 10560 11092 10566 11104
rect 12253 11101 12265 11135
rect 12299 11101 12311 11135
rect 12253 11095 12311 11101
rect 9508 11064 9536 11092
rect 9140 11036 9536 11064
rect 12268 11064 12296 11095
rect 12434 11064 12440 11076
rect 12268 11036 12440 11064
rect 12434 11024 12440 11036
rect 12492 11024 12498 11076
rect 8849 10999 8907 11005
rect 8849 10965 8861 10999
rect 8895 10965 8907 10999
rect 8849 10959 8907 10965
rect 10134 10956 10140 11008
rect 10192 10956 10198 11008
rect 11514 10956 11520 11008
rect 11572 10996 11578 11008
rect 12544 10996 12572 11172
rect 13909 11169 13921 11203
rect 13955 11169 13967 11203
rect 13909 11163 13967 11169
rect 13998 11160 14004 11212
rect 14056 11160 14062 11212
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11200 14335 11203
rect 15102 11200 15108 11212
rect 14323 11172 15108 11200
rect 14323 11169 14335 11172
rect 14277 11163 14335 11169
rect 15102 11160 15108 11172
rect 15160 11160 15166 11212
rect 16393 11203 16451 11209
rect 16393 11200 16405 11203
rect 15212 11172 16405 11200
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 12676 11104 14381 11132
rect 12676 11092 12682 11104
rect 14369 11101 14381 11104
rect 14415 11132 14427 11135
rect 14415 11104 14780 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 14752 11073 14780 11104
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 15212 11132 15240 11172
rect 16393 11169 16405 11172
rect 16439 11200 16451 11203
rect 16758 11200 16764 11212
rect 16439 11172 16764 11200
rect 16439 11169 16451 11172
rect 16393 11163 16451 11169
rect 16758 11160 16764 11172
rect 16816 11160 16822 11212
rect 18049 11203 18107 11209
rect 18049 11169 18061 11203
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 14976 11104 15240 11132
rect 14976 11092 14982 11104
rect 15562 11092 15568 11144
rect 15620 11092 15626 11144
rect 17310 11092 17316 11144
rect 17368 11092 17374 11144
rect 18064 11132 18092 11163
rect 20162 11160 20168 11212
rect 20220 11160 20226 11212
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 21637 11203 21695 11209
rect 21637 11200 21649 11203
rect 20312 11172 21649 11200
rect 20312 11160 20318 11172
rect 21637 11169 21649 11172
rect 21683 11169 21695 11203
rect 21637 11163 21695 11169
rect 22094 11160 22100 11212
rect 22152 11160 22158 11212
rect 22281 11203 22339 11209
rect 22281 11169 22293 11203
rect 22327 11200 22339 11203
rect 22370 11200 22376 11212
rect 22327 11172 22376 11200
rect 22327 11169 22339 11172
rect 22281 11163 22339 11169
rect 22370 11160 22376 11172
rect 22428 11160 22434 11212
rect 24872 11209 24900 11240
rect 25130 11228 25136 11280
rect 25188 11268 25194 11280
rect 25406 11268 25412 11280
rect 25188 11240 25412 11268
rect 25188 11228 25194 11240
rect 25406 11228 25412 11240
rect 25464 11228 25470 11280
rect 26878 11228 26884 11280
rect 26936 11228 26942 11280
rect 27154 11228 27160 11280
rect 27212 11228 27218 11280
rect 28626 11228 28632 11280
rect 28684 11268 28690 11280
rect 29104 11277 29132 11308
rect 29362 11296 29368 11308
rect 29420 11296 29426 11348
rect 30374 11296 30380 11348
rect 30432 11296 30438 11348
rect 30742 11296 30748 11348
rect 30800 11296 30806 11348
rect 30834 11296 30840 11348
rect 30892 11296 30898 11348
rect 30929 11339 30987 11345
rect 30929 11305 30941 11339
rect 30975 11336 30987 11339
rect 31294 11336 31300 11348
rect 30975 11308 31300 11336
rect 30975 11305 30987 11308
rect 30929 11299 30987 11305
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 31570 11296 31576 11348
rect 31628 11296 31634 11348
rect 28997 11271 29055 11277
rect 28997 11268 29009 11271
rect 28684 11240 29009 11268
rect 28684 11228 28690 11240
rect 28997 11237 29009 11240
rect 29043 11237 29055 11271
rect 28997 11231 29055 11237
rect 29089 11271 29147 11277
rect 29089 11237 29101 11271
rect 29135 11237 29147 11271
rect 29089 11231 29147 11237
rect 24857 11203 24915 11209
rect 24857 11169 24869 11203
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 26234 11160 26240 11212
rect 26292 11160 26298 11212
rect 26896 11200 26924 11228
rect 26973 11203 27031 11209
rect 26973 11200 26985 11203
rect 26896 11172 26985 11200
rect 26973 11169 26985 11172
rect 27019 11200 27031 11203
rect 29273 11203 29331 11209
rect 29273 11200 29285 11203
rect 27019 11172 29285 11200
rect 27019 11169 27031 11172
rect 26973 11163 27031 11169
rect 29273 11169 29285 11172
rect 29319 11169 29331 11203
rect 29273 11163 29331 11169
rect 29730 11160 29736 11212
rect 29788 11200 29794 11212
rect 30009 11203 30067 11209
rect 30009 11200 30021 11203
rect 29788 11172 30021 11200
rect 29788 11160 29794 11172
rect 30009 11169 30021 11172
rect 30055 11169 30067 11203
rect 30009 11163 30067 11169
rect 30098 11160 30104 11212
rect 30156 11160 30162 11212
rect 30282 11160 30288 11212
rect 30340 11160 30346 11212
rect 30392 11200 30420 11296
rect 30852 11268 30880 11296
rect 30852 11240 31064 11268
rect 31036 11209 31064 11240
rect 30837 11203 30895 11209
rect 30837 11200 30849 11203
rect 30392 11172 30849 11200
rect 30837 11169 30849 11172
rect 30883 11169 30895 11203
rect 30837 11163 30895 11169
rect 31021 11203 31079 11209
rect 31021 11169 31033 11203
rect 31067 11169 31079 11203
rect 31021 11163 31079 11169
rect 31386 11160 31392 11212
rect 31444 11160 31450 11212
rect 31662 11160 31668 11212
rect 31720 11160 31726 11212
rect 19242 11132 19248 11144
rect 18064 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 20806 11092 20812 11144
rect 20864 11132 20870 11144
rect 21821 11135 21879 11141
rect 21821 11132 21833 11135
rect 20864 11104 21833 11132
rect 20864 11092 20870 11104
rect 21821 11101 21833 11104
rect 21867 11101 21879 11135
rect 21821 11095 21879 11101
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 25130 11092 25136 11144
rect 25188 11092 25194 11144
rect 26605 11135 26663 11141
rect 26605 11101 26617 11135
rect 26651 11132 26663 11135
rect 26697 11135 26755 11141
rect 26697 11132 26709 11135
rect 26651 11104 26709 11132
rect 26651 11101 26663 11104
rect 26605 11095 26663 11101
rect 26697 11101 26709 11104
rect 26743 11101 26755 11135
rect 26697 11095 26755 11101
rect 27062 11092 27068 11144
rect 27120 11132 27126 11144
rect 28169 11135 28227 11141
rect 28169 11132 28181 11135
rect 27120 11104 28181 11132
rect 27120 11092 27126 11104
rect 28169 11101 28181 11104
rect 28215 11101 28227 11135
rect 28169 11095 28227 11101
rect 13725 11067 13783 11073
rect 13725 11064 13737 11067
rect 13504 11036 13737 11064
rect 13504 11024 13510 11036
rect 13725 11033 13737 11036
rect 13771 11033 13783 11067
rect 13725 11027 13783 11033
rect 14737 11067 14795 11073
rect 14737 11033 14749 11067
rect 14783 11064 14795 11067
rect 16850 11064 16856 11076
rect 14783 11036 16856 11064
rect 14783 11033 14795 11036
rect 14737 11027 14795 11033
rect 16850 11024 16856 11036
rect 16908 11024 16914 11076
rect 18414 11024 18420 11076
rect 18472 11024 18478 11076
rect 21269 11067 21327 11073
rect 21269 11033 21281 11067
rect 21315 11064 21327 11067
rect 21358 11064 21364 11076
rect 21315 11036 21364 11064
rect 21315 11033 21327 11036
rect 21269 11027 21327 11033
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 29457 11067 29515 11073
rect 29457 11064 29469 11067
rect 27172 11036 29469 11064
rect 11572 10968 12572 10996
rect 11572 10956 11578 10968
rect 16666 10956 16672 11008
rect 16724 10996 16730 11008
rect 16761 10999 16819 11005
rect 16761 10996 16773 10999
rect 16724 10968 16773 10996
rect 16724 10956 16730 10968
rect 16761 10965 16773 10968
rect 16807 10965 16819 10999
rect 16761 10959 16819 10965
rect 18782 10956 18788 11008
rect 18840 10996 18846 11008
rect 24394 10996 24400 11008
rect 18840 10968 24400 10996
rect 18840 10956 18846 10968
rect 24394 10956 24400 10968
rect 24452 10956 24458 11008
rect 25314 10956 25320 11008
rect 25372 10996 25378 11008
rect 27172 10996 27200 11036
rect 29457 11033 29469 11036
rect 29503 11033 29515 11067
rect 29457 11027 29515 11033
rect 30285 11067 30343 11073
rect 30285 11033 30297 11067
rect 30331 11064 30343 11067
rect 31478 11064 31484 11076
rect 30331 11036 31484 11064
rect 30331 11033 30343 11036
rect 30285 11027 30343 11033
rect 31478 11024 31484 11036
rect 31536 11024 31542 11076
rect 25372 10968 27200 10996
rect 27617 10999 27675 11005
rect 25372 10956 25378 10968
rect 27617 10965 27629 10999
rect 27663 10996 27675 10999
rect 27706 10996 27712 11008
rect 27663 10968 27712 10996
rect 27663 10965 27675 10968
rect 27617 10959 27675 10965
rect 27706 10956 27712 10968
rect 27764 10956 27770 11008
rect 28629 10999 28687 11005
rect 28629 10965 28641 10999
rect 28675 10996 28687 10999
rect 28718 10996 28724 11008
rect 28675 10968 28724 10996
rect 28675 10965 28687 10968
rect 28629 10959 28687 10965
rect 28718 10956 28724 10968
rect 28776 10956 28782 11008
rect 28810 10956 28816 11008
rect 28868 10956 28874 11008
rect 31018 10956 31024 11008
rect 31076 10996 31082 11008
rect 31205 10999 31263 11005
rect 31205 10996 31217 10999
rect 31076 10968 31217 10996
rect 31076 10956 31082 10968
rect 31205 10965 31217 10968
rect 31251 10965 31263 10999
rect 31205 10959 31263 10965
rect 2760 10906 32200 10928
rect 2760 10854 6286 10906
rect 6338 10854 6350 10906
rect 6402 10854 6414 10906
rect 6466 10854 6478 10906
rect 6530 10854 6542 10906
rect 6594 10854 13646 10906
rect 13698 10854 13710 10906
rect 13762 10854 13774 10906
rect 13826 10854 13838 10906
rect 13890 10854 13902 10906
rect 13954 10854 21006 10906
rect 21058 10854 21070 10906
rect 21122 10854 21134 10906
rect 21186 10854 21198 10906
rect 21250 10854 21262 10906
rect 21314 10854 28366 10906
rect 28418 10854 28430 10906
rect 28482 10854 28494 10906
rect 28546 10854 28558 10906
rect 28610 10854 28622 10906
rect 28674 10854 32200 10906
rect 2760 10832 32200 10854
rect 5902 10752 5908 10804
rect 5960 10792 5966 10804
rect 6362 10792 6368 10804
rect 5960 10764 6368 10792
rect 5960 10752 5966 10764
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 8570 10752 8576 10804
rect 8628 10752 8634 10804
rect 12986 10792 12992 10804
rect 12360 10764 12992 10792
rect 5920 10724 5948 10752
rect 5644 10696 5948 10724
rect 6181 10727 6239 10733
rect 5644 10665 5672 10696
rect 6181 10693 6193 10727
rect 6227 10724 6239 10727
rect 6227 10696 6868 10724
rect 6227 10693 6239 10696
rect 6181 10687 6239 10693
rect 5629 10659 5687 10665
rect 5629 10625 5641 10659
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10656 5779 10659
rect 5994 10656 6000 10668
rect 5767 10628 6000 10656
rect 5767 10625 5779 10628
rect 5721 10619 5779 10625
rect 5994 10616 6000 10628
rect 6052 10616 6058 10668
rect 6840 10665 6868 10696
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 8018 10616 8024 10668
rect 8076 10616 8082 10668
rect 10134 10616 10140 10668
rect 10192 10616 10198 10668
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 12161 10659 12219 10665
rect 12161 10625 12173 10659
rect 12207 10656 12219 10659
rect 12360 10656 12388 10764
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13998 10792 14004 10804
rect 13228 10764 14004 10792
rect 13228 10752 13234 10764
rect 13998 10752 14004 10764
rect 14056 10752 14062 10804
rect 18874 10752 18880 10804
rect 18932 10792 18938 10804
rect 18969 10795 19027 10801
rect 18969 10792 18981 10795
rect 18932 10764 18981 10792
rect 18932 10752 18938 10764
rect 18969 10761 18981 10764
rect 19015 10761 19027 10795
rect 18969 10755 19027 10761
rect 20254 10752 20260 10804
rect 20312 10752 20318 10804
rect 20714 10752 20720 10804
rect 20772 10752 20778 10804
rect 20898 10752 20904 10804
rect 20956 10792 20962 10804
rect 23569 10795 23627 10801
rect 23569 10792 23581 10795
rect 20956 10764 23581 10792
rect 20956 10752 20962 10764
rect 23569 10761 23581 10764
rect 23615 10761 23627 10795
rect 23569 10755 23627 10761
rect 23750 10752 23756 10804
rect 23808 10752 23814 10804
rect 25130 10752 25136 10804
rect 25188 10792 25194 10804
rect 25225 10795 25283 10801
rect 25225 10792 25237 10795
rect 25188 10764 25237 10792
rect 25188 10752 25194 10764
rect 25225 10761 25237 10764
rect 25271 10761 25283 10795
rect 25225 10755 25283 10761
rect 26053 10795 26111 10801
rect 26053 10761 26065 10795
rect 26099 10792 26111 10795
rect 27062 10792 27068 10804
rect 26099 10764 27068 10792
rect 26099 10761 26111 10764
rect 26053 10755 26111 10761
rect 27062 10752 27068 10764
rect 27120 10752 27126 10804
rect 29273 10795 29331 10801
rect 29273 10761 29285 10795
rect 29319 10792 29331 10795
rect 29454 10792 29460 10804
rect 29319 10764 29460 10792
rect 29319 10761 29331 10764
rect 29273 10755 29331 10761
rect 29454 10752 29460 10764
rect 29512 10792 29518 10804
rect 30098 10792 30104 10804
rect 29512 10764 30104 10792
rect 29512 10752 29518 10764
rect 30098 10752 30104 10764
rect 30156 10752 30162 10804
rect 30190 10752 30196 10804
rect 30248 10752 30254 10804
rect 30282 10752 30288 10804
rect 30340 10752 30346 10804
rect 14829 10727 14887 10733
rect 14829 10693 14841 10727
rect 14875 10724 14887 10727
rect 15654 10724 15660 10736
rect 14875 10696 15660 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 15654 10684 15660 10696
rect 15712 10684 15718 10736
rect 18785 10727 18843 10733
rect 18785 10693 18797 10727
rect 18831 10724 18843 10727
rect 19334 10724 19340 10736
rect 18831 10696 19340 10724
rect 18831 10693 18843 10696
rect 18785 10687 18843 10693
rect 19334 10684 19340 10696
rect 19392 10724 19398 10736
rect 20272 10724 20300 10752
rect 22922 10724 22928 10736
rect 19392 10696 20300 10724
rect 21008 10696 22928 10724
rect 19392 10684 19398 10696
rect 12207 10628 12388 10656
rect 12437 10659 12495 10665
rect 12207 10625 12219 10628
rect 12161 10619 12219 10625
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12526 10656 12532 10668
rect 12483 10628 12532 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12526 10616 12532 10628
rect 12584 10656 12590 10668
rect 13357 10659 13415 10665
rect 12584 10628 13124 10656
rect 12584 10616 12590 10628
rect 13096 10600 13124 10628
rect 13357 10625 13369 10659
rect 13403 10656 13415 10659
rect 13446 10656 13452 10668
rect 13403 10628 13452 10656
rect 13403 10625 13415 10628
rect 13357 10619 13415 10625
rect 13446 10616 13452 10628
rect 13504 10616 13510 10668
rect 15010 10656 15016 10668
rect 14660 10628 15016 10656
rect 14660 10600 14688 10628
rect 15010 10616 15016 10628
rect 15068 10656 15074 10668
rect 16298 10656 16304 10668
rect 15068 10628 16304 10656
rect 15068 10616 15074 10628
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 16577 10659 16635 10665
rect 16577 10625 16589 10659
rect 16623 10656 16635 10659
rect 16666 10656 16672 10668
rect 16623 10628 16672 10656
rect 16623 10625 16635 10628
rect 16577 10619 16635 10625
rect 16666 10616 16672 10628
rect 16724 10616 16730 10668
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10656 18107 10659
rect 18141 10659 18199 10665
rect 18141 10656 18153 10659
rect 18095 10628 18153 10656
rect 18095 10625 18107 10628
rect 18049 10619 18107 10625
rect 18141 10625 18153 10628
rect 18187 10625 18199 10659
rect 19242 10656 19248 10668
rect 18141 10619 18199 10625
rect 18892 10628 19248 10656
rect 4338 10548 4344 10600
rect 4396 10588 4402 10600
rect 4617 10591 4675 10597
rect 4617 10588 4629 10591
rect 4396 10560 4629 10588
rect 4396 10548 4402 10560
rect 4617 10557 4629 10560
rect 4663 10557 4675 10591
rect 4617 10551 4675 10557
rect 12713 10591 12771 10597
rect 12713 10557 12725 10591
rect 12759 10557 12771 10591
rect 12713 10551 12771 10557
rect 5261 10523 5319 10529
rect 5261 10489 5273 10523
rect 5307 10520 5319 10523
rect 5813 10523 5871 10529
rect 5813 10520 5825 10523
rect 5307 10492 5825 10520
rect 5307 10489 5319 10492
rect 5261 10483 5319 10489
rect 5813 10489 5825 10492
rect 5859 10489 5871 10523
rect 5813 10483 5871 10489
rect 9674 10480 9680 10532
rect 9732 10480 9738 10532
rect 11730 10492 12434 10520
rect 6270 10412 6276 10464
rect 6328 10412 6334 10464
rect 8662 10412 8668 10464
rect 8720 10412 8726 10464
rect 10689 10455 10747 10461
rect 10689 10421 10701 10455
rect 10735 10452 10747 10455
rect 11514 10452 11520 10464
rect 10735 10424 11520 10452
rect 10735 10421 10747 10424
rect 10689 10415 10747 10421
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 12406 10452 12434 10492
rect 12728 10464 12756 10551
rect 13078 10548 13084 10600
rect 13136 10548 13142 10600
rect 14642 10548 14648 10600
rect 14700 10548 14706 10600
rect 15194 10548 15200 10600
rect 15252 10548 15258 10600
rect 18892 10597 18920 10628
rect 19242 10616 19248 10628
rect 19300 10616 19306 10668
rect 21008 10597 21036 10696
rect 22922 10684 22928 10696
rect 22980 10684 22986 10736
rect 23109 10727 23167 10733
rect 23109 10693 23121 10727
rect 23155 10693 23167 10727
rect 23109 10687 23167 10693
rect 29089 10727 29147 10733
rect 29089 10693 29101 10727
rect 29135 10724 29147 10727
rect 30208 10724 30236 10752
rect 29135 10696 30236 10724
rect 29135 10693 29147 10696
rect 29089 10687 29147 10693
rect 15473 10591 15531 10597
rect 15473 10557 15485 10591
rect 15519 10588 15531 10591
rect 18877 10591 18935 10597
rect 15519 10560 15976 10588
rect 15519 10557 15531 10560
rect 15473 10551 15531 10557
rect 14090 10480 14096 10532
rect 14148 10480 14154 10532
rect 15562 10520 15568 10532
rect 14936 10492 15568 10520
rect 12621 10455 12679 10461
rect 12621 10452 12633 10455
rect 12406 10424 12633 10452
rect 12621 10421 12633 10424
rect 12667 10421 12679 10455
rect 12621 10415 12679 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 14936 10452 14964 10492
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 15948 10464 15976 10560
rect 18877 10557 18889 10591
rect 18923 10557 18935 10591
rect 20993 10591 21051 10597
rect 20993 10588 21005 10591
rect 18877 10551 18935 10557
rect 19260 10560 21005 10588
rect 18414 10520 18420 10532
rect 17802 10492 18420 10520
rect 18414 10480 18420 10492
rect 18472 10480 18478 10532
rect 19260 10464 19288 10560
rect 20993 10557 21005 10560
rect 21039 10557 21051 10591
rect 22189 10591 22247 10597
rect 22189 10588 22201 10591
rect 20993 10551 21051 10557
rect 21376 10560 22201 10588
rect 20714 10480 20720 10532
rect 20772 10520 20778 10532
rect 21376 10520 21404 10560
rect 22189 10557 22201 10560
rect 22235 10557 22247 10591
rect 22189 10551 22247 10557
rect 22278 10548 22284 10600
rect 22336 10548 22342 10600
rect 20772 10492 21404 10520
rect 20772 10480 20778 10492
rect 21450 10480 21456 10532
rect 21508 10480 21514 10532
rect 22002 10480 22008 10532
rect 22060 10520 22066 10532
rect 23124 10520 23152 10687
rect 25222 10616 25228 10668
rect 25280 10656 25286 10668
rect 25777 10659 25835 10665
rect 25777 10656 25789 10659
rect 25280 10628 25789 10656
rect 25280 10616 25286 10628
rect 25777 10625 25789 10628
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 27154 10616 27160 10668
rect 27212 10656 27218 10668
rect 27801 10659 27859 10665
rect 27801 10656 27813 10659
rect 27212 10628 27813 10656
rect 27212 10616 27218 10628
rect 27801 10625 27813 10628
rect 27847 10656 27859 10659
rect 29362 10656 29368 10668
rect 27847 10628 29368 10656
rect 27847 10625 27859 10628
rect 27801 10619 27859 10625
rect 29362 10616 29368 10628
rect 29420 10616 29426 10668
rect 29472 10628 30788 10656
rect 23198 10548 23204 10600
rect 23256 10588 23262 10600
rect 23753 10591 23811 10597
rect 23753 10588 23765 10591
rect 23256 10560 23765 10588
rect 23256 10548 23262 10560
rect 23753 10557 23765 10560
rect 23799 10557 23811 10591
rect 23753 10551 23811 10557
rect 23937 10591 23995 10597
rect 23937 10557 23949 10591
rect 23983 10557 23995 10591
rect 23937 10551 23995 10557
rect 24029 10591 24087 10597
rect 24029 10557 24041 10591
rect 24075 10588 24087 10591
rect 24118 10588 24124 10600
rect 24075 10560 24124 10588
rect 24075 10557 24087 10560
rect 24029 10551 24087 10557
rect 22060 10492 23152 10520
rect 23477 10523 23535 10529
rect 22060 10480 22066 10492
rect 23477 10489 23489 10523
rect 23523 10520 23535 10523
rect 23658 10520 23664 10532
rect 23523 10492 23664 10520
rect 23523 10489 23535 10492
rect 23477 10483 23535 10489
rect 23658 10480 23664 10492
rect 23716 10480 23722 10532
rect 23952 10520 23980 10551
rect 24118 10548 24124 10560
rect 24176 10548 24182 10600
rect 24213 10591 24271 10597
rect 24213 10557 24225 10591
rect 24259 10557 24271 10591
rect 24213 10551 24271 10557
rect 24228 10520 24256 10551
rect 26418 10548 26424 10600
rect 26476 10548 26482 10600
rect 28537 10591 28595 10597
rect 28537 10557 28549 10591
rect 28583 10588 28595 10591
rect 28718 10588 28724 10600
rect 28583 10560 28724 10588
rect 28583 10557 28595 10560
rect 28537 10551 28595 10557
rect 28718 10548 28724 10560
rect 28776 10548 28782 10600
rect 29472 10588 29500 10628
rect 30760 10600 30788 10628
rect 29380 10560 29500 10588
rect 24854 10520 24860 10532
rect 23952 10492 24164 10520
rect 24228 10492 24860 10520
rect 12768 10424 14964 10452
rect 15013 10455 15071 10461
rect 12768 10412 12774 10424
rect 15013 10421 15025 10455
rect 15059 10452 15071 10455
rect 15286 10452 15292 10464
rect 15059 10424 15292 10452
rect 15059 10421 15071 10424
rect 15013 10415 15071 10421
rect 15286 10412 15292 10424
rect 15344 10412 15350 10464
rect 15378 10412 15384 10464
rect 15436 10412 15442 10464
rect 15930 10412 15936 10464
rect 15988 10412 15994 10464
rect 19242 10412 19248 10464
rect 19300 10412 19306 10464
rect 20990 10412 20996 10464
rect 21048 10452 21054 10464
rect 21085 10455 21143 10461
rect 21085 10452 21097 10455
rect 21048 10424 21097 10452
rect 21048 10412 21054 10424
rect 21085 10421 21097 10424
rect 21131 10421 21143 10455
rect 21085 10415 21143 10421
rect 22370 10412 22376 10464
rect 22428 10452 22434 10464
rect 22465 10455 22523 10461
rect 22465 10452 22477 10455
rect 22428 10424 22477 10452
rect 22428 10412 22434 10424
rect 22465 10421 22477 10424
rect 22511 10421 22523 10455
rect 22465 10415 22523 10421
rect 23014 10412 23020 10464
rect 23072 10412 23078 10464
rect 24136 10461 24164 10492
rect 24854 10480 24860 10492
rect 24912 10480 24918 10532
rect 27525 10523 27583 10529
rect 27525 10489 27537 10523
rect 27571 10520 27583 10523
rect 27893 10523 27951 10529
rect 27893 10520 27905 10523
rect 27571 10492 27905 10520
rect 27571 10489 27583 10492
rect 27525 10483 27583 10489
rect 27893 10489 27905 10492
rect 27939 10489 27951 10523
rect 29380 10520 29408 10560
rect 29546 10548 29552 10600
rect 29604 10548 29610 10600
rect 30742 10548 30748 10600
rect 30800 10548 30806 10600
rect 30926 10548 30932 10600
rect 30984 10548 30990 10600
rect 31205 10591 31263 10597
rect 31205 10557 31217 10591
rect 31251 10557 31263 10591
rect 31205 10551 31263 10557
rect 27893 10483 27951 10489
rect 28000 10492 29408 10520
rect 29457 10523 29515 10529
rect 24121 10455 24179 10461
rect 24121 10421 24133 10455
rect 24167 10452 24179 10455
rect 24302 10452 24308 10464
rect 24167 10424 24308 10452
rect 24167 10421 24179 10424
rect 24121 10415 24179 10421
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 24394 10412 24400 10464
rect 24452 10452 24458 10464
rect 28000 10452 28028 10492
rect 29457 10489 29469 10523
rect 29503 10520 29515 10523
rect 29638 10520 29644 10532
rect 29503 10492 29644 10520
rect 29503 10489 29515 10492
rect 29457 10483 29515 10489
rect 29638 10480 29644 10492
rect 29696 10520 29702 10532
rect 30282 10520 30288 10532
rect 29696 10492 30288 10520
rect 29696 10480 29702 10492
rect 30282 10480 30288 10492
rect 30340 10480 30346 10532
rect 30760 10520 30788 10548
rect 31220 10520 31248 10551
rect 30760 10492 31248 10520
rect 31386 10480 31392 10532
rect 31444 10520 31450 10532
rect 31481 10523 31539 10529
rect 31481 10520 31493 10523
rect 31444 10492 31493 10520
rect 31444 10480 31450 10492
rect 31481 10489 31493 10492
rect 31527 10489 31539 10523
rect 31481 10483 31539 10489
rect 24452 10424 28028 10452
rect 29257 10455 29315 10461
rect 24452 10412 24458 10424
rect 29257 10421 29269 10455
rect 29303 10452 29315 10455
rect 29730 10452 29736 10464
rect 29303 10424 29736 10452
rect 29303 10421 29315 10424
rect 29257 10415 29315 10421
rect 29730 10412 29736 10424
rect 29788 10412 29794 10464
rect 29914 10412 29920 10464
rect 29972 10452 29978 10464
rect 30193 10455 30251 10461
rect 30193 10452 30205 10455
rect 29972 10424 30205 10452
rect 29972 10412 29978 10424
rect 30193 10421 30205 10424
rect 30239 10421 30251 10455
rect 30193 10415 30251 10421
rect 2760 10362 32200 10384
rect 2760 10310 6946 10362
rect 6998 10310 7010 10362
rect 7062 10310 7074 10362
rect 7126 10310 7138 10362
rect 7190 10310 7202 10362
rect 7254 10310 14306 10362
rect 14358 10310 14370 10362
rect 14422 10310 14434 10362
rect 14486 10310 14498 10362
rect 14550 10310 14562 10362
rect 14614 10310 21666 10362
rect 21718 10310 21730 10362
rect 21782 10310 21794 10362
rect 21846 10310 21858 10362
rect 21910 10310 21922 10362
rect 21974 10310 29026 10362
rect 29078 10310 29090 10362
rect 29142 10310 29154 10362
rect 29206 10310 29218 10362
rect 29270 10310 29282 10362
rect 29334 10310 32200 10362
rect 2760 10288 32200 10310
rect 6270 10208 6276 10260
rect 6328 10208 6334 10260
rect 6362 10208 6368 10260
rect 6420 10208 6426 10260
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 9364 10220 9505 10248
rect 9364 10208 9370 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 9732 10220 10149 10248
rect 9732 10208 9738 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 10137 10211 10195 10217
rect 10502 10208 10508 10260
rect 10560 10208 10566 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 12897 10251 12955 10257
rect 12897 10248 12909 10251
rect 12492 10220 12909 10248
rect 12492 10208 12498 10220
rect 12897 10217 12909 10220
rect 12943 10217 12955 10251
rect 12897 10211 12955 10217
rect 14090 10208 14096 10260
rect 14148 10208 14154 10260
rect 14553 10251 14611 10257
rect 14553 10217 14565 10251
rect 14599 10248 14611 10251
rect 14918 10248 14924 10260
rect 14599 10220 14924 10248
rect 14599 10217 14611 10220
rect 14553 10211 14611 10217
rect 5534 10180 5540 10192
rect 5382 10152 5540 10180
rect 5534 10140 5540 10152
rect 5592 10140 5598 10192
rect 5813 10183 5871 10189
rect 5813 10149 5825 10183
rect 5859 10180 5871 10183
rect 6288 10180 6316 10208
rect 5859 10152 6316 10180
rect 5859 10149 5871 10152
rect 5813 10143 5871 10149
rect 9766 10140 9772 10192
rect 9824 10180 9830 10192
rect 9861 10183 9919 10189
rect 9861 10180 9873 10183
rect 9824 10152 9873 10180
rect 9824 10140 9830 10152
rect 9861 10149 9873 10152
rect 9907 10149 9919 10183
rect 9861 10143 9919 10149
rect 3050 10072 3056 10124
rect 3108 10072 3114 10124
rect 10229 10115 10287 10121
rect 10229 10081 10241 10115
rect 10275 10112 10287 10115
rect 12710 10112 12716 10124
rect 10275 10084 12716 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 12710 10072 12716 10084
rect 12768 10072 12774 10124
rect 14001 10115 14059 10121
rect 14001 10081 14013 10115
rect 14047 10112 14059 10115
rect 14568 10112 14596 10211
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 16853 10251 16911 10257
rect 15620 10220 16712 10248
rect 15620 10208 15626 10220
rect 16577 10183 16635 10189
rect 16577 10180 16589 10183
rect 16146 10152 16589 10180
rect 16577 10149 16589 10152
rect 16623 10149 16635 10183
rect 16577 10143 16635 10149
rect 16684 10121 16712 10220
rect 16853 10217 16865 10251
rect 16899 10248 16911 10251
rect 17310 10248 17316 10260
rect 16899 10220 17316 10248
rect 16899 10217 16911 10220
rect 16853 10211 16911 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18414 10208 18420 10260
rect 18472 10208 18478 10260
rect 18782 10208 18788 10260
rect 18840 10208 18846 10260
rect 19334 10208 19340 10260
rect 19392 10208 19398 10260
rect 20533 10251 20591 10257
rect 20533 10217 20545 10251
rect 20579 10248 20591 10251
rect 22278 10248 22284 10260
rect 20579 10220 22284 10248
rect 20579 10217 20591 10220
rect 20533 10211 20591 10217
rect 22278 10208 22284 10220
rect 22336 10208 22342 10260
rect 22741 10251 22799 10257
rect 22741 10217 22753 10251
rect 22787 10248 22799 10251
rect 24213 10251 24271 10257
rect 24213 10248 24225 10251
rect 22787 10220 24225 10248
rect 22787 10217 22799 10220
rect 22741 10211 22799 10217
rect 24213 10217 24225 10220
rect 24259 10217 24271 10251
rect 25777 10251 25835 10257
rect 24213 10211 24271 10217
rect 24320 10220 24624 10248
rect 17221 10183 17279 10189
rect 17221 10149 17233 10183
rect 17267 10180 17279 10183
rect 19352 10180 19380 10208
rect 17267 10152 19380 10180
rect 17267 10149 17279 10152
rect 17221 10143 17279 10149
rect 20990 10140 20996 10192
rect 21048 10140 21054 10192
rect 22005 10183 22063 10189
rect 22005 10149 22017 10183
rect 22051 10180 22063 10183
rect 23477 10183 23535 10189
rect 23477 10180 23489 10183
rect 22051 10152 23489 10180
rect 22051 10149 22063 10152
rect 22005 10143 22063 10149
rect 23477 10149 23489 10152
rect 23523 10149 23535 10183
rect 23477 10143 23535 10149
rect 24118 10140 24124 10192
rect 24176 10180 24182 10192
rect 24320 10180 24348 10220
rect 24596 10189 24624 10220
rect 25777 10217 25789 10251
rect 25823 10248 25835 10251
rect 26234 10248 26240 10260
rect 25823 10220 26240 10248
rect 25823 10217 25835 10220
rect 25777 10211 25835 10217
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 26418 10208 26424 10260
rect 26476 10208 26482 10260
rect 27249 10251 27307 10257
rect 27249 10217 27261 10251
rect 27295 10248 27307 10251
rect 28074 10248 28080 10260
rect 27295 10220 28080 10248
rect 27295 10217 27307 10220
rect 27249 10211 27307 10217
rect 28074 10208 28080 10220
rect 28132 10208 28138 10260
rect 29273 10251 29331 10257
rect 29273 10217 29285 10251
rect 29319 10248 29331 10251
rect 29546 10248 29552 10260
rect 29319 10220 29552 10248
rect 29319 10217 29331 10220
rect 29273 10211 29331 10217
rect 29546 10208 29552 10220
rect 29604 10208 29610 10260
rect 29914 10208 29920 10260
rect 29972 10208 29978 10260
rect 30926 10208 30932 10260
rect 30984 10248 30990 10260
rect 31113 10251 31171 10257
rect 31113 10248 31125 10251
rect 30984 10220 31125 10248
rect 30984 10208 30990 10220
rect 31113 10217 31125 10220
rect 31159 10217 31171 10251
rect 31113 10211 31171 10217
rect 24176 10152 24348 10180
rect 24381 10183 24439 10189
rect 24176 10140 24182 10152
rect 24381 10149 24393 10183
rect 24427 10180 24439 10183
rect 24581 10183 24639 10189
rect 24427 10152 24532 10180
rect 24427 10149 24439 10152
rect 24381 10143 24439 10149
rect 14047 10084 14596 10112
rect 16669 10115 16727 10121
rect 14047 10081 14059 10084
rect 14001 10075 14059 10081
rect 16669 10081 16681 10115
rect 16715 10112 16727 10115
rect 16758 10112 16764 10124
rect 16715 10084 16764 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 16758 10072 16764 10084
rect 16816 10072 16822 10124
rect 18509 10115 18567 10121
rect 18509 10081 18521 10115
rect 18555 10112 18567 10115
rect 18782 10112 18788 10124
rect 18555 10084 18788 10112
rect 18555 10081 18567 10084
rect 18509 10075 18567 10081
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 6086 10004 6092 10056
rect 6144 10004 6150 10056
rect 14642 10004 14648 10056
rect 14700 10004 14706 10056
rect 14918 10004 14924 10056
rect 14976 10004 14982 10056
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 16393 10047 16451 10053
rect 15436 10016 16344 10044
rect 15436 10004 15442 10016
rect 16316 9976 16344 10016
rect 16393 10013 16405 10047
rect 16439 10044 16451 10047
rect 16574 10044 16580 10056
rect 16439 10016 16580 10044
rect 16439 10013 16451 10016
rect 16393 10007 16451 10013
rect 16574 10004 16580 10016
rect 16632 10004 16638 10056
rect 17313 10047 17371 10053
rect 17313 10013 17325 10047
rect 17359 10013 17371 10047
rect 17313 10007 17371 10013
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 19242 10044 19248 10056
rect 17543 10016 18000 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 17328 9976 17356 10007
rect 16316 9948 17356 9976
rect 17972 9920 18000 10016
rect 18524 10016 19248 10044
rect 18524 9920 18552 10016
rect 19242 10004 19248 10016
rect 19300 10044 19306 10056
rect 19812 10044 19840 10075
rect 23382 10072 23388 10124
rect 23440 10112 23446 10124
rect 24504 10112 24532 10152
rect 24581 10149 24593 10183
rect 24627 10180 24639 10183
rect 25498 10180 25504 10192
rect 24627 10152 25504 10180
rect 24627 10149 24639 10152
rect 24581 10143 24639 10149
rect 25498 10140 25504 10152
rect 25556 10140 25562 10192
rect 27614 10180 27620 10192
rect 26988 10152 27620 10180
rect 24854 10112 24860 10124
rect 23440 10084 24860 10112
rect 23440 10072 23446 10084
rect 24854 10072 24860 10084
rect 24912 10112 24918 10124
rect 25406 10112 25412 10124
rect 24912 10084 25412 10112
rect 24912 10072 24918 10084
rect 25406 10072 25412 10084
rect 25464 10072 25470 10124
rect 25685 10115 25743 10121
rect 25685 10081 25697 10115
rect 25731 10112 25743 10115
rect 25774 10112 25780 10124
rect 25731 10084 25780 10112
rect 25731 10081 25743 10084
rect 25685 10075 25743 10081
rect 25774 10072 25780 10084
rect 25832 10112 25838 10124
rect 26329 10115 26387 10121
rect 26329 10112 26341 10115
rect 25832 10084 26341 10112
rect 25832 10072 25838 10084
rect 26329 10081 26341 10084
rect 26375 10081 26387 10115
rect 26329 10075 26387 10081
rect 26878 10072 26884 10124
rect 26936 10072 26942 10124
rect 26988 10121 27016 10152
rect 27614 10140 27620 10152
rect 27672 10140 27678 10192
rect 27798 10140 27804 10192
rect 27856 10180 27862 10192
rect 27985 10183 28043 10189
rect 27985 10180 27997 10183
rect 27856 10152 27997 10180
rect 27856 10140 27862 10152
rect 27985 10149 27997 10152
rect 28031 10149 28043 10183
rect 27985 10143 28043 10149
rect 28166 10140 28172 10192
rect 28224 10180 28230 10192
rect 29641 10183 29699 10189
rect 28224 10152 28304 10180
rect 28224 10140 28230 10152
rect 26973 10115 27031 10121
rect 26973 10081 26985 10115
rect 27019 10081 27031 10115
rect 26973 10075 27031 10081
rect 27065 10115 27123 10121
rect 27065 10081 27077 10115
rect 27111 10112 27123 10115
rect 27246 10112 27252 10124
rect 27111 10084 27252 10112
rect 27111 10081 27123 10084
rect 27065 10075 27123 10081
rect 27246 10072 27252 10084
rect 27304 10072 27310 10124
rect 28276 10121 28304 10152
rect 29641 10149 29653 10183
rect 29687 10180 29699 10183
rect 29932 10180 29960 10208
rect 31297 10183 31355 10189
rect 31297 10180 31309 10183
rect 29687 10152 29960 10180
rect 30866 10152 31309 10180
rect 29687 10149 29699 10152
rect 29641 10143 29699 10149
rect 31297 10149 31309 10152
rect 31343 10149 31355 10183
rect 31297 10143 31355 10149
rect 27525 10115 27583 10121
rect 27525 10081 27537 10115
rect 27571 10081 27583 10115
rect 27525 10075 27583 10081
rect 28261 10115 28319 10121
rect 28261 10081 28273 10115
rect 28307 10081 28319 10115
rect 28261 10075 28319 10081
rect 28721 10115 28779 10121
rect 28721 10081 28733 10115
rect 28767 10112 28779 10115
rect 28767 10084 28856 10112
rect 28767 10081 28779 10084
rect 28721 10075 28779 10081
rect 19300 10016 19840 10044
rect 22281 10047 22339 10053
rect 19300 10004 19306 10016
rect 22281 10013 22293 10047
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 3234 9868 3240 9920
rect 3292 9868 3298 9920
rect 4338 9868 4344 9920
rect 4396 9868 4402 9920
rect 17954 9868 17960 9920
rect 18012 9868 18018 9920
rect 18506 9868 18512 9920
rect 18564 9868 18570 9920
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 20714 9908 20720 9920
rect 19935 9880 20720 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 21450 9868 21456 9920
rect 21508 9908 21514 9920
rect 22296 9908 22324 10007
rect 22370 10004 22376 10056
rect 22428 10044 22434 10056
rect 22465 10047 22523 10053
rect 22465 10044 22477 10047
rect 22428 10016 22477 10044
rect 22428 10004 22434 10016
rect 22465 10013 22477 10016
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10044 22707 10047
rect 23566 10044 23572 10056
rect 22695 10016 23572 10044
rect 22695 10013 22707 10016
rect 22649 10007 22707 10013
rect 23566 10004 23572 10016
rect 23624 10004 23630 10056
rect 24029 10047 24087 10053
rect 24029 10013 24041 10047
rect 24075 10013 24087 10047
rect 24029 10007 24087 10013
rect 26789 10047 26847 10053
rect 26789 10013 26801 10047
rect 26835 10013 26847 10047
rect 26896 10044 26924 10072
rect 27540 10044 27568 10075
rect 26896 10016 27568 10044
rect 26789 10007 26847 10013
rect 23109 9979 23167 9985
rect 23109 9945 23121 9979
rect 23155 9976 23167 9979
rect 24044 9976 24072 10007
rect 23155 9948 24072 9976
rect 26804 9976 26832 10007
rect 27706 10004 27712 10056
rect 27764 10004 27770 10056
rect 27982 10004 27988 10056
rect 28040 10044 28046 10056
rect 28077 10047 28135 10053
rect 28077 10044 28089 10047
rect 28040 10016 28089 10044
rect 28040 10004 28046 10016
rect 28077 10013 28089 10016
rect 28123 10013 28135 10047
rect 28077 10007 28135 10013
rect 27724 9976 27752 10004
rect 26804 9948 27752 9976
rect 23155 9945 23167 9948
rect 23109 9939 23167 9945
rect 21508 9880 22324 9908
rect 21508 9868 21514 9880
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 24397 9911 24455 9917
rect 24397 9908 24409 9911
rect 23532 9880 24409 9908
rect 23532 9868 23538 9880
rect 24397 9877 24409 9880
rect 24443 9877 24455 9911
rect 24397 9871 24455 9877
rect 27341 9911 27399 9917
rect 27341 9877 27353 9911
rect 27387 9908 27399 9911
rect 27430 9908 27436 9920
rect 27387 9880 27436 9908
rect 27387 9877 27399 9880
rect 27341 9871 27399 9877
rect 27430 9868 27436 9880
rect 27488 9908 27494 9920
rect 27890 9908 27896 9920
rect 27488 9880 27896 9908
rect 27488 9868 27494 9880
rect 27890 9868 27896 9880
rect 27948 9868 27954 9920
rect 28258 9868 28264 9920
rect 28316 9868 28322 9920
rect 28445 9911 28503 9917
rect 28445 9877 28457 9911
rect 28491 9908 28503 9911
rect 28718 9908 28724 9920
rect 28491 9880 28724 9908
rect 28491 9877 28503 9880
rect 28445 9871 28503 9877
rect 28718 9868 28724 9880
rect 28776 9868 28782 9920
rect 28828 9908 28856 10084
rect 28902 10072 28908 10124
rect 28960 10072 28966 10124
rect 28997 10115 29055 10121
rect 28997 10081 29009 10115
rect 29043 10081 29055 10115
rect 28997 10075 29055 10081
rect 29012 10044 29040 10075
rect 29086 10072 29092 10124
rect 29144 10072 29150 10124
rect 31386 10072 31392 10124
rect 31444 10072 31450 10124
rect 31478 10072 31484 10124
rect 31536 10072 31542 10124
rect 31665 10115 31723 10121
rect 31665 10081 31677 10115
rect 31711 10081 31723 10115
rect 31665 10075 31723 10081
rect 29012 10016 29132 10044
rect 29104 9976 29132 10016
rect 29362 10004 29368 10056
rect 29420 10004 29426 10056
rect 29638 10044 29644 10056
rect 29472 10016 29644 10044
rect 29472 9976 29500 10016
rect 29638 10004 29644 10016
rect 29696 10004 29702 10056
rect 30190 10004 30196 10056
rect 30248 10044 30254 10056
rect 31680 10044 31708 10075
rect 30248 10016 31708 10044
rect 30248 10004 30254 10016
rect 29104 9948 29500 9976
rect 31481 9911 31539 9917
rect 31481 9908 31493 9911
rect 28828 9880 31493 9908
rect 31481 9877 31493 9880
rect 31527 9877 31539 9911
rect 31481 9871 31539 9877
rect 2760 9818 32200 9840
rect 2760 9766 6286 9818
rect 6338 9766 6350 9818
rect 6402 9766 6414 9818
rect 6466 9766 6478 9818
rect 6530 9766 6542 9818
rect 6594 9766 13646 9818
rect 13698 9766 13710 9818
rect 13762 9766 13774 9818
rect 13826 9766 13838 9818
rect 13890 9766 13902 9818
rect 13954 9766 21006 9818
rect 21058 9766 21070 9818
rect 21122 9766 21134 9818
rect 21186 9766 21198 9818
rect 21250 9766 21262 9818
rect 21314 9766 28366 9818
rect 28418 9766 28430 9818
rect 28482 9766 28494 9818
rect 28546 9766 28558 9818
rect 28610 9766 28622 9818
rect 28674 9766 32200 9818
rect 2760 9744 32200 9766
rect 14553 9707 14611 9713
rect 14553 9673 14565 9707
rect 14599 9673 14611 9707
rect 14553 9667 14611 9673
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 8757 9571 8815 9577
rect 8757 9568 8769 9571
rect 8720 9540 8769 9568
rect 8720 9528 8726 9540
rect 8757 9537 8769 9540
rect 8803 9537 8815 9571
rect 14568 9568 14596 9667
rect 14918 9664 14924 9716
rect 14976 9664 14982 9716
rect 15194 9664 15200 9716
rect 15252 9664 15258 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15436 9676 15945 9704
rect 15436 9664 15442 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 15933 9667 15991 9673
rect 21637 9707 21695 9713
rect 21637 9673 21649 9707
rect 21683 9704 21695 9707
rect 21818 9704 21824 9716
rect 21683 9676 21824 9704
rect 21683 9673 21695 9676
rect 21637 9667 21695 9673
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 22554 9704 22560 9716
rect 21928 9676 22560 9704
rect 14737 9639 14795 9645
rect 14737 9605 14749 9639
rect 14783 9636 14795 9639
rect 15212 9636 15240 9664
rect 21928 9648 21956 9676
rect 22554 9664 22560 9676
rect 22612 9704 22618 9716
rect 23198 9704 23204 9716
rect 22612 9676 23204 9704
rect 22612 9664 22618 9676
rect 23198 9664 23204 9676
rect 23256 9664 23262 9716
rect 24118 9704 24124 9716
rect 23492 9676 24124 9704
rect 14783 9608 15240 9636
rect 14783 9605 14795 9608
rect 14737 9599 14795 9605
rect 15838 9596 15844 9648
rect 15896 9636 15902 9648
rect 19150 9636 19156 9648
rect 15896 9608 19156 9636
rect 15896 9596 15902 9608
rect 19150 9596 19156 9608
rect 19208 9596 19214 9648
rect 21085 9639 21143 9645
rect 21085 9636 21097 9639
rect 20364 9608 21097 9636
rect 15010 9568 15016 9580
rect 14568 9540 15016 9568
rect 8757 9531 8815 9537
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 15473 9571 15531 9577
rect 15473 9568 15485 9571
rect 15344 9540 15485 9568
rect 15344 9528 15350 9540
rect 15473 9537 15485 9540
rect 15519 9537 15531 9571
rect 15473 9531 15531 9537
rect 16574 9528 16580 9580
rect 16632 9528 16638 9580
rect 20254 9528 20260 9580
rect 20312 9528 20318 9580
rect 20364 9512 20392 9608
rect 21085 9605 21097 9608
rect 21131 9636 21143 9639
rect 21910 9636 21916 9648
rect 21131 9608 21916 9636
rect 21131 9605 21143 9608
rect 21085 9599 21143 9605
rect 20717 9571 20775 9577
rect 20717 9537 20729 9571
rect 20763 9568 20775 9571
rect 20898 9568 20904 9580
rect 20763 9540 20904 9568
rect 20763 9537 20775 9540
rect 20717 9531 20775 9537
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 13998 9460 14004 9512
rect 14056 9500 14062 9512
rect 14185 9503 14243 9509
rect 14185 9500 14197 9503
rect 14056 9472 14197 9500
rect 14056 9460 14062 9472
rect 14185 9469 14197 9472
rect 14231 9500 14243 9503
rect 14231 9472 15976 9500
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 15948 9376 15976 9472
rect 16666 9460 16672 9512
rect 16724 9460 16730 9512
rect 18046 9460 18052 9512
rect 18104 9460 18110 9512
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 20027 9472 20085 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 20346 9460 20352 9512
rect 20404 9460 20410 9512
rect 20806 9460 20812 9512
rect 20864 9460 20870 9512
rect 18598 9392 18604 9444
rect 18656 9432 18662 9444
rect 18656 9404 20208 9432
rect 18656 9392 18662 9404
rect 20180 9376 20208 9404
rect 8205 9367 8263 9373
rect 8205 9333 8217 9367
rect 8251 9364 8263 9367
rect 8294 9364 8300 9376
rect 8251 9336 8300 9364
rect 8251 9333 8263 9336
rect 8205 9327 8263 9333
rect 8294 9324 8300 9336
rect 8352 9364 8358 9376
rect 9582 9364 9588 9376
rect 8352 9336 9588 9364
rect 8352 9324 8358 9336
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 13538 9324 13544 9376
rect 13596 9364 13602 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13596 9336 14013 9364
rect 13596 9324 13602 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 14001 9327 14059 9333
rect 14090 9324 14096 9376
rect 14148 9364 14154 9376
rect 14553 9367 14611 9373
rect 14553 9364 14565 9367
rect 14148 9336 14565 9364
rect 14148 9324 14154 9336
rect 14553 9333 14565 9336
rect 14599 9333 14611 9367
rect 14553 9327 14611 9333
rect 15930 9324 15936 9376
rect 15988 9324 15994 9376
rect 17313 9367 17371 9373
rect 17313 9333 17325 9367
rect 17359 9364 17371 9367
rect 17678 9364 17684 9376
rect 17359 9336 17684 9364
rect 17359 9333 17371 9336
rect 17313 9327 17371 9333
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 18966 9324 18972 9376
rect 19024 9324 19030 9376
rect 19337 9367 19395 9373
rect 19337 9333 19349 9367
rect 19383 9364 19395 9367
rect 19610 9364 19616 9376
rect 19383 9336 19616 9364
rect 19383 9333 19395 9336
rect 19337 9327 19395 9333
rect 19610 9324 19616 9336
rect 19668 9324 19674 9376
rect 20162 9324 20168 9376
rect 20220 9324 20226 9376
rect 20824 9364 20852 9460
rect 21100 9432 21128 9599
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 22005 9639 22063 9645
rect 22005 9605 22017 9639
rect 22051 9636 22063 9639
rect 22462 9636 22468 9648
rect 22051 9608 22468 9636
rect 22051 9605 22063 9608
rect 22005 9599 22063 9605
rect 22462 9596 22468 9608
rect 22520 9596 22526 9648
rect 22649 9639 22707 9645
rect 22649 9605 22661 9639
rect 22695 9636 22707 9639
rect 22738 9636 22744 9648
rect 22695 9608 22744 9636
rect 22695 9605 22707 9608
rect 22649 9599 22707 9605
rect 22738 9596 22744 9608
rect 22796 9596 22802 9648
rect 23492 9636 23520 9676
rect 24118 9664 24124 9676
rect 24176 9664 24182 9716
rect 24302 9664 24308 9716
rect 24360 9704 24366 9716
rect 25133 9707 25191 9713
rect 25133 9704 25145 9707
rect 24360 9676 25145 9704
rect 24360 9664 24366 9676
rect 25133 9673 25145 9676
rect 25179 9673 25191 9707
rect 25133 9667 25191 9673
rect 26602 9664 26608 9716
rect 26660 9704 26666 9716
rect 27246 9704 27252 9716
rect 26660 9676 27252 9704
rect 26660 9664 26666 9676
rect 27246 9664 27252 9676
rect 27304 9664 27310 9716
rect 27525 9707 27583 9713
rect 27525 9704 27537 9707
rect 27356 9676 27537 9704
rect 22848 9608 23520 9636
rect 22848 9568 22876 9608
rect 23566 9596 23572 9648
rect 23624 9636 23630 9648
rect 25225 9639 25283 9645
rect 25225 9636 25237 9639
rect 23624 9608 25237 9636
rect 23624 9596 23630 9608
rect 25225 9605 25237 9608
rect 25271 9605 25283 9639
rect 25225 9599 25283 9605
rect 25406 9596 25412 9648
rect 25464 9636 25470 9648
rect 27356 9636 27384 9676
rect 27525 9673 27537 9676
rect 27571 9673 27583 9707
rect 27525 9667 27583 9673
rect 27798 9664 27804 9716
rect 27856 9664 27862 9716
rect 27890 9664 27896 9716
rect 27948 9704 27954 9716
rect 28169 9707 28227 9713
rect 28169 9704 28181 9707
rect 27948 9676 28181 9704
rect 27948 9664 27954 9676
rect 28169 9673 28181 9676
rect 28215 9673 28227 9707
rect 29454 9704 29460 9716
rect 28169 9667 28227 9673
rect 28644 9676 29460 9704
rect 25464 9608 27384 9636
rect 25464 9596 25470 9608
rect 27430 9596 27436 9648
rect 27488 9596 27494 9648
rect 27816 9636 27844 9664
rect 28353 9639 28411 9645
rect 27540 9608 27844 9636
rect 27908 9608 28212 9636
rect 25317 9571 25375 9577
rect 25317 9568 25329 9571
rect 21284 9540 22140 9568
rect 21284 9512 21312 9540
rect 22112 9512 22140 9540
rect 22204 9540 22876 9568
rect 23492 9540 25084 9568
rect 21266 9460 21272 9512
rect 21324 9460 21330 9512
rect 21910 9460 21916 9512
rect 21968 9460 21974 9512
rect 22094 9460 22100 9512
rect 22152 9460 22158 9512
rect 22204 9509 22232 9540
rect 23492 9512 23520 9540
rect 22189 9503 22247 9509
rect 22189 9469 22201 9503
rect 22235 9469 22247 9503
rect 22189 9463 22247 9469
rect 22278 9460 22284 9512
rect 22336 9500 22342 9512
rect 22373 9503 22431 9509
rect 22373 9500 22385 9503
rect 22336 9472 22385 9500
rect 22336 9460 22342 9472
rect 22373 9469 22385 9472
rect 22419 9469 22431 9503
rect 23474 9500 23480 9512
rect 22373 9463 22431 9469
rect 22848 9472 23480 9500
rect 21453 9435 21511 9441
rect 21453 9432 21465 9435
rect 21100 9404 21465 9432
rect 21453 9401 21465 9404
rect 21499 9401 21511 9435
rect 22848 9432 22876 9472
rect 23474 9460 23480 9472
rect 23532 9460 23538 9512
rect 23658 9460 23664 9512
rect 23716 9460 23722 9512
rect 23753 9503 23811 9509
rect 23753 9469 23765 9503
rect 23799 9500 23811 9503
rect 23842 9500 23848 9512
rect 23799 9472 23848 9500
rect 23799 9469 23811 9472
rect 23753 9463 23811 9469
rect 23842 9460 23848 9472
rect 23900 9460 23906 9512
rect 24762 9500 24768 9512
rect 24044 9472 24768 9500
rect 21453 9395 21511 9401
rect 22112 9404 22876 9432
rect 21174 9364 21180 9376
rect 20824 9336 21180 9364
rect 21174 9324 21180 9336
rect 21232 9364 21238 9376
rect 21653 9367 21711 9373
rect 21653 9364 21665 9367
rect 21232 9336 21665 9364
rect 21232 9324 21238 9336
rect 21653 9333 21665 9336
rect 21699 9333 21711 9367
rect 21653 9327 21711 9333
rect 21821 9367 21879 9373
rect 21821 9333 21833 9367
rect 21867 9364 21879 9367
rect 22112 9364 22140 9404
rect 22922 9392 22928 9444
rect 22980 9392 22986 9444
rect 23382 9432 23388 9444
rect 23032 9404 23388 9432
rect 21867 9336 22140 9364
rect 22281 9367 22339 9373
rect 21867 9333 21879 9336
rect 21821 9327 21879 9333
rect 22281 9333 22293 9367
rect 22327 9364 22339 9367
rect 23032 9364 23060 9404
rect 23382 9392 23388 9404
rect 23440 9392 23446 9444
rect 22327 9336 23060 9364
rect 23676 9364 23704 9460
rect 23934 9392 23940 9444
rect 23992 9392 23998 9444
rect 24044 9373 24072 9472
rect 24762 9460 24768 9472
rect 24820 9460 24826 9512
rect 25056 9509 25084 9540
rect 25148 9540 25329 9568
rect 25041 9503 25099 9509
rect 25041 9469 25053 9503
rect 25087 9469 25099 9503
rect 25041 9463 25099 9469
rect 25148 9444 25176 9540
rect 25317 9537 25329 9540
rect 25363 9537 25375 9571
rect 27448 9568 27476 9596
rect 25317 9531 25375 9537
rect 26804 9540 27476 9568
rect 25222 9460 25228 9512
rect 25280 9500 25286 9512
rect 25409 9503 25467 9509
rect 25409 9500 25421 9503
rect 25280 9472 25421 9500
rect 25280 9460 25286 9472
rect 25409 9469 25421 9472
rect 25455 9469 25467 9503
rect 25409 9463 25467 9469
rect 25593 9503 25651 9509
rect 25593 9469 25605 9503
rect 25639 9469 25651 9503
rect 25593 9463 25651 9469
rect 24578 9392 24584 9444
rect 24636 9392 24642 9444
rect 25130 9392 25136 9444
rect 25188 9392 25194 9444
rect 25608 9432 25636 9463
rect 25682 9460 25688 9512
rect 25740 9460 25746 9512
rect 25869 9503 25927 9509
rect 25869 9469 25881 9503
rect 25915 9500 25927 9503
rect 25915 9472 26556 9500
rect 25915 9469 25927 9472
rect 25869 9463 25927 9469
rect 25332 9404 25636 9432
rect 25777 9435 25835 9441
rect 24029 9367 24087 9373
rect 24029 9364 24041 9367
rect 23676 9336 24041 9364
rect 22327 9333 22339 9336
rect 22281 9327 22339 9333
rect 24029 9333 24041 9336
rect 24075 9333 24087 9367
rect 24029 9327 24087 9333
rect 24394 9324 24400 9376
rect 24452 9324 24458 9376
rect 24949 9367 25007 9373
rect 24949 9333 24961 9367
rect 24995 9364 25007 9367
rect 25332 9364 25360 9404
rect 25777 9401 25789 9435
rect 25823 9432 25835 9435
rect 25823 9404 26188 9432
rect 25823 9401 25835 9404
rect 25777 9395 25835 9401
rect 24995 9336 25360 9364
rect 24995 9333 25007 9336
rect 24949 9327 25007 9333
rect 25406 9324 25412 9376
rect 25464 9324 25470 9376
rect 25866 9324 25872 9376
rect 25924 9364 25930 9376
rect 26053 9367 26111 9373
rect 26053 9364 26065 9367
rect 25924 9336 26065 9364
rect 25924 9324 25930 9336
rect 26053 9333 26065 9336
rect 26099 9333 26111 9367
rect 26160 9364 26188 9404
rect 26234 9392 26240 9444
rect 26292 9392 26298 9444
rect 26326 9392 26332 9444
rect 26384 9432 26390 9444
rect 26421 9435 26479 9441
rect 26421 9432 26433 9435
rect 26384 9404 26433 9432
rect 26384 9392 26390 9404
rect 26421 9401 26433 9404
rect 26467 9401 26479 9435
rect 26528 9432 26556 9472
rect 26602 9460 26608 9512
rect 26660 9460 26666 9512
rect 26804 9509 26832 9540
rect 27540 9509 27568 9608
rect 27706 9528 27712 9580
rect 27764 9528 27770 9580
rect 27908 9577 27936 9608
rect 28184 9580 28212 9608
rect 28353 9605 28365 9639
rect 28399 9636 28411 9639
rect 28644 9636 28672 9676
rect 29454 9664 29460 9676
rect 29512 9664 29518 9716
rect 29638 9664 29644 9716
rect 29696 9704 29702 9716
rect 29733 9707 29791 9713
rect 29733 9704 29745 9707
rect 29696 9676 29745 9704
rect 29696 9664 29702 9676
rect 29733 9673 29745 9676
rect 29779 9673 29791 9707
rect 29733 9667 29791 9673
rect 28399 9608 28672 9636
rect 28399 9605 28411 9608
rect 28353 9599 28411 9605
rect 28994 9596 29000 9648
rect 29052 9636 29058 9648
rect 29549 9639 29607 9645
rect 29549 9636 29561 9639
rect 29052 9608 29561 9636
rect 29052 9596 29058 9608
rect 29549 9605 29561 9608
rect 29595 9605 29607 9639
rect 29549 9599 29607 9605
rect 27893 9571 27951 9577
rect 27893 9537 27905 9571
rect 27939 9537 27951 9571
rect 27893 9531 27951 9537
rect 28166 9528 28172 9580
rect 28224 9568 28230 9580
rect 28224 9540 28396 9568
rect 28224 9528 28230 9540
rect 26789 9503 26847 9509
rect 26789 9469 26801 9503
rect 26835 9469 26847 9503
rect 27279 9503 27337 9509
rect 27279 9500 27291 9503
rect 26789 9463 26847 9469
rect 26988 9472 27291 9500
rect 26988 9444 27016 9472
rect 27279 9469 27291 9472
rect 27325 9469 27337 9503
rect 27279 9463 27337 9469
rect 27433 9503 27491 9509
rect 27433 9469 27445 9503
rect 27479 9469 27491 9503
rect 27433 9463 27491 9469
rect 27525 9503 27583 9509
rect 27525 9469 27537 9503
rect 27571 9469 27583 9503
rect 27525 9463 27583 9469
rect 27801 9503 27859 9509
rect 27801 9469 27813 9503
rect 27847 9500 27859 9503
rect 28258 9500 28264 9512
rect 27847 9472 28264 9500
rect 27847 9469 27859 9472
rect 27801 9463 27859 9469
rect 26970 9432 26976 9444
rect 26528 9404 26976 9432
rect 26421 9395 26479 9401
rect 26970 9392 26976 9404
rect 27028 9392 27034 9444
rect 26878 9364 26884 9376
rect 26160 9336 26884 9364
rect 26053 9327 26111 9333
rect 26878 9324 26884 9336
rect 26936 9324 26942 9376
rect 27062 9324 27068 9376
rect 27120 9324 27126 9376
rect 27448 9364 27476 9463
rect 28258 9460 28264 9472
rect 28316 9460 28322 9512
rect 27614 9392 27620 9444
rect 27672 9432 27678 9444
rect 27985 9435 28043 9441
rect 27985 9432 27997 9435
rect 27672 9404 27997 9432
rect 27672 9392 27678 9404
rect 27985 9401 27997 9404
rect 28031 9401 28043 9435
rect 28368 9432 28396 9540
rect 28534 9528 28540 9580
rect 28592 9568 28598 9580
rect 29108 9571 29166 9577
rect 29108 9568 29120 9571
rect 28592 9540 29120 9568
rect 28592 9528 28598 9540
rect 29108 9537 29120 9540
rect 29154 9537 29166 9571
rect 30466 9568 30472 9580
rect 29108 9531 29166 9537
rect 29748 9540 30472 9568
rect 28442 9460 28448 9512
rect 28500 9460 28506 9512
rect 28629 9503 28687 9509
rect 28629 9469 28641 9503
rect 28675 9500 28687 9503
rect 28718 9500 28724 9512
rect 28675 9472 28724 9500
rect 28675 9469 28687 9472
rect 28629 9463 28687 9469
rect 28718 9460 28724 9472
rect 28776 9500 28782 9512
rect 28905 9503 28963 9509
rect 28905 9500 28917 9503
rect 28776 9472 28917 9500
rect 28776 9460 28782 9472
rect 28905 9469 28917 9472
rect 28951 9469 28963 9503
rect 28905 9463 28963 9469
rect 28997 9503 29055 9509
rect 28997 9469 29009 9503
rect 29043 9500 29055 9503
rect 29546 9500 29552 9512
rect 29043 9472 29552 9500
rect 29043 9469 29055 9472
rect 28997 9463 29055 9469
rect 29546 9460 29552 9472
rect 29604 9460 29610 9512
rect 29748 9509 29776 9540
rect 30466 9528 30472 9540
rect 30524 9528 30530 9580
rect 29733 9503 29791 9509
rect 29733 9469 29745 9503
rect 29779 9469 29791 9503
rect 29733 9463 29791 9469
rect 30101 9503 30159 9509
rect 30101 9469 30113 9503
rect 30147 9469 30159 9503
rect 30101 9463 30159 9469
rect 30193 9503 30251 9509
rect 30193 9469 30205 9503
rect 30239 9500 30251 9503
rect 30374 9500 30380 9512
rect 30239 9472 30380 9500
rect 30239 9469 30251 9472
rect 30193 9463 30251 9469
rect 29178 9441 29184 9444
rect 28368 9404 29040 9432
rect 27985 9395 28043 9401
rect 29012 9376 29040 9404
rect 29177 9395 29184 9441
rect 29178 9392 29184 9395
rect 29236 9392 29242 9444
rect 30116 9432 30144 9463
rect 30374 9460 30380 9472
rect 30432 9460 30438 9512
rect 30650 9460 30656 9512
rect 30708 9500 30714 9512
rect 30929 9503 30987 9509
rect 30929 9500 30941 9503
rect 30708 9472 30941 9500
rect 30708 9460 30714 9472
rect 30929 9469 30941 9472
rect 30975 9469 30987 9503
rect 30929 9463 30987 9469
rect 31202 9460 31208 9512
rect 31260 9460 31266 9512
rect 30282 9432 30288 9444
rect 30116 9404 30288 9432
rect 30282 9392 30288 9404
rect 30340 9392 30346 9444
rect 27522 9364 27528 9376
rect 27448 9336 27528 9364
rect 27522 9324 27528 9336
rect 27580 9324 27586 9376
rect 27798 9324 27804 9376
rect 27856 9364 27862 9376
rect 28185 9367 28243 9373
rect 28185 9364 28197 9367
rect 27856 9336 28197 9364
rect 27856 9324 27862 9336
rect 28185 9333 28197 9336
rect 28231 9333 28243 9367
rect 28185 9327 28243 9333
rect 28350 9324 28356 9376
rect 28408 9364 28414 9376
rect 28813 9367 28871 9373
rect 28813 9364 28825 9367
rect 28408 9336 28825 9364
rect 28408 9324 28414 9336
rect 28813 9333 28825 9336
rect 28859 9364 28871 9367
rect 28902 9364 28908 9376
rect 28859 9336 28908 9364
rect 28859 9333 28871 9336
rect 28813 9327 28871 9333
rect 28902 9324 28908 9336
rect 28960 9324 28966 9376
rect 28994 9324 29000 9376
rect 29052 9324 29058 9376
rect 30098 9324 30104 9376
rect 30156 9364 30162 9376
rect 30377 9367 30435 9373
rect 30377 9364 30389 9367
rect 30156 9336 30389 9364
rect 30156 9324 30162 9336
rect 30377 9333 30389 9336
rect 30423 9333 30435 9367
rect 30377 9327 30435 9333
rect 31849 9367 31907 9373
rect 31849 9333 31861 9367
rect 31895 9364 31907 9367
rect 31895 9336 32260 9364
rect 31895 9333 31907 9336
rect 31849 9327 31907 9333
rect 2760 9274 32200 9296
rect 2760 9222 6946 9274
rect 6998 9222 7010 9274
rect 7062 9222 7074 9274
rect 7126 9222 7138 9274
rect 7190 9222 7202 9274
rect 7254 9222 14306 9274
rect 14358 9222 14370 9274
rect 14422 9222 14434 9274
rect 14486 9222 14498 9274
rect 14550 9222 14562 9274
rect 14614 9222 21666 9274
rect 21718 9222 21730 9274
rect 21782 9222 21794 9274
rect 21846 9222 21858 9274
rect 21910 9222 21922 9274
rect 21974 9222 29026 9274
rect 29078 9222 29090 9274
rect 29142 9222 29154 9274
rect 29206 9222 29218 9274
rect 29270 9222 29282 9274
rect 29334 9222 32200 9274
rect 2760 9200 32200 9222
rect 6365 9163 6423 9169
rect 6365 9129 6377 9163
rect 6411 9160 6423 9163
rect 6730 9160 6736 9172
rect 6411 9132 6736 9160
rect 6411 9129 6423 9132
rect 6365 9123 6423 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 10505 9163 10563 9169
rect 10505 9160 10517 9163
rect 7524 9132 10517 9160
rect 7524 9120 7530 9132
rect 10505 9129 10517 9132
rect 10551 9129 10563 9163
rect 10505 9123 10563 9129
rect 12529 9163 12587 9169
rect 12529 9129 12541 9163
rect 12575 9160 12587 9163
rect 14090 9160 14096 9172
rect 12575 9132 14096 9160
rect 12575 9129 12587 9132
rect 12529 9123 12587 9129
rect 10520 9024 10548 9123
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 15838 9160 15844 9172
rect 14292 9132 15844 9160
rect 13541 9095 13599 9101
rect 13541 9061 13553 9095
rect 13587 9092 13599 9095
rect 14292 9092 14320 9132
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 16393 9163 16451 9169
rect 16393 9129 16405 9163
rect 16439 9160 16451 9163
rect 16666 9160 16672 9172
rect 16439 9132 16672 9160
rect 16439 9129 16451 9132
rect 16393 9123 16451 9129
rect 16666 9120 16672 9132
rect 16724 9120 16730 9172
rect 17589 9163 17647 9169
rect 17589 9129 17601 9163
rect 17635 9160 17647 9163
rect 18598 9160 18604 9172
rect 17635 9132 18604 9160
rect 17635 9129 17647 9132
rect 17589 9123 17647 9129
rect 18598 9120 18604 9132
rect 18656 9120 18662 9172
rect 23201 9163 23259 9169
rect 19444 9132 21496 9160
rect 13587 9064 14320 9092
rect 13587 9061 13599 9064
rect 13541 9055 13599 9061
rect 14366 9052 14372 9104
rect 14424 9052 14430 9104
rect 17954 9092 17960 9104
rect 17880 9064 17960 9092
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10520 8996 10701 9024
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 10870 8984 10876 9036
rect 10928 8984 10934 9036
rect 13998 8984 14004 9036
rect 14056 8984 14062 9036
rect 16666 9024 16672 9036
rect 16054 8996 16672 9024
rect 16666 8984 16672 8996
rect 16724 8984 16730 9036
rect 11606 8916 11612 8968
rect 11664 8916 11670 8968
rect 11698 8916 11704 8968
rect 11756 8965 11762 8968
rect 11756 8959 11784 8965
rect 11772 8925 11784 8959
rect 11756 8919 11784 8925
rect 11885 8959 11943 8965
rect 11885 8925 11897 8959
rect 11931 8956 11943 8959
rect 13538 8956 13544 8968
rect 11931 8928 13544 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 11756 8916 11762 8919
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 14090 8916 14096 8968
rect 14148 8956 14154 8968
rect 14642 8956 14648 8968
rect 14148 8928 14648 8956
rect 14148 8916 14154 8928
rect 14642 8916 14648 8928
rect 14700 8916 14706 8968
rect 14918 8916 14924 8968
rect 14976 8916 14982 8968
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16356 8928 17049 8956
rect 16356 8916 16362 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 17880 8965 17908 9064
rect 17954 9052 17960 9064
rect 18012 9092 18018 9104
rect 18966 9092 18972 9104
rect 18012 9064 18972 9092
rect 18012 9052 18018 9064
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 18506 8984 18512 9036
rect 18564 8984 18570 9036
rect 19444 9033 19472 9132
rect 19610 9052 19616 9104
rect 19668 9092 19674 9104
rect 19705 9095 19763 9101
rect 19705 9092 19717 9095
rect 19668 9064 19717 9092
rect 19668 9052 19674 9064
rect 19705 9061 19717 9064
rect 19751 9061 19763 9095
rect 19705 9055 19763 9061
rect 20714 9052 20720 9104
rect 20772 9052 20778 9104
rect 21266 9052 21272 9104
rect 21324 9052 21330 9104
rect 19429 9027 19487 9033
rect 19429 9024 19441 9027
rect 18800 8996 19441 9024
rect 18800 8968 18828 8996
rect 19429 8993 19441 8996
rect 19475 8993 19487 9027
rect 19429 8987 19487 8993
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 18782 8916 18788 8968
rect 18840 8916 18846 8968
rect 19242 8916 19248 8968
rect 19300 8916 19306 8968
rect 21177 8959 21235 8965
rect 21177 8925 21189 8959
rect 21223 8956 21235 8959
rect 21284 8956 21312 9052
rect 21468 9036 21496 9132
rect 23201 9129 23213 9163
rect 23247 9160 23259 9163
rect 23934 9160 23940 9172
rect 23247 9132 23940 9160
rect 23247 9129 23259 9132
rect 23201 9123 23259 9129
rect 23934 9120 23940 9132
rect 23992 9120 23998 9172
rect 25041 9163 25099 9169
rect 25041 9160 25053 9163
rect 24044 9132 25053 9160
rect 24044 9092 24072 9132
rect 25041 9129 25053 9132
rect 25087 9129 25099 9163
rect 25041 9123 25099 9129
rect 25406 9120 25412 9172
rect 25464 9120 25470 9172
rect 26602 9160 26608 9172
rect 25884 9132 26608 9160
rect 22954 9064 24072 9092
rect 24394 9052 24400 9104
rect 24452 9052 24458 9104
rect 25424 9092 25452 9120
rect 24504 9064 25452 9092
rect 21450 8984 21456 9036
rect 21508 8984 21514 9036
rect 23842 8984 23848 9036
rect 23900 9024 23906 9036
rect 24412 9024 24440 9052
rect 24504 9033 24532 9064
rect 23900 8996 24440 9024
rect 24489 9027 24547 9033
rect 23900 8984 23906 8996
rect 24489 8993 24501 9027
rect 24535 8993 24547 9027
rect 24489 8987 24547 8993
rect 24762 8984 24768 9036
rect 24820 8984 24826 9036
rect 24946 8984 24952 9036
rect 25004 9024 25010 9036
rect 25133 9027 25191 9033
rect 25133 9024 25145 9027
rect 25004 8996 25145 9024
rect 25004 8984 25010 8996
rect 25133 8993 25145 8996
rect 25179 8993 25191 9027
rect 25133 8987 25191 8993
rect 25682 8984 25688 9036
rect 25740 8984 25746 9036
rect 25777 9027 25835 9033
rect 25777 8993 25789 9027
rect 25823 9024 25835 9027
rect 25884 9024 25912 9132
rect 26602 9120 26608 9132
rect 26660 9120 26666 9172
rect 27062 9120 27068 9172
rect 27120 9120 27126 9172
rect 27246 9120 27252 9172
rect 27304 9160 27310 9172
rect 27341 9163 27399 9169
rect 27341 9160 27353 9163
rect 27304 9132 27353 9160
rect 27304 9120 27310 9132
rect 27341 9129 27353 9132
rect 27387 9129 27399 9163
rect 27341 9123 27399 9129
rect 27430 9120 27436 9172
rect 27488 9120 27494 9172
rect 27525 9163 27583 9169
rect 27525 9129 27537 9163
rect 27571 9160 27583 9163
rect 27798 9160 27804 9172
rect 27571 9132 27804 9160
rect 27571 9129 27583 9132
rect 27525 9123 27583 9129
rect 27798 9120 27804 9132
rect 27856 9120 27862 9172
rect 27890 9120 27896 9172
rect 27948 9160 27954 9172
rect 28350 9160 28356 9172
rect 27948 9132 28356 9160
rect 27948 9120 27954 9132
rect 28350 9120 28356 9132
rect 28408 9120 28414 9172
rect 28442 9120 28448 9172
rect 28500 9160 28506 9172
rect 29546 9160 29552 9172
rect 28500 9132 29552 9160
rect 28500 9120 28506 9132
rect 29546 9120 29552 9132
rect 29604 9120 29610 9172
rect 30098 9160 30104 9172
rect 29840 9132 30104 9160
rect 27080 9092 27108 9120
rect 25976 9064 27108 9092
rect 28905 9095 28963 9101
rect 25976 9033 26004 9064
rect 28905 9061 28917 9095
rect 28951 9092 28963 9095
rect 29454 9092 29460 9104
rect 28951 9064 29460 9092
rect 28951 9061 28963 9064
rect 28905 9055 28963 9061
rect 29454 9052 29460 9064
rect 29512 9052 29518 9104
rect 29840 9101 29868 9132
rect 30098 9120 30104 9132
rect 30156 9120 30162 9172
rect 31202 9120 31208 9172
rect 31260 9160 31266 9172
rect 31297 9163 31355 9169
rect 31297 9160 31309 9163
rect 31260 9132 31309 9160
rect 31260 9120 31266 9132
rect 31297 9129 31309 9132
rect 31343 9129 31355 9163
rect 32232 9160 32260 9336
rect 31297 9123 31355 9129
rect 31726 9132 32260 9160
rect 29825 9095 29883 9101
rect 29825 9061 29837 9095
rect 29871 9061 29883 9095
rect 31110 9092 31116 9104
rect 31050 9064 31116 9092
rect 29825 9055 29883 9061
rect 31110 9052 31116 9064
rect 31168 9052 31174 9104
rect 25823 8996 25912 9024
rect 25961 9027 26019 9033
rect 25823 8993 25835 8996
rect 25777 8987 25835 8993
rect 25961 8993 25973 9027
rect 26007 8993 26019 9027
rect 25961 8987 26019 8993
rect 26418 8984 26424 9036
rect 26476 8984 26482 9036
rect 26602 8984 26608 9036
rect 26660 8984 26666 9036
rect 27985 9027 28043 9033
rect 27985 9024 27997 9027
rect 27540 8996 27997 9024
rect 21223 8928 21312 8956
rect 21729 8959 21787 8965
rect 21223 8925 21235 8928
rect 21177 8919 21235 8925
rect 21729 8925 21741 8959
rect 21775 8956 21787 8959
rect 23477 8959 23535 8965
rect 23477 8956 23489 8959
rect 21775 8928 23489 8956
rect 21775 8925 21787 8928
rect 21729 8919 21787 8925
rect 23477 8925 23489 8928
rect 23523 8925 23535 8959
rect 23477 8919 23535 8925
rect 24121 8959 24179 8965
rect 24121 8925 24133 8959
rect 24167 8925 24179 8959
rect 24121 8919 24179 8925
rect 11333 8891 11391 8897
rect 11333 8857 11345 8891
rect 11379 8857 11391 8891
rect 17954 8888 17960 8900
rect 11333 8851 11391 8857
rect 14384 8860 14780 8888
rect 11348 8820 11376 8851
rect 12897 8823 12955 8829
rect 12897 8820 12909 8823
rect 11348 8792 12909 8820
rect 12897 8789 12909 8792
rect 12943 8820 12955 8823
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 12943 8792 13921 8820
rect 12943 8789 12955 8792
rect 12897 8783 12955 8789
rect 13909 8789 13921 8792
rect 13955 8820 13967 8823
rect 13998 8820 14004 8832
rect 13955 8792 14004 8820
rect 13955 8789 13967 8792
rect 13909 8783 13967 8789
rect 13998 8780 14004 8792
rect 14056 8780 14062 8832
rect 14384 8829 14412 8860
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8789 14427 8823
rect 14369 8783 14427 8789
rect 14553 8823 14611 8829
rect 14553 8789 14565 8823
rect 14599 8820 14611 8823
rect 14642 8820 14648 8832
rect 14599 8792 14648 8820
rect 14599 8789 14611 8792
rect 14553 8783 14611 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14752 8820 14780 8860
rect 16132 8860 17960 8888
rect 16132 8832 16160 8860
rect 17954 8848 17960 8860
rect 18012 8888 18018 8900
rect 18874 8888 18880 8900
rect 18012 8860 18880 8888
rect 18012 8848 18018 8860
rect 18874 8848 18880 8860
rect 18932 8848 18938 8900
rect 24136 8888 24164 8919
rect 24302 8916 24308 8968
rect 24360 8956 24366 8968
rect 24397 8959 24455 8965
rect 24397 8956 24409 8959
rect 24360 8928 24409 8956
rect 24360 8916 24366 8928
rect 24397 8925 24409 8928
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 24670 8916 24676 8968
rect 24728 8956 24734 8968
rect 24857 8959 24915 8965
rect 24857 8956 24869 8959
rect 24728 8928 24869 8956
rect 24728 8916 24734 8928
rect 24857 8925 24869 8928
rect 24903 8925 24915 8959
rect 25866 8956 25872 8968
rect 24857 8919 24915 8925
rect 25792 8928 25872 8956
rect 24213 8891 24271 8897
rect 24213 8888 24225 8891
rect 24136 8860 24225 8888
rect 24213 8857 24225 8860
rect 24259 8857 24271 8891
rect 24872 8888 24900 8919
rect 25792 8888 25820 8928
rect 25866 8916 25872 8928
rect 25924 8916 25930 8968
rect 26620 8956 26648 8984
rect 27540 8956 27568 8996
rect 27985 8993 27997 8996
rect 28031 8993 28043 9027
rect 29114 9027 29172 9033
rect 29114 9024 29126 9027
rect 27985 8987 28043 8993
rect 28920 8996 29126 9024
rect 28920 8968 28948 8996
rect 29114 8993 29126 8996
rect 29160 8993 29172 9027
rect 29114 8987 29172 8993
rect 31573 9027 31631 9033
rect 31573 8993 31585 9027
rect 31619 9024 31631 9027
rect 31726 9024 31754 9132
rect 33134 9092 33140 9104
rect 31864 9064 33140 9092
rect 31864 9033 31892 9064
rect 33134 9052 33140 9064
rect 33192 9052 33198 9104
rect 31619 8996 31754 9024
rect 31849 9027 31907 9033
rect 31619 8993 31631 8996
rect 31573 8987 31631 8993
rect 31849 8993 31861 9027
rect 31895 8993 31907 9027
rect 31849 8987 31907 8993
rect 26620 8928 27568 8956
rect 28074 8916 28080 8968
rect 28132 8956 28138 8968
rect 28169 8959 28227 8965
rect 28169 8956 28181 8959
rect 28132 8928 28181 8956
rect 28132 8916 28138 8928
rect 28169 8925 28181 8928
rect 28215 8925 28227 8959
rect 28169 8919 28227 8925
rect 28626 8916 28632 8968
rect 28684 8916 28690 8968
rect 28902 8916 28908 8968
rect 28960 8916 28966 8968
rect 28997 8959 29055 8965
rect 28997 8925 29009 8959
rect 29043 8925 29055 8959
rect 28997 8919 29055 8925
rect 27062 8888 27068 8900
rect 24872 8860 25820 8888
rect 26068 8860 27068 8888
rect 24213 8851 24271 8857
rect 15010 8820 15016 8832
rect 14752 8792 15016 8820
rect 15010 8780 15016 8792
rect 15068 8820 15074 8832
rect 15378 8820 15384 8832
rect 15068 8792 15384 8820
rect 15068 8780 15074 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 16114 8780 16120 8832
rect 16172 8780 16178 8832
rect 16482 8780 16488 8832
rect 16540 8780 16546 8832
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 17221 8823 17279 8829
rect 17221 8820 17233 8823
rect 17000 8792 17233 8820
rect 17000 8780 17006 8792
rect 17221 8789 17233 8792
rect 17267 8789 17279 8823
rect 17221 8783 17279 8789
rect 18414 8780 18420 8832
rect 18472 8780 18478 8832
rect 18690 8780 18696 8832
rect 18748 8780 18754 8832
rect 21174 8780 21180 8832
rect 21232 8820 21238 8832
rect 21726 8820 21732 8832
rect 21232 8792 21732 8820
rect 21232 8780 21238 8792
rect 21726 8780 21732 8792
rect 21784 8780 21790 8832
rect 21910 8780 21916 8832
rect 21968 8820 21974 8832
rect 23750 8820 23756 8832
rect 21968 8792 23756 8820
rect 21968 8780 21974 8792
rect 23750 8780 23756 8792
rect 23808 8820 23814 8832
rect 25222 8820 25228 8832
rect 23808 8792 25228 8820
rect 23808 8780 23814 8792
rect 25222 8780 25228 8792
rect 25280 8780 25286 8832
rect 25774 8780 25780 8832
rect 25832 8820 25838 8832
rect 26068 8820 26096 8860
rect 27062 8848 27068 8860
rect 27120 8888 27126 8900
rect 27157 8891 27215 8897
rect 27157 8888 27169 8891
rect 27120 8860 27169 8888
rect 27120 8848 27126 8860
rect 27157 8857 27169 8860
rect 27203 8888 27215 8891
rect 28442 8888 28448 8900
rect 27203 8860 28448 8888
rect 27203 8857 27215 8860
rect 27157 8851 27215 8857
rect 28442 8848 28448 8860
rect 28500 8848 28506 8900
rect 29012 8888 29040 8919
rect 29362 8916 29368 8968
rect 29420 8956 29426 8968
rect 29549 8959 29607 8965
rect 29549 8956 29561 8959
rect 29420 8928 29561 8956
rect 29420 8916 29426 8928
rect 29549 8925 29561 8928
rect 29595 8925 29607 8959
rect 31588 8956 31616 8987
rect 29549 8919 29607 8925
rect 29656 8928 31616 8956
rect 29454 8888 29460 8900
rect 29012 8860 29460 8888
rect 29454 8848 29460 8860
rect 29512 8848 29518 8900
rect 29656 8832 29684 8928
rect 31662 8848 31668 8900
rect 31720 8848 31726 8900
rect 25832 8792 26096 8820
rect 25832 8780 25838 8792
rect 26142 8780 26148 8832
rect 26200 8780 26206 8832
rect 26326 8780 26332 8832
rect 26384 8820 26390 8832
rect 27522 8820 27528 8832
rect 26384 8792 27528 8820
rect 26384 8780 26390 8792
rect 27522 8780 27528 8792
rect 27580 8780 27586 8832
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 27709 8823 27767 8829
rect 27709 8820 27721 8823
rect 27672 8792 27721 8820
rect 27672 8780 27678 8792
rect 27709 8789 27721 8792
rect 27755 8789 27767 8823
rect 27709 8783 27767 8789
rect 29270 8780 29276 8832
rect 29328 8780 29334 8832
rect 29638 8780 29644 8832
rect 29696 8780 29702 8832
rect 30282 8780 30288 8832
rect 30340 8820 30346 8832
rect 31478 8820 31484 8832
rect 30340 8792 31484 8820
rect 30340 8780 30346 8792
rect 31478 8780 31484 8792
rect 31536 8780 31542 8832
rect 2760 8730 32200 8752
rect 2760 8678 6286 8730
rect 6338 8678 6350 8730
rect 6402 8678 6414 8730
rect 6466 8678 6478 8730
rect 6530 8678 6542 8730
rect 6594 8678 13646 8730
rect 13698 8678 13710 8730
rect 13762 8678 13774 8730
rect 13826 8678 13838 8730
rect 13890 8678 13902 8730
rect 13954 8678 21006 8730
rect 21058 8678 21070 8730
rect 21122 8678 21134 8730
rect 21186 8678 21198 8730
rect 21250 8678 21262 8730
rect 21314 8678 28366 8730
rect 28418 8678 28430 8730
rect 28482 8678 28494 8730
rect 28546 8678 28558 8730
rect 28610 8678 28622 8730
rect 28674 8678 32200 8730
rect 2760 8656 32200 8678
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 12897 8619 12955 8625
rect 3384 8588 12434 8616
rect 3384 8576 3390 8588
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8548 6239 8551
rect 6227 8520 6868 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8480 5687 8483
rect 6730 8480 6736 8492
rect 5675 8452 6736 8480
rect 5675 8449 5687 8452
rect 5629 8443 5687 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 6840 8489 6868 8520
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 12406 8480 12434 8588
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 14366 8616 14372 8628
rect 12943 8588 14372 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 14366 8576 14372 8588
rect 14424 8576 14430 8628
rect 14734 8576 14740 8628
rect 14792 8576 14798 8628
rect 14918 8576 14924 8628
rect 14976 8576 14982 8628
rect 15838 8576 15844 8628
rect 15896 8576 15902 8628
rect 16482 8576 16488 8628
rect 16540 8576 16546 8628
rect 16942 8576 16948 8628
rect 17000 8576 17006 8628
rect 17037 8619 17095 8625
rect 17037 8585 17049 8619
rect 17083 8616 17095 8619
rect 18322 8616 18328 8628
rect 17083 8588 18328 8616
rect 17083 8585 17095 8588
rect 17037 8579 17095 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 18690 8576 18696 8628
rect 18748 8576 18754 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 19242 8616 19248 8628
rect 18923 8588 19248 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 19242 8576 19248 8588
rect 19300 8576 19306 8628
rect 21358 8576 21364 8628
rect 21416 8576 21422 8628
rect 21821 8619 21879 8625
rect 21821 8585 21833 8619
rect 21867 8616 21879 8619
rect 21910 8616 21916 8628
rect 21867 8588 21916 8616
rect 21867 8585 21879 8588
rect 21821 8579 21879 8585
rect 21910 8576 21916 8588
rect 21968 8576 21974 8628
rect 22002 8576 22008 8628
rect 22060 8576 22066 8628
rect 25130 8616 25136 8628
rect 22664 8588 25136 8616
rect 13998 8508 14004 8560
rect 14056 8548 14062 8560
rect 14093 8551 14151 8557
rect 14093 8548 14105 8551
rect 14056 8520 14105 8548
rect 14056 8508 14062 8520
rect 14093 8517 14105 8520
rect 14139 8548 14151 8551
rect 14752 8548 14780 8576
rect 14139 8520 14780 8548
rect 14139 8517 14151 8520
rect 14093 8511 14151 8517
rect 13679 8483 13737 8489
rect 13679 8480 13691 8483
rect 12406 8452 13691 8480
rect 6825 8443 6883 8449
rect 13679 8449 13691 8452
rect 13725 8449 13737 8483
rect 13679 8443 13737 8449
rect 14737 8483 14795 8489
rect 14737 8449 14749 8483
rect 14783 8480 14795 8483
rect 15856 8480 15884 8576
rect 16500 8548 16528 8576
rect 14783 8452 15884 8480
rect 15948 8520 16528 8548
rect 14783 8449 14795 8452
rect 14737 8443 14795 8449
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 8294 8412 8300 8424
rect 5767 8384 8300 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 13538 8372 13544 8424
rect 13596 8372 13602 8424
rect 13814 8372 13820 8424
rect 13872 8372 13878 8424
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8381 14611 8415
rect 14553 8375 14611 8381
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 4264 8316 5825 8344
rect 4264 8288 4292 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 14568 8344 14596 8375
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 15948 8421 15976 8520
rect 16960 8489 16988 8576
rect 16945 8483 17003 8489
rect 16040 8452 16252 8480
rect 16040 8424 16068 8452
rect 15473 8415 15531 8421
rect 15473 8412 15485 8415
rect 14976 8384 15485 8412
rect 14976 8372 14982 8384
rect 15473 8381 15485 8384
rect 15519 8381 15531 8415
rect 15473 8375 15531 8381
rect 15933 8415 15991 8421
rect 15933 8381 15945 8415
rect 15979 8381 15991 8415
rect 15933 8375 15991 8381
rect 16022 8372 16028 8424
rect 16080 8372 16086 8424
rect 16114 8372 16120 8424
rect 16172 8372 16178 8424
rect 16224 8421 16252 8452
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18708 8480 18736 8576
rect 18966 8508 18972 8560
rect 19024 8548 19030 8560
rect 19024 8520 19564 8548
rect 19024 8508 19030 8520
rect 18555 8452 18736 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 18874 8440 18880 8492
rect 18932 8480 18938 8492
rect 19536 8489 19564 8520
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 18932 8452 19349 8480
rect 18932 8440 18938 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 19567 8452 20024 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 16209 8415 16267 8421
rect 16209 8381 16221 8415
rect 16255 8381 16267 8415
rect 16209 8375 16267 8381
rect 18782 8372 18788 8424
rect 18840 8372 18846 8424
rect 16301 8347 16359 8353
rect 14568 8316 16252 8344
rect 5813 8307 5871 8313
rect 4246 8236 4252 8288
rect 4304 8236 4310 8288
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6273 8279 6331 8285
rect 6273 8276 6285 8279
rect 6236 8248 6285 8276
rect 6236 8236 6242 8248
rect 6273 8245 6285 8248
rect 6319 8245 6331 8279
rect 6273 8239 6331 8245
rect 12713 8279 12771 8285
rect 12713 8245 12725 8279
rect 12759 8276 12771 8279
rect 13538 8276 13544 8288
rect 12759 8248 13544 8276
rect 12759 8245 12771 8248
rect 12713 8239 12771 8245
rect 13538 8236 13544 8248
rect 13596 8276 13602 8288
rect 14826 8276 14832 8288
rect 13596 8248 14832 8276
rect 13596 8236 13602 8248
rect 14826 8236 14832 8248
rect 14884 8236 14890 8288
rect 15746 8236 15752 8288
rect 15804 8236 15810 8288
rect 16224 8276 16252 8316
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 16574 8344 16580 8356
rect 16347 8316 16580 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 18230 8344 18236 8356
rect 16684 8316 17264 8344
rect 18078 8316 18236 8344
rect 16684 8276 16712 8316
rect 16224 8248 16712 8276
rect 17236 8276 17264 8316
rect 18230 8304 18236 8316
rect 18288 8304 18294 8356
rect 19702 8344 19708 8356
rect 18340 8316 19708 8344
rect 18340 8276 18368 8316
rect 19702 8304 19708 8316
rect 19760 8304 19766 8356
rect 17236 8248 18368 8276
rect 19242 8236 19248 8288
rect 19300 8236 19306 8288
rect 19996 8285 20024 8452
rect 20346 8372 20352 8424
rect 20404 8412 20410 8424
rect 20993 8415 21051 8421
rect 20993 8412 21005 8415
rect 20404 8384 21005 8412
rect 20404 8372 20410 8384
rect 20993 8381 21005 8384
rect 21039 8381 21051 8415
rect 20993 8375 21051 8381
rect 21151 8415 21209 8421
rect 21151 8381 21163 8415
rect 21197 8412 21209 8415
rect 21376 8412 21404 8576
rect 21637 8551 21695 8557
rect 21637 8517 21649 8551
rect 21683 8548 21695 8551
rect 22020 8548 22048 8576
rect 21683 8520 22048 8548
rect 21683 8517 21695 8520
rect 21637 8511 21695 8517
rect 22186 8480 22192 8492
rect 21468 8452 22192 8480
rect 21468 8421 21496 8452
rect 22186 8440 22192 8452
rect 22244 8440 22250 8492
rect 21197 8384 21404 8412
rect 21453 8415 21511 8421
rect 21197 8381 21209 8384
rect 21151 8375 21209 8381
rect 21453 8381 21465 8415
rect 21499 8381 21511 8415
rect 21453 8375 21511 8381
rect 21726 8372 21732 8424
rect 21784 8372 21790 8424
rect 22664 8421 22692 8588
rect 25130 8576 25136 8588
rect 25188 8576 25194 8628
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 27433 8619 27491 8625
rect 27433 8616 27445 8619
rect 25740 8588 27445 8616
rect 25740 8576 25746 8588
rect 27433 8585 27445 8588
rect 27479 8585 27491 8619
rect 27433 8579 27491 8585
rect 27890 8576 27896 8628
rect 27948 8576 27954 8628
rect 27982 8576 27988 8628
rect 28040 8616 28046 8628
rect 28353 8619 28411 8625
rect 28353 8616 28365 8619
rect 28040 8588 28365 8616
rect 28040 8576 28046 8588
rect 28353 8585 28365 8588
rect 28399 8585 28411 8619
rect 28353 8579 28411 8585
rect 28810 8576 28816 8628
rect 28868 8576 28874 8628
rect 29089 8619 29147 8625
rect 29089 8585 29101 8619
rect 29135 8616 29147 8619
rect 29730 8616 29736 8628
rect 29135 8588 29736 8616
rect 29135 8585 29147 8588
rect 29089 8579 29147 8585
rect 29730 8576 29736 8588
rect 29788 8576 29794 8628
rect 30469 8619 30527 8625
rect 30469 8585 30481 8619
rect 30515 8616 30527 8619
rect 30650 8616 30656 8628
rect 30515 8588 30656 8616
rect 30515 8585 30527 8588
rect 30469 8579 30527 8585
rect 30650 8576 30656 8588
rect 30708 8576 30714 8628
rect 31110 8576 31116 8628
rect 31168 8616 31174 8628
rect 31297 8619 31355 8625
rect 31297 8616 31309 8619
rect 31168 8588 31309 8616
rect 31168 8576 31174 8588
rect 31297 8585 31309 8588
rect 31343 8585 31355 8619
rect 31297 8579 31355 8585
rect 24305 8551 24363 8557
rect 24305 8548 24317 8551
rect 22848 8520 24317 8548
rect 22848 8489 22876 8520
rect 24305 8517 24317 8520
rect 24351 8517 24363 8551
rect 24305 8511 24363 8517
rect 26878 8508 26884 8560
rect 26936 8548 26942 8560
rect 27522 8548 27528 8560
rect 26936 8520 27528 8548
rect 26936 8508 26942 8520
rect 27522 8508 27528 8520
rect 27580 8548 27586 8560
rect 28828 8548 28856 8576
rect 27580 8520 28856 8548
rect 27580 8508 27586 8520
rect 29638 8508 29644 8560
rect 29696 8508 29702 8560
rect 30929 8551 30987 8557
rect 30929 8548 30941 8551
rect 30852 8520 30941 8548
rect 22833 8483 22891 8489
rect 22833 8449 22845 8483
rect 22879 8449 22891 8483
rect 22833 8443 22891 8449
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 24670 8480 24676 8492
rect 23707 8452 24676 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 21913 8415 21971 8421
rect 21913 8381 21925 8415
rect 21959 8381 21971 8415
rect 21913 8375 21971 8381
rect 22649 8415 22707 8421
rect 22649 8381 22661 8415
rect 22695 8381 22707 8415
rect 22649 8375 22707 8381
rect 20898 8304 20904 8356
rect 20956 8344 20962 8356
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 20956 8316 21281 8344
rect 20956 8304 20962 8316
rect 21269 8313 21281 8316
rect 21315 8313 21327 8347
rect 21269 8307 21327 8313
rect 21361 8347 21419 8353
rect 21361 8313 21373 8347
rect 21407 8344 21419 8347
rect 21542 8344 21548 8356
rect 21407 8316 21548 8344
rect 21407 8313 21419 8316
rect 21361 8307 21419 8313
rect 19981 8279 20039 8285
rect 19981 8245 19993 8279
rect 20027 8276 20039 8279
rect 20438 8276 20444 8288
rect 20027 8248 20444 8276
rect 20027 8245 20039 8248
rect 19981 8239 20039 8245
rect 20438 8236 20444 8248
rect 20496 8236 20502 8288
rect 21284 8276 21312 8307
rect 21542 8304 21548 8316
rect 21600 8304 21606 8356
rect 21928 8344 21956 8375
rect 22002 8344 22008 8356
rect 21928 8316 22008 8344
rect 22002 8304 22008 8316
rect 22060 8304 22066 8356
rect 22848 8344 22876 8443
rect 24670 8440 24676 8452
rect 24728 8440 24734 8492
rect 26142 8440 26148 8492
rect 26200 8440 26206 8492
rect 27062 8440 27068 8492
rect 27120 8440 27126 8492
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8480 27307 8483
rect 29917 8483 29975 8489
rect 27295 8452 28120 8480
rect 27295 8449 27307 8452
rect 27249 8443 27307 8449
rect 28092 8424 28120 8452
rect 28276 8452 29408 8480
rect 23290 8372 23296 8424
rect 23348 8372 23354 8424
rect 23385 8415 23443 8421
rect 23385 8381 23397 8415
rect 23431 8412 23443 8415
rect 24302 8412 24308 8424
rect 23431 8384 24308 8412
rect 23431 8381 23443 8384
rect 23385 8375 23443 8381
rect 23400 8344 23428 8375
rect 24302 8372 24308 8384
rect 24360 8372 24366 8424
rect 24489 8415 24547 8421
rect 24489 8381 24501 8415
rect 24535 8412 24547 8415
rect 24578 8412 24584 8424
rect 24535 8384 24584 8412
rect 24535 8381 24547 8384
rect 24489 8375 24547 8381
rect 24578 8372 24584 8384
rect 24636 8412 24642 8424
rect 24636 8384 24808 8412
rect 24636 8372 24642 8384
rect 22112 8316 22876 8344
rect 23032 8316 23428 8344
rect 23753 8347 23811 8353
rect 22112 8276 22140 8316
rect 21284 8248 22140 8276
rect 22186 8236 22192 8288
rect 22244 8276 22250 8288
rect 22281 8279 22339 8285
rect 22281 8276 22293 8279
rect 22244 8248 22293 8276
rect 22244 8236 22250 8248
rect 22281 8245 22293 8248
rect 22327 8245 22339 8279
rect 22281 8239 22339 8245
rect 22741 8279 22799 8285
rect 22741 8245 22753 8279
rect 22787 8276 22799 8279
rect 23032 8276 23060 8316
rect 23753 8313 23765 8347
rect 23799 8344 23811 8347
rect 24673 8347 24731 8353
rect 24673 8344 24685 8347
rect 23799 8316 24685 8344
rect 23799 8313 23811 8316
rect 23753 8307 23811 8313
rect 24673 8313 24685 8316
rect 24719 8313 24731 8347
rect 24673 8307 24731 8313
rect 22787 8248 23060 8276
rect 22787 8245 22799 8248
rect 22741 8239 22799 8245
rect 23106 8236 23112 8288
rect 23164 8236 23170 8288
rect 23382 8236 23388 8288
rect 23440 8276 23446 8288
rect 24780 8276 24808 8384
rect 25314 8372 25320 8424
rect 25372 8372 25378 8424
rect 25866 8372 25872 8424
rect 25924 8372 25930 8424
rect 26970 8372 26976 8424
rect 27028 8372 27034 8424
rect 27157 8415 27215 8421
rect 27157 8381 27169 8415
rect 27203 8381 27215 8415
rect 27157 8375 27215 8381
rect 27433 8415 27491 8421
rect 27433 8381 27445 8415
rect 27479 8412 27491 8415
rect 27522 8412 27528 8424
rect 27479 8384 27528 8412
rect 27479 8381 27491 8384
rect 27433 8375 27491 8381
rect 26602 8304 26608 8356
rect 26660 8344 26666 8356
rect 27172 8344 27200 8375
rect 27522 8372 27528 8384
rect 27580 8372 27586 8424
rect 27617 8415 27675 8421
rect 27617 8381 27629 8415
rect 27663 8412 27675 8415
rect 27709 8415 27767 8421
rect 27709 8412 27721 8415
rect 27663 8384 27721 8412
rect 27663 8381 27675 8384
rect 27617 8375 27675 8381
rect 27709 8381 27721 8384
rect 27755 8381 27767 8415
rect 27709 8375 27767 8381
rect 27632 8344 27660 8375
rect 28074 8372 28080 8424
rect 28132 8372 28138 8424
rect 28169 8415 28227 8421
rect 28169 8381 28181 8415
rect 28215 8412 28227 8415
rect 28276 8412 28304 8452
rect 28215 8384 28304 8412
rect 28215 8381 28227 8384
rect 28169 8375 28227 8381
rect 26660 8316 27660 8344
rect 26660 8304 26666 8316
rect 28276 8288 28304 8384
rect 28442 8372 28448 8424
rect 28500 8412 28506 8424
rect 28718 8412 28724 8424
rect 28500 8384 28724 8412
rect 28500 8372 28506 8384
rect 28718 8372 28724 8384
rect 28776 8412 28782 8424
rect 28813 8415 28871 8421
rect 28813 8412 28825 8415
rect 28776 8384 28825 8412
rect 28776 8372 28782 8384
rect 28813 8381 28825 8384
rect 28859 8381 28871 8415
rect 28813 8375 28871 8381
rect 28997 8415 29055 8421
rect 28997 8381 29009 8415
rect 29043 8412 29055 8415
rect 29270 8412 29276 8424
rect 29043 8384 29276 8412
rect 29043 8381 29055 8384
rect 28997 8375 29055 8381
rect 29270 8372 29276 8384
rect 29328 8372 29334 8424
rect 29380 8421 29408 8452
rect 29917 8449 29929 8483
rect 29963 8480 29975 8483
rect 30852 8480 30880 8520
rect 30929 8517 30941 8520
rect 30975 8517 30987 8551
rect 30929 8511 30987 8517
rect 29963 8452 30880 8480
rect 29963 8449 29975 8452
rect 29917 8443 29975 8449
rect 29365 8415 29423 8421
rect 29365 8381 29377 8415
rect 29411 8381 29423 8415
rect 29365 8375 29423 8381
rect 29454 8372 29460 8424
rect 29512 8412 29518 8424
rect 29822 8412 29828 8424
rect 29512 8384 29828 8412
rect 29512 8372 29518 8384
rect 29822 8372 29828 8384
rect 29880 8372 29886 8424
rect 30101 8415 30159 8421
rect 30101 8381 30113 8415
rect 30147 8412 30159 8415
rect 30282 8412 30288 8424
rect 30147 8384 30288 8412
rect 30147 8381 30159 8384
rect 30101 8375 30159 8381
rect 30282 8372 30288 8384
rect 30340 8372 30346 8424
rect 30561 8415 30619 8421
rect 30561 8381 30573 8415
rect 30607 8381 30619 8415
rect 30561 8375 30619 8381
rect 28905 8347 28963 8353
rect 28905 8313 28917 8347
rect 28951 8344 28963 8347
rect 29638 8344 29644 8356
rect 28951 8316 29644 8344
rect 28951 8313 28963 8316
rect 28905 8307 28963 8313
rect 29638 8304 29644 8316
rect 29696 8304 29702 8356
rect 30576 8288 30604 8375
rect 30650 8372 30656 8424
rect 30708 8372 30714 8424
rect 30745 8415 30803 8421
rect 30745 8381 30757 8415
rect 30791 8381 30803 8415
rect 30745 8375 30803 8381
rect 30760 8344 30788 8375
rect 30834 8372 30840 8424
rect 30892 8372 30898 8424
rect 31021 8415 31079 8421
rect 31021 8381 31033 8415
rect 31067 8412 31079 8415
rect 31110 8412 31116 8424
rect 31067 8384 31116 8412
rect 31067 8381 31079 8384
rect 31021 8375 31079 8381
rect 31110 8372 31116 8384
rect 31168 8372 31174 8424
rect 31202 8372 31208 8424
rect 31260 8412 31266 8424
rect 31386 8412 31392 8424
rect 31260 8384 31392 8412
rect 31260 8372 31266 8384
rect 31386 8372 31392 8384
rect 31444 8372 31450 8424
rect 31478 8372 31484 8424
rect 31536 8372 31542 8424
rect 31496 8344 31524 8372
rect 30760 8316 31524 8344
rect 23440 8248 24808 8276
rect 23440 8236 23446 8248
rect 25774 8236 25780 8288
rect 25832 8236 25838 8288
rect 26694 8236 26700 8288
rect 26752 8236 26758 8288
rect 26789 8279 26847 8285
rect 26789 8245 26801 8279
rect 26835 8276 26847 8279
rect 27430 8276 27436 8288
rect 26835 8248 27436 8276
rect 26835 8245 26847 8248
rect 26789 8239 26847 8245
rect 27430 8236 27436 8248
rect 27488 8236 27494 8288
rect 28258 8236 28264 8288
rect 28316 8236 28322 8288
rect 28718 8236 28724 8288
rect 28776 8236 28782 8288
rect 28810 8236 28816 8288
rect 28868 8276 28874 8288
rect 29273 8279 29331 8285
rect 29273 8276 29285 8279
rect 28868 8248 29285 8276
rect 28868 8236 28874 8248
rect 29273 8245 29285 8248
rect 29319 8245 29331 8279
rect 29273 8239 29331 8245
rect 29454 8236 29460 8288
rect 29512 8236 29518 8288
rect 30009 8279 30067 8285
rect 30009 8245 30021 8279
rect 30055 8276 30067 8279
rect 30466 8276 30472 8288
rect 30055 8248 30472 8276
rect 30055 8245 30067 8248
rect 30009 8239 30067 8245
rect 30466 8236 30472 8248
rect 30524 8236 30530 8288
rect 30558 8236 30564 8288
rect 30616 8276 30622 8288
rect 31665 8279 31723 8285
rect 31665 8276 31677 8279
rect 30616 8248 31677 8276
rect 30616 8236 30622 8248
rect 31665 8245 31677 8248
rect 31711 8245 31723 8279
rect 31665 8239 31723 8245
rect 2760 8186 32200 8208
rect 2760 8134 6946 8186
rect 6998 8134 7010 8186
rect 7062 8134 7074 8186
rect 7126 8134 7138 8186
rect 7190 8134 7202 8186
rect 7254 8134 14306 8186
rect 14358 8134 14370 8186
rect 14422 8134 14434 8186
rect 14486 8134 14498 8186
rect 14550 8134 14562 8186
rect 14614 8134 21666 8186
rect 21718 8134 21730 8186
rect 21782 8134 21794 8186
rect 21846 8134 21858 8186
rect 21910 8134 21922 8186
rect 21974 8134 29026 8186
rect 29078 8134 29090 8186
rect 29142 8134 29154 8186
rect 29206 8134 29218 8186
rect 29270 8134 29282 8186
rect 29334 8134 32200 8186
rect 2760 8112 32200 8134
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 14182 8072 14188 8084
rect 3292 8044 14188 8072
rect 3292 8032 3298 8044
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 16224 8044 16804 8072
rect 6181 8007 6239 8013
rect 6181 8004 6193 8007
rect 5290 7976 6193 8004
rect 6181 7973 6193 7976
rect 6227 7973 6239 8007
rect 6181 7967 6239 7973
rect 1302 7896 1308 7948
rect 1360 7936 1366 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 1360 7908 3065 7936
rect 1360 7896 1366 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 6273 7939 6331 7945
rect 6273 7905 6285 7939
rect 6319 7936 6331 7939
rect 6319 7908 6868 7936
rect 6319 7905 6331 7908
rect 6273 7899 6331 7905
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 5997 7871 6055 7877
rect 5767 7840 5948 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 5920 7800 5948 7840
rect 5997 7837 6009 7871
rect 6043 7868 6055 7871
rect 6086 7868 6092 7880
rect 6043 7840 6092 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6086 7828 6092 7840
rect 6144 7828 6150 7880
rect 6178 7828 6184 7880
rect 6236 7828 6242 7880
rect 6196 7800 6224 7828
rect 6840 7812 6868 7908
rect 14182 7896 14188 7948
rect 14240 7945 14246 7948
rect 14240 7939 14268 7945
rect 14256 7905 14268 7939
rect 14240 7899 14268 7905
rect 14240 7896 14246 7899
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16224 7945 16252 8044
rect 16776 8016 16804 8044
rect 18046 8032 18052 8084
rect 18104 8072 18110 8084
rect 18141 8075 18199 8081
rect 18141 8072 18153 8075
rect 18104 8044 18153 8072
rect 18104 8032 18110 8044
rect 18141 8041 18153 8044
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 18969 8075 19027 8081
rect 18969 8041 18981 8075
rect 19015 8072 19027 8075
rect 19242 8072 19248 8084
rect 19015 8044 19248 8072
rect 19015 8041 19027 8044
rect 18969 8035 19027 8041
rect 19242 8032 19248 8044
rect 19300 8032 19306 8084
rect 22189 8075 22247 8081
rect 22189 8041 22201 8075
rect 22235 8041 22247 8075
rect 22189 8035 22247 8041
rect 22833 8075 22891 8081
rect 22833 8041 22845 8075
rect 22879 8072 22891 8075
rect 23290 8072 23296 8084
rect 22879 8044 23296 8072
rect 22879 8041 22891 8044
rect 22833 8035 22891 8041
rect 16574 7964 16580 8016
rect 16632 8004 16638 8016
rect 16669 8007 16727 8013
rect 16669 8004 16681 8007
rect 16632 7976 16681 8004
rect 16632 7964 16638 7976
rect 16669 7973 16681 7976
rect 16715 7973 16727 8007
rect 16669 7967 16727 7973
rect 16758 7964 16764 8016
rect 16816 7964 16822 8016
rect 18414 8004 18420 8016
rect 17894 7976 18420 8004
rect 18414 7964 18420 7976
rect 18472 7964 18478 8016
rect 20993 8007 21051 8013
rect 20993 7973 21005 8007
rect 21039 8004 21051 8007
rect 21821 8007 21879 8013
rect 21821 8004 21833 8007
rect 21039 7976 21833 8004
rect 21039 7973 21051 7976
rect 20993 7967 21051 7973
rect 21821 7973 21833 7976
rect 21867 7973 21879 8007
rect 21821 7967 21879 7973
rect 21913 8007 21971 8013
rect 21913 7973 21925 8007
rect 21959 8004 21971 8007
rect 22094 8004 22100 8016
rect 21959 7976 22100 8004
rect 21959 7973 21971 7976
rect 21913 7967 21971 7973
rect 22094 7964 22100 7976
rect 22152 7964 22158 8016
rect 22204 8004 22232 8035
rect 23290 8032 23296 8044
rect 23348 8032 23354 8084
rect 25041 8075 25099 8081
rect 25041 8041 25053 8075
rect 25087 8072 25099 8075
rect 26418 8072 26424 8084
rect 25087 8044 26424 8072
rect 25087 8041 25099 8044
rect 25041 8035 25099 8041
rect 26418 8032 26424 8044
rect 26476 8032 26482 8084
rect 26694 8072 26700 8084
rect 26528 8044 26700 8072
rect 22204 7976 22784 8004
rect 15841 7939 15899 7945
rect 15841 7936 15853 7939
rect 15804 7908 15853 7936
rect 15804 7896 15810 7908
rect 15841 7905 15853 7908
rect 15887 7905 15899 7939
rect 15841 7899 15899 7905
rect 16209 7939 16267 7945
rect 16209 7905 16221 7939
rect 16255 7905 16267 7939
rect 16209 7899 16267 7905
rect 18322 7896 18328 7948
rect 18380 7936 18386 7948
rect 19153 7939 19211 7945
rect 19153 7936 19165 7939
rect 18380 7908 19165 7936
rect 18380 7896 18386 7908
rect 19153 7905 19165 7908
rect 19199 7905 19211 7939
rect 19153 7899 19211 7905
rect 20162 7896 20168 7948
rect 20220 7945 20226 7948
rect 20220 7939 20248 7945
rect 20236 7905 20248 7939
rect 20220 7899 20248 7905
rect 20220 7896 20226 7899
rect 20346 7896 20352 7948
rect 20404 7896 20410 7948
rect 21637 7939 21695 7945
rect 21637 7905 21649 7939
rect 21683 7905 21695 7939
rect 21637 7899 21695 7905
rect 22005 7939 22063 7945
rect 22005 7905 22017 7939
rect 22051 7936 22063 7939
rect 22051 7908 22324 7936
rect 22051 7905 22063 7908
rect 22005 7899 22063 7905
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 13964 7840 14105 7868
rect 13964 7828 13970 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14369 7871 14427 7877
rect 14369 7837 14381 7871
rect 14415 7868 14427 7871
rect 14415 7840 14872 7868
rect 14415 7837 14427 7840
rect 14369 7831 14427 7837
rect 3283 7772 4752 7800
rect 5920 7772 6224 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 4246 7692 4252 7744
rect 4304 7692 4310 7744
rect 4724 7732 4752 7772
rect 6822 7760 6828 7812
rect 6880 7760 6886 7812
rect 13817 7803 13875 7809
rect 13817 7769 13829 7803
rect 13863 7769 13875 7803
rect 13817 7763 13875 7769
rect 13722 7732 13728 7744
rect 4724 7704 13728 7732
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 13832 7732 13860 7763
rect 14844 7744 14872 7840
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 16117 7871 16175 7877
rect 16117 7868 16129 7871
rect 15252 7840 16129 7868
rect 15252 7828 15258 7840
rect 16117 7837 16129 7840
rect 16163 7837 16175 7871
rect 16117 7831 16175 7837
rect 16390 7828 16396 7880
rect 16448 7828 16454 7880
rect 19334 7828 19340 7880
rect 19392 7828 19398 7880
rect 20070 7828 20076 7880
rect 20128 7828 20134 7880
rect 21652 7868 21680 7899
rect 21910 7868 21916 7880
rect 21652 7840 21916 7868
rect 21910 7828 21916 7840
rect 21968 7828 21974 7880
rect 15013 7803 15071 7809
rect 15013 7769 15025 7803
rect 15059 7800 15071 7803
rect 15562 7800 15568 7812
rect 15059 7772 15568 7800
rect 15059 7769 15071 7772
rect 15013 7763 15071 7769
rect 15562 7760 15568 7772
rect 15620 7760 15626 7812
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7769 19855 7803
rect 19797 7763 19855 7769
rect 14182 7732 14188 7744
rect 13832 7704 14188 7732
rect 14182 7692 14188 7704
rect 14240 7732 14246 7744
rect 14734 7732 14740 7744
rect 14240 7704 14740 7732
rect 14240 7692 14246 7704
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 14826 7692 14832 7744
rect 14884 7692 14890 7744
rect 15286 7692 15292 7744
rect 15344 7692 15350 7744
rect 19812 7732 19840 7763
rect 20898 7732 20904 7744
rect 19812 7704 20904 7732
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 21928 7732 21956 7828
rect 22296 7809 22324 7908
rect 22554 7896 22560 7948
rect 22612 7896 22618 7948
rect 22756 7945 22784 7976
rect 25774 7964 25780 8016
rect 25832 7964 25838 8016
rect 26528 8013 26556 8044
rect 26694 8032 26700 8044
rect 26752 8032 26758 8084
rect 28074 8032 28080 8084
rect 28132 8072 28138 8084
rect 28261 8075 28319 8081
rect 28261 8072 28273 8075
rect 28132 8044 28273 8072
rect 28132 8032 28138 8044
rect 28261 8041 28273 8044
rect 28307 8041 28319 8075
rect 28261 8035 28319 8041
rect 28718 8032 28724 8084
rect 28776 8072 28782 8084
rect 29914 8072 29920 8084
rect 28776 8044 29920 8072
rect 28776 8032 28782 8044
rect 26513 8007 26571 8013
rect 26513 7973 26525 8007
rect 26559 7973 26571 8007
rect 26513 7967 26571 7973
rect 27632 7976 28948 8004
rect 27632 7948 27660 7976
rect 22649 7939 22707 7945
rect 22649 7905 22661 7939
rect 22695 7905 22707 7939
rect 22649 7899 22707 7905
rect 22741 7939 22799 7945
rect 22741 7905 22753 7939
rect 22787 7905 22799 7939
rect 22741 7899 22799 7905
rect 22925 7939 22983 7945
rect 22925 7905 22937 7939
rect 22971 7936 22983 7939
rect 23014 7936 23020 7948
rect 22971 7908 23020 7936
rect 22971 7905 22983 7908
rect 22925 7899 22983 7905
rect 22664 7868 22692 7899
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 23106 7896 23112 7948
rect 23164 7936 23170 7948
rect 23661 7939 23719 7945
rect 23661 7936 23673 7939
rect 23164 7908 23673 7936
rect 23164 7896 23170 7908
rect 23661 7905 23673 7908
rect 23707 7905 23719 7939
rect 23661 7899 23719 7905
rect 24397 7939 24455 7945
rect 24397 7905 24409 7939
rect 24443 7936 24455 7939
rect 24762 7936 24768 7948
rect 24443 7908 24768 7936
rect 24443 7905 24455 7908
rect 24397 7899 24455 7905
rect 23474 7868 23480 7880
rect 22664 7840 23480 7868
rect 23474 7828 23480 7840
rect 23532 7828 23538 7880
rect 22281 7803 22339 7809
rect 22281 7769 22293 7803
rect 22327 7769 22339 7803
rect 22281 7763 22339 7769
rect 22922 7760 22928 7812
rect 22980 7800 22986 7812
rect 24412 7800 24440 7899
rect 24762 7896 24768 7908
rect 24820 7896 24826 7948
rect 27614 7896 27620 7948
rect 27672 7896 27678 7948
rect 28166 7896 28172 7948
rect 28224 7936 28230 7948
rect 28920 7945 28948 7976
rect 29104 7945 29132 8044
rect 29914 8032 29920 8044
rect 29972 8072 29978 8084
rect 30558 8072 30564 8084
rect 29972 8044 30564 8072
rect 29972 8032 29978 8044
rect 30558 8032 30564 8044
rect 30616 8032 30622 8084
rect 31021 8075 31079 8081
rect 31021 8041 31033 8075
rect 31067 8072 31079 8075
rect 31110 8072 31116 8084
rect 31067 8044 31116 8072
rect 31067 8041 31079 8044
rect 31021 8035 31079 8041
rect 29454 7964 29460 8016
rect 29512 8004 29518 8016
rect 30374 8004 30380 8016
rect 29512 7976 30380 8004
rect 29512 7964 29518 7976
rect 30374 7964 30380 7976
rect 30432 8004 30438 8016
rect 31036 8004 31064 8035
rect 31110 8032 31116 8044
rect 31168 8032 31174 8084
rect 30432 7976 31064 8004
rect 30432 7964 30438 7976
rect 28813 7939 28871 7945
rect 28813 7936 28825 7939
rect 28224 7908 28825 7936
rect 28224 7896 28230 7908
rect 28813 7905 28825 7908
rect 28859 7905 28871 7939
rect 28813 7899 28871 7905
rect 28905 7939 28963 7945
rect 28905 7905 28917 7939
rect 28951 7905 28963 7939
rect 28905 7899 28963 7905
rect 29089 7939 29147 7945
rect 29089 7905 29101 7939
rect 29135 7905 29147 7939
rect 29089 7899 29147 7905
rect 26789 7871 26847 7877
rect 26789 7837 26801 7871
rect 26835 7837 26847 7871
rect 26789 7831 26847 7837
rect 22980 7772 24440 7800
rect 22980 7760 22986 7772
rect 22462 7732 22468 7744
rect 21928 7704 22468 7732
rect 22462 7692 22468 7704
rect 22520 7692 22526 7744
rect 24118 7692 24124 7744
rect 24176 7732 24182 7744
rect 24305 7735 24363 7741
rect 24305 7732 24317 7735
rect 24176 7704 24317 7732
rect 24176 7692 24182 7704
rect 24305 7701 24317 7704
rect 24351 7701 24363 7735
rect 24305 7695 24363 7701
rect 24486 7692 24492 7744
rect 24544 7692 24550 7744
rect 26326 7692 26332 7744
rect 26384 7732 26390 7744
rect 26804 7732 26832 7831
rect 27430 7828 27436 7880
rect 27488 7828 27494 7880
rect 27706 7828 27712 7880
rect 27764 7828 27770 7880
rect 27798 7828 27804 7880
rect 27856 7868 27862 7880
rect 29472 7877 29500 7964
rect 29641 7939 29699 7945
rect 29641 7905 29653 7939
rect 29687 7936 29699 7939
rect 29730 7936 29736 7948
rect 29687 7908 29736 7936
rect 29687 7905 29699 7908
rect 29641 7899 29699 7905
rect 29730 7896 29736 7908
rect 29788 7936 29794 7948
rect 30742 7936 30748 7948
rect 29788 7908 30748 7936
rect 29788 7896 29794 7908
rect 30742 7896 30748 7908
rect 30800 7896 30806 7948
rect 30834 7896 30840 7948
rect 30892 7896 30898 7948
rect 31849 7939 31907 7945
rect 31849 7905 31861 7939
rect 31895 7936 31907 7939
rect 33134 7936 33140 7948
rect 31895 7908 33140 7936
rect 31895 7905 31907 7908
rect 31849 7899 31907 7905
rect 33134 7896 33140 7908
rect 33192 7896 33198 7948
rect 28997 7871 29055 7877
rect 28997 7868 29009 7871
rect 27856 7840 29009 7868
rect 27856 7828 27862 7840
rect 28997 7837 29009 7840
rect 29043 7837 29055 7871
rect 28997 7831 29055 7837
rect 29457 7871 29515 7877
rect 29457 7837 29469 7871
rect 29503 7837 29515 7871
rect 29457 7831 29515 7837
rect 29549 7871 29607 7877
rect 29549 7837 29561 7871
rect 29595 7837 29607 7871
rect 29549 7831 29607 7837
rect 30653 7871 30711 7877
rect 30653 7837 30665 7871
rect 30699 7837 30711 7871
rect 30653 7831 30711 7837
rect 26970 7760 26976 7812
rect 27028 7800 27034 7812
rect 27028 7772 28994 7800
rect 27028 7760 27034 7772
rect 26384 7704 26832 7732
rect 26384 7692 26390 7704
rect 26878 7692 26884 7744
rect 26936 7692 26942 7744
rect 28718 7692 28724 7744
rect 28776 7692 28782 7744
rect 28966 7732 28994 7772
rect 29454 7732 29460 7744
rect 28966 7704 29460 7732
rect 29454 7692 29460 7704
rect 29512 7692 29518 7744
rect 29564 7732 29592 7831
rect 30009 7803 30067 7809
rect 30009 7769 30021 7803
rect 30055 7800 30067 7803
rect 30668 7800 30696 7831
rect 30055 7772 30696 7800
rect 30055 7769 30067 7772
rect 30009 7763 30067 7769
rect 29638 7732 29644 7744
rect 29564 7704 29644 7732
rect 29638 7692 29644 7704
rect 29696 7692 29702 7744
rect 30098 7692 30104 7744
rect 30156 7692 30162 7744
rect 31662 7692 31668 7744
rect 31720 7692 31726 7744
rect 2760 7642 32200 7664
rect 2760 7590 6286 7642
rect 6338 7590 6350 7642
rect 6402 7590 6414 7642
rect 6466 7590 6478 7642
rect 6530 7590 6542 7642
rect 6594 7590 13646 7642
rect 13698 7590 13710 7642
rect 13762 7590 13774 7642
rect 13826 7590 13838 7642
rect 13890 7590 13902 7642
rect 13954 7590 21006 7642
rect 21058 7590 21070 7642
rect 21122 7590 21134 7642
rect 21186 7590 21198 7642
rect 21250 7590 21262 7642
rect 21314 7590 28366 7642
rect 28418 7590 28430 7642
rect 28482 7590 28494 7642
rect 28546 7590 28558 7642
rect 28610 7590 28622 7642
rect 28674 7590 32200 7642
rect 2760 7568 32200 7590
rect 7650 7488 7656 7540
rect 7708 7528 7714 7540
rect 9398 7528 9404 7540
rect 7708 7500 9404 7528
rect 7708 7488 7714 7500
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13630 7528 13636 7540
rect 13320 7500 13636 7528
rect 13320 7488 13326 7500
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 14080 7531 14138 7537
rect 14080 7497 14092 7531
rect 14126 7528 14138 7531
rect 15286 7528 15292 7540
rect 14126 7500 15292 7528
rect 14126 7497 14138 7500
rect 14080 7491 14138 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 15749 7531 15807 7537
rect 15749 7528 15761 7531
rect 15396 7500 15761 7528
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 15396 7460 15424 7500
rect 15749 7497 15761 7500
rect 15795 7497 15807 7531
rect 15749 7491 15807 7497
rect 16577 7531 16635 7537
rect 16577 7497 16589 7531
rect 16623 7528 16635 7531
rect 16666 7528 16672 7540
rect 16623 7500 16672 7528
rect 16623 7497 16635 7500
rect 16577 7491 16635 7497
rect 16666 7488 16672 7500
rect 16724 7488 16730 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18141 7531 18199 7537
rect 18141 7528 18153 7531
rect 18012 7500 18153 7528
rect 18012 7488 18018 7500
rect 18141 7497 18153 7500
rect 18187 7497 18199 7531
rect 18141 7491 18199 7497
rect 18230 7488 18236 7540
rect 18288 7528 18294 7540
rect 18417 7531 18475 7537
rect 18417 7528 18429 7531
rect 18288 7500 18429 7528
rect 18288 7488 18294 7500
rect 18417 7497 18429 7500
rect 18463 7497 18475 7531
rect 22554 7528 22560 7540
rect 18417 7491 18475 7497
rect 18524 7500 22560 7528
rect 18524 7460 18552 7500
rect 22554 7488 22560 7500
rect 22612 7488 22618 7540
rect 23382 7488 23388 7540
rect 23440 7488 23446 7540
rect 27706 7488 27712 7540
rect 27764 7528 27770 7540
rect 27801 7531 27859 7537
rect 27801 7528 27813 7531
rect 27764 7500 27813 7528
rect 27764 7488 27770 7500
rect 27801 7497 27813 7500
rect 27847 7497 27859 7531
rect 27801 7491 27859 7497
rect 28718 7488 28724 7540
rect 28776 7488 28782 7540
rect 28813 7531 28871 7537
rect 28813 7497 28825 7531
rect 28859 7528 28871 7531
rect 28902 7528 28908 7540
rect 28859 7500 28908 7528
rect 28859 7497 28871 7500
rect 28813 7491 28871 7497
rect 15160 7432 15424 7460
rect 15488 7432 18552 7460
rect 15160 7420 15166 7432
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7361 13875 7395
rect 13817 7355 13875 7361
rect 13832 7256 13860 7355
rect 15194 7284 15200 7336
rect 15252 7284 15258 7336
rect 14090 7256 14096 7268
rect 13832 7228 14096 7256
rect 14090 7216 14096 7228
rect 14148 7216 14154 7268
rect 13170 7148 13176 7200
rect 13228 7188 13234 7200
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 13228 7160 13737 7188
rect 13228 7148 13234 7160
rect 13725 7157 13737 7160
rect 13771 7188 13783 7191
rect 15488 7188 15516 7432
rect 15565 7395 15623 7401
rect 15565 7361 15577 7395
rect 15611 7392 15623 7395
rect 17497 7395 17555 7401
rect 17497 7392 17509 7395
rect 15611 7364 17509 7392
rect 15611 7361 15623 7364
rect 15565 7355 15623 7361
rect 17497 7361 17509 7364
rect 17543 7361 17555 7395
rect 17497 7355 17555 7361
rect 21450 7352 21456 7404
rect 21508 7392 21514 7404
rect 21637 7395 21695 7401
rect 21637 7392 21649 7395
rect 21508 7364 21649 7392
rect 21508 7352 21514 7364
rect 21637 7361 21649 7364
rect 21683 7392 21695 7395
rect 21910 7392 21916 7404
rect 21683 7364 21916 7392
rect 21683 7361 21695 7364
rect 21637 7355 21695 7361
rect 21910 7352 21916 7364
rect 21968 7352 21974 7404
rect 23753 7395 23811 7401
rect 23753 7361 23765 7395
rect 23799 7392 23811 7395
rect 26053 7395 26111 7401
rect 26053 7392 26065 7395
rect 23799 7364 26065 7392
rect 23799 7361 23811 7364
rect 23753 7355 23811 7361
rect 26053 7361 26065 7364
rect 26099 7361 26111 7395
rect 28736 7392 28764 7488
rect 26053 7355 26111 7361
rect 27448 7364 28764 7392
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7293 16359 7327
rect 16301 7287 16359 7293
rect 16669 7327 16727 7333
rect 16669 7293 16681 7327
rect 16715 7324 16727 7327
rect 16758 7324 16764 7336
rect 16715 7296 16764 7324
rect 16715 7293 16727 7296
rect 16669 7287 16727 7293
rect 15654 7216 15660 7268
rect 15712 7256 15718 7268
rect 16316 7256 16344 7287
rect 16758 7284 16764 7296
rect 16816 7324 16822 7336
rect 17034 7324 17040 7336
rect 16816 7296 17040 7324
rect 16816 7284 16822 7296
rect 17034 7284 17040 7296
rect 17092 7284 17098 7336
rect 17310 7284 17316 7336
rect 17368 7284 17374 7336
rect 18506 7324 18512 7336
rect 18248 7296 18512 7324
rect 18248 7268 18276 7296
rect 18506 7284 18512 7296
rect 18564 7284 18570 7336
rect 24118 7284 24124 7336
rect 24176 7284 24182 7336
rect 15712 7228 16344 7256
rect 15712 7216 15718 7228
rect 18230 7216 18236 7268
rect 18288 7216 18294 7268
rect 21913 7259 21971 7265
rect 21913 7225 21925 7259
rect 21959 7256 21971 7259
rect 22186 7256 22192 7268
rect 21959 7228 22192 7256
rect 21959 7225 21971 7228
rect 21913 7219 21971 7225
rect 22186 7216 22192 7228
rect 22244 7216 22250 7268
rect 22646 7216 22652 7268
rect 22704 7216 22710 7268
rect 24486 7216 24492 7268
rect 24544 7216 24550 7268
rect 26068 7256 26096 7355
rect 27448 7310 27476 7364
rect 28258 7284 28264 7336
rect 28316 7324 28322 7336
rect 28316 7296 28396 7324
rect 28316 7284 28322 7296
rect 26234 7256 26240 7268
rect 25240 7228 25912 7256
rect 26068 7228 26240 7256
rect 13771 7160 15516 7188
rect 13771 7157 13783 7160
rect 13725 7151 13783 7157
rect 16758 7148 16764 7200
rect 16816 7148 16822 7200
rect 20438 7148 20444 7200
rect 20496 7188 20502 7200
rect 20625 7191 20683 7197
rect 20625 7188 20637 7191
rect 20496 7160 20637 7188
rect 20496 7148 20502 7160
rect 20625 7157 20637 7160
rect 20671 7157 20683 7191
rect 20625 7151 20683 7157
rect 22554 7148 22560 7200
rect 22612 7188 22618 7200
rect 25240 7188 25268 7228
rect 22612 7160 25268 7188
rect 22612 7148 22618 7160
rect 25314 7148 25320 7200
rect 25372 7188 25378 7200
rect 25547 7191 25605 7197
rect 25547 7188 25559 7191
rect 25372 7160 25559 7188
rect 25372 7148 25378 7160
rect 25547 7157 25559 7160
rect 25593 7188 25605 7191
rect 25774 7188 25780 7200
rect 25593 7160 25780 7188
rect 25593 7157 25605 7160
rect 25547 7151 25605 7157
rect 25774 7148 25780 7160
rect 25832 7148 25838 7200
rect 25884 7188 25912 7228
rect 26234 7216 26240 7228
rect 26292 7216 26298 7268
rect 26326 7216 26332 7268
rect 26384 7216 26390 7268
rect 27614 7216 27620 7268
rect 27672 7256 27678 7268
rect 28368 7256 28396 7296
rect 28442 7284 28448 7336
rect 28500 7284 28506 7336
rect 28828 7324 28856 7491
rect 28902 7488 28908 7500
rect 28960 7488 28966 7540
rect 29352 7531 29410 7537
rect 29352 7497 29364 7531
rect 29398 7528 29410 7531
rect 30098 7528 30104 7540
rect 29398 7500 30104 7528
rect 29398 7497 29410 7500
rect 29352 7491 29410 7497
rect 30098 7488 30104 7500
rect 30156 7488 30162 7540
rect 30834 7488 30840 7540
rect 30892 7488 30898 7540
rect 29362 7392 29368 7404
rect 29104 7364 29368 7392
rect 28552 7296 28856 7324
rect 28552 7256 28580 7296
rect 28994 7284 29000 7336
rect 29052 7324 29058 7336
rect 29104 7333 29132 7364
rect 29362 7352 29368 7364
rect 29420 7352 29426 7404
rect 29089 7327 29147 7333
rect 29089 7324 29101 7327
rect 29052 7296 29101 7324
rect 29052 7284 29058 7296
rect 29089 7293 29101 7296
rect 29135 7293 29147 7327
rect 29089 7287 29147 7293
rect 30466 7284 30472 7336
rect 30524 7284 30530 7336
rect 27672 7228 28304 7256
rect 28368 7228 28580 7256
rect 28629 7259 28687 7265
rect 27672 7216 27678 7228
rect 26970 7188 26976 7200
rect 25884 7160 26976 7188
rect 26970 7148 26976 7160
rect 27028 7148 27034 7200
rect 27246 7148 27252 7200
rect 27304 7188 27310 7200
rect 27893 7191 27951 7197
rect 27893 7188 27905 7191
rect 27304 7160 27905 7188
rect 27304 7148 27310 7160
rect 27893 7157 27905 7160
rect 27939 7157 27951 7191
rect 28276 7188 28304 7228
rect 28629 7225 28641 7259
rect 28675 7256 28687 7259
rect 28718 7256 28724 7268
rect 28675 7228 28724 7256
rect 28675 7225 28687 7228
rect 28629 7219 28687 7225
rect 28718 7216 28724 7228
rect 28776 7216 28782 7268
rect 28829 7191 28887 7197
rect 28829 7188 28841 7191
rect 28276 7160 28841 7188
rect 27893 7151 27951 7157
rect 28829 7157 28841 7160
rect 28875 7157 28887 7191
rect 28829 7151 28887 7157
rect 28997 7191 29055 7197
rect 28997 7157 29009 7191
rect 29043 7188 29055 7191
rect 29362 7188 29368 7200
rect 29043 7160 29368 7188
rect 29043 7157 29055 7160
rect 28997 7151 29055 7157
rect 29362 7148 29368 7160
rect 29420 7188 29426 7200
rect 29730 7188 29736 7200
rect 29420 7160 29736 7188
rect 29420 7148 29426 7160
rect 29730 7148 29736 7160
rect 29788 7148 29794 7200
rect 2760 7098 32200 7120
rect 2760 7046 6946 7098
rect 6998 7046 7010 7098
rect 7062 7046 7074 7098
rect 7126 7046 7138 7098
rect 7190 7046 7202 7098
rect 7254 7046 14306 7098
rect 14358 7046 14370 7098
rect 14422 7046 14434 7098
rect 14486 7046 14498 7098
rect 14550 7046 14562 7098
rect 14614 7046 21666 7098
rect 21718 7046 21730 7098
rect 21782 7046 21794 7098
rect 21846 7046 21858 7098
rect 21910 7046 21922 7098
rect 21974 7046 29026 7098
rect 29078 7046 29090 7098
rect 29142 7046 29154 7098
rect 29206 7046 29218 7098
rect 29270 7046 29282 7098
rect 29334 7046 32200 7098
rect 2760 7024 32200 7046
rect 13538 6984 13544 6996
rect 12452 6956 13544 6984
rect 7285 6919 7343 6925
rect 7285 6885 7297 6919
rect 7331 6916 7343 6919
rect 7650 6916 7656 6928
rect 7331 6888 7656 6916
rect 7331 6885 7343 6888
rect 7285 6879 7343 6885
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 8297 6919 8355 6925
rect 8297 6885 8309 6919
rect 8343 6916 8355 6919
rect 8343 6888 9674 6916
rect 8343 6885 8355 6888
rect 8297 6879 8355 6885
rect 7101 6851 7159 6857
rect 7101 6817 7113 6851
rect 7147 6817 7159 6851
rect 7101 6811 7159 6817
rect 7116 6780 7144 6811
rect 7190 6808 7196 6860
rect 7248 6808 7254 6860
rect 7469 6851 7527 6857
rect 7469 6817 7481 6851
rect 7515 6848 7527 6851
rect 8312 6848 8340 6879
rect 7515 6820 8340 6848
rect 9646 6848 9674 6888
rect 11882 6848 11888 6860
rect 9646 6820 11888 6848
rect 7515 6817 7527 6820
rect 7469 6811 7527 6817
rect 11882 6808 11888 6820
rect 11940 6808 11946 6860
rect 7116 6752 7788 6780
rect 6914 6604 6920 6656
rect 6972 6604 6978 6656
rect 7760 6653 7788 6752
rect 9398 6740 9404 6792
rect 9456 6780 9462 6792
rect 12452 6780 12480 6956
rect 13538 6944 13544 6956
rect 13596 6984 13602 6996
rect 15470 6984 15476 6996
rect 13596 6956 15476 6984
rect 13596 6944 13602 6956
rect 15470 6944 15476 6956
rect 15528 6944 15534 6996
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 16117 6987 16175 6993
rect 16117 6984 16129 6987
rect 15620 6956 16129 6984
rect 15620 6944 15626 6956
rect 16117 6953 16129 6956
rect 16163 6953 16175 6987
rect 16117 6947 16175 6953
rect 16298 6944 16304 6996
rect 16356 6944 16362 6996
rect 19334 6944 19340 6996
rect 19392 6984 19398 6996
rect 20165 6987 20223 6993
rect 20165 6984 20177 6987
rect 19392 6956 20177 6984
rect 19392 6944 19398 6956
rect 20165 6953 20177 6956
rect 20211 6984 20223 6987
rect 20625 6987 20683 6993
rect 20625 6984 20637 6987
rect 20211 6956 20637 6984
rect 20211 6953 20223 6956
rect 20165 6947 20223 6953
rect 20625 6953 20637 6956
rect 20671 6953 20683 6987
rect 20625 6947 20683 6953
rect 22646 6944 22652 6996
rect 22704 6984 22710 6996
rect 22741 6987 22799 6993
rect 22741 6984 22753 6987
rect 22704 6956 22753 6984
rect 22704 6944 22710 6956
rect 22741 6953 22753 6956
rect 22787 6953 22799 6987
rect 22741 6947 22799 6953
rect 23474 6944 23480 6996
rect 23532 6944 23538 6996
rect 26326 6944 26332 6996
rect 26384 6984 26390 6996
rect 26513 6987 26571 6993
rect 26513 6984 26525 6987
rect 26384 6956 26525 6984
rect 26384 6944 26390 6956
rect 26513 6953 26525 6956
rect 26559 6953 26571 6987
rect 26513 6947 26571 6953
rect 26878 6944 26884 6996
rect 26936 6944 26942 6996
rect 27614 6944 27620 6996
rect 27672 6944 27678 6996
rect 27798 6944 27804 6996
rect 27856 6944 27862 6996
rect 27985 6987 28043 6993
rect 27985 6953 27997 6987
rect 28031 6984 28043 6987
rect 28350 6984 28356 6996
rect 28031 6956 28356 6984
rect 28031 6953 28043 6956
rect 27985 6947 28043 6953
rect 28350 6944 28356 6956
rect 28408 6944 28414 6996
rect 28718 6984 28724 6996
rect 28460 6956 28724 6984
rect 12526 6876 12532 6928
rect 12584 6916 12590 6928
rect 15194 6916 15200 6928
rect 12584 6888 15200 6916
rect 12584 6876 12590 6888
rect 15194 6876 15200 6888
rect 15252 6876 15258 6928
rect 15378 6876 15384 6928
rect 15436 6876 15442 6928
rect 16669 6919 16727 6925
rect 16669 6885 16681 6919
rect 16715 6916 16727 6919
rect 16758 6916 16764 6928
rect 16715 6888 16764 6916
rect 16715 6885 16727 6888
rect 16669 6879 16727 6885
rect 16758 6876 16764 6888
rect 16816 6876 16822 6928
rect 20070 6876 20076 6928
rect 20128 6876 20134 6928
rect 22922 6916 22928 6928
rect 22664 6888 22928 6916
rect 13262 6848 13268 6860
rect 13096 6820 13268 6848
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 9456 6752 12541 6780
rect 9456 6740 9462 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 12529 6743 12587 6749
rect 7745 6647 7803 6653
rect 7745 6613 7757 6647
rect 7791 6644 7803 6647
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 7791 6616 12909 6644
rect 7791 6613 7803 6616
rect 7745 6607 7803 6613
rect 12897 6613 12909 6616
rect 12943 6644 12955 6647
rect 13096 6644 13124 6820
rect 13262 6808 13268 6820
rect 13320 6848 13326 6860
rect 13357 6851 13415 6857
rect 13357 6848 13369 6851
rect 13320 6820 13369 6848
rect 13320 6808 13326 6820
rect 13357 6817 13369 6820
rect 13403 6817 13415 6851
rect 13357 6811 13415 6817
rect 13446 6808 13452 6860
rect 13504 6808 13510 6860
rect 13538 6808 13544 6860
rect 13596 6808 13602 6860
rect 13630 6808 13636 6860
rect 13688 6848 13694 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13688 6820 13737 6848
rect 13688 6808 13694 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 14461 6851 14519 6857
rect 14461 6817 14473 6851
rect 14507 6817 14519 6851
rect 14461 6811 14519 6817
rect 14553 6851 14611 6857
rect 14553 6817 14565 6851
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 14476 6712 14504 6811
rect 14568 6780 14596 6811
rect 14642 6808 14648 6860
rect 14700 6848 14706 6860
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 14700 6820 14749 6848
rect 14700 6808 14706 6820
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 14737 6811 14795 6817
rect 14918 6808 14924 6860
rect 14976 6808 14982 6860
rect 15010 6808 15016 6860
rect 15068 6808 15074 6860
rect 15212 6848 15240 6876
rect 16390 6848 16396 6860
rect 15212 6820 16396 6848
rect 16390 6808 16396 6820
rect 16448 6808 16454 6860
rect 18414 6848 18420 6860
rect 17802 6820 18420 6848
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18969 6851 19027 6857
rect 18969 6817 18981 6851
rect 19015 6848 19027 6851
rect 20088 6848 20116 6876
rect 19015 6820 20116 6848
rect 20257 6851 20315 6857
rect 19015 6817 19027 6820
rect 18969 6811 19027 6817
rect 20257 6817 20269 6851
rect 20303 6848 20315 6851
rect 20622 6848 20628 6860
rect 20303 6820 20628 6848
rect 20303 6817 20315 6820
rect 20257 6811 20315 6817
rect 16666 6780 16672 6792
rect 14568 6752 15424 6780
rect 15010 6712 15016 6724
rect 14476 6684 15016 6712
rect 15010 6672 15016 6684
rect 15068 6672 15074 6724
rect 15396 6712 15424 6752
rect 15580 6752 16672 6780
rect 15580 6721 15608 6752
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 18141 6783 18199 6789
rect 18141 6749 18153 6783
rect 18187 6780 18199 6783
rect 18325 6783 18383 6789
rect 18325 6780 18337 6783
rect 18187 6752 18337 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 18325 6749 18337 6752
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 15565 6715 15623 6721
rect 15396 6684 15516 6712
rect 12943 6616 13124 6644
rect 12943 6613 12955 6616
rect 12897 6607 12955 6613
rect 13170 6604 13176 6656
rect 13228 6604 13234 6656
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 14826 6644 14832 6656
rect 14415 6616 14832 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 14826 6604 14832 6616
rect 14884 6604 14890 6656
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 15381 6647 15439 6653
rect 15381 6644 15393 6647
rect 15344 6616 15393 6644
rect 15344 6604 15350 6616
rect 15381 6613 15393 6616
rect 15427 6613 15439 6647
rect 15488 6644 15516 6684
rect 15565 6681 15577 6715
rect 15611 6681 15623 6715
rect 15565 6675 15623 6681
rect 15749 6715 15807 6721
rect 15749 6681 15761 6715
rect 15795 6712 15807 6715
rect 15930 6712 15936 6724
rect 15795 6684 15936 6712
rect 15795 6681 15807 6684
rect 15749 6675 15807 6681
rect 15930 6672 15936 6684
rect 15988 6672 15994 6724
rect 16040 6684 16528 6712
rect 16040 6644 16068 6684
rect 15488 6616 16068 6644
rect 16117 6647 16175 6653
rect 15381 6607 15439 6613
rect 16117 6613 16129 6647
rect 16163 6644 16175 6647
rect 16206 6644 16212 6656
rect 16163 6616 16212 6644
rect 16163 6613 16175 6616
rect 16117 6607 16175 6613
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 16500 6644 16528 6684
rect 17954 6672 17960 6724
rect 18012 6712 18018 6724
rect 18984 6712 19012 6811
rect 20622 6808 20628 6820
rect 20680 6808 20686 6860
rect 21542 6808 21548 6860
rect 21600 6848 21606 6860
rect 22664 6857 22692 6888
rect 22922 6876 22928 6888
rect 22980 6876 22986 6928
rect 24228 6888 24440 6916
rect 22649 6851 22707 6857
rect 22649 6848 22661 6851
rect 21600 6820 22661 6848
rect 21600 6808 21606 6820
rect 22649 6817 22661 6820
rect 22695 6817 22707 6851
rect 22649 6811 22707 6817
rect 23842 6808 23848 6860
rect 23900 6808 23906 6860
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6848 23995 6851
rect 24228 6848 24256 6888
rect 23983 6820 24256 6848
rect 24305 6851 24363 6857
rect 23983 6817 23995 6820
rect 23937 6811 23995 6817
rect 24305 6817 24317 6851
rect 24351 6817 24363 6851
rect 24412 6848 24440 6888
rect 24489 6851 24547 6857
rect 24489 6848 24501 6851
rect 24412 6820 24501 6848
rect 24305 6811 24363 6817
rect 24489 6817 24501 6820
rect 24535 6848 24547 6851
rect 26237 6851 26295 6857
rect 24535 6820 25084 6848
rect 24535 6817 24547 6820
rect 24489 6811 24547 6817
rect 19705 6783 19763 6789
rect 19705 6749 19717 6783
rect 19751 6780 19763 6783
rect 19751 6752 19840 6780
rect 19751 6749 19763 6752
rect 19705 6743 19763 6749
rect 19812 6721 19840 6752
rect 20438 6740 20444 6792
rect 20496 6740 20502 6792
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 21177 6783 21235 6789
rect 21177 6780 21189 6783
rect 20772 6752 21189 6780
rect 20772 6740 20778 6752
rect 21177 6749 21189 6752
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 23382 6740 23388 6792
rect 23440 6780 23446 6792
rect 24029 6783 24087 6789
rect 24029 6780 24041 6783
rect 23440 6752 24041 6780
rect 23440 6740 23446 6752
rect 24029 6749 24041 6752
rect 24075 6749 24087 6783
rect 24029 6743 24087 6749
rect 18012 6684 19012 6712
rect 19797 6715 19855 6721
rect 18012 6672 18018 6684
rect 19797 6681 19809 6715
rect 19843 6681 19855 6715
rect 19797 6675 19855 6681
rect 20254 6672 20260 6724
rect 20312 6712 20318 6724
rect 20456 6712 20484 6740
rect 24320 6712 24348 6811
rect 20312 6684 24992 6712
rect 20312 6672 20318 6684
rect 24964 6656 24992 6684
rect 25056 6656 25084 6820
rect 26237 6817 26249 6851
rect 26283 6848 26295 6851
rect 26896 6848 26924 6944
rect 27525 6919 27583 6925
rect 27525 6885 27537 6919
rect 27571 6916 27583 6919
rect 27816 6916 27844 6944
rect 28460 6925 28488 6956
rect 28718 6944 28724 6956
rect 28776 6944 28782 6996
rect 27571 6888 27844 6916
rect 28445 6919 28503 6925
rect 27571 6885 27583 6888
rect 27525 6879 27583 6885
rect 28445 6885 28457 6919
rect 28491 6885 28503 6919
rect 28445 6879 28503 6885
rect 27540 6848 27568 6879
rect 26283 6820 26924 6848
rect 27356 6820 27568 6848
rect 26283 6817 26295 6820
rect 26237 6811 26295 6817
rect 26053 6783 26111 6789
rect 26053 6749 26065 6783
rect 26099 6749 26111 6783
rect 26053 6743 26111 6749
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6780 26479 6783
rect 27065 6783 27123 6789
rect 27065 6780 27077 6783
rect 26467 6752 27077 6780
rect 26467 6749 26479 6752
rect 26421 6743 26479 6749
rect 27065 6749 27077 6752
rect 27111 6749 27123 6783
rect 27065 6743 27123 6749
rect 26068 6712 26096 6743
rect 27356 6712 27384 6820
rect 27614 6808 27620 6860
rect 27672 6848 27678 6860
rect 28169 6851 28227 6857
rect 28169 6848 28181 6851
rect 27672 6820 28181 6848
rect 27672 6808 27678 6820
rect 28169 6817 28181 6820
rect 28215 6817 28227 6851
rect 28169 6811 28227 6817
rect 28258 6808 28264 6860
rect 28316 6848 28322 6860
rect 29917 6851 29975 6857
rect 29917 6848 29929 6851
rect 28316 6820 29929 6848
rect 28316 6808 28322 6820
rect 29917 6817 29929 6820
rect 29963 6817 29975 6851
rect 31481 6851 31539 6857
rect 31481 6848 31493 6851
rect 29917 6811 29975 6817
rect 30300 6820 31493 6848
rect 27433 6783 27491 6789
rect 27433 6749 27445 6783
rect 27479 6780 27491 6783
rect 27890 6780 27896 6792
rect 27479 6752 27896 6780
rect 27479 6749 27491 6752
rect 27433 6743 27491 6749
rect 27890 6740 27896 6752
rect 27948 6780 27954 6792
rect 28629 6783 28687 6789
rect 28629 6780 28641 6783
rect 27948 6752 28212 6780
rect 27948 6740 27954 6752
rect 26068 6684 27384 6712
rect 17678 6644 17684 6656
rect 16500 6616 17684 6644
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 19058 6604 19064 6656
rect 19116 6604 19122 6656
rect 24670 6604 24676 6656
rect 24728 6604 24734 6656
rect 24946 6604 24952 6656
rect 25004 6604 25010 6656
rect 25038 6604 25044 6656
rect 25096 6604 25102 6656
rect 28184 6644 28212 6752
rect 28460 6752 28641 6780
rect 28460 6721 28488 6752
rect 28629 6749 28641 6752
rect 28675 6749 28687 6783
rect 28629 6743 28687 6749
rect 28718 6740 28724 6792
rect 28776 6780 28782 6792
rect 28776 6752 29500 6780
rect 28776 6740 28782 6752
rect 28445 6715 28503 6721
rect 28445 6681 28457 6715
rect 28491 6681 28503 6715
rect 29365 6715 29423 6721
rect 29365 6712 29377 6715
rect 28445 6675 28503 6681
rect 28552 6684 29377 6712
rect 28552 6644 28580 6684
rect 29365 6681 29377 6684
rect 29411 6681 29423 6715
rect 29472 6712 29500 6752
rect 29822 6740 29828 6792
rect 29880 6780 29886 6792
rect 30300 6780 30328 6820
rect 31481 6817 31493 6820
rect 31527 6817 31539 6851
rect 31481 6811 31539 6817
rect 29880 6752 30328 6780
rect 29880 6740 29886 6752
rect 30650 6740 30656 6792
rect 30708 6740 30714 6792
rect 31297 6715 31355 6721
rect 31297 6712 31309 6715
rect 29472 6684 31309 6712
rect 29365 6675 29423 6681
rect 31297 6681 31309 6684
rect 31343 6681 31355 6715
rect 31297 6675 31355 6681
rect 28184 6616 28580 6644
rect 28810 6604 28816 6656
rect 28868 6644 28874 6656
rect 29273 6647 29331 6653
rect 29273 6644 29285 6647
rect 28868 6616 29285 6644
rect 28868 6604 28874 6616
rect 29273 6613 29285 6616
rect 29319 6613 29331 6647
rect 29273 6607 29331 6613
rect 30098 6604 30104 6656
rect 30156 6604 30162 6656
rect 2760 6554 32200 6576
rect 2760 6502 6286 6554
rect 6338 6502 6350 6554
rect 6402 6502 6414 6554
rect 6466 6502 6478 6554
rect 6530 6502 6542 6554
rect 6594 6502 13646 6554
rect 13698 6502 13710 6554
rect 13762 6502 13774 6554
rect 13826 6502 13838 6554
rect 13890 6502 13902 6554
rect 13954 6502 21006 6554
rect 21058 6502 21070 6554
rect 21122 6502 21134 6554
rect 21186 6502 21198 6554
rect 21250 6502 21262 6554
rect 21314 6502 28366 6554
rect 28418 6502 28430 6554
rect 28482 6502 28494 6554
rect 28546 6502 28558 6554
rect 28610 6502 28622 6554
rect 28674 6502 32200 6554
rect 2760 6480 32200 6502
rect 6914 6400 6920 6452
rect 6972 6400 6978 6452
rect 13170 6400 13176 6452
rect 13228 6400 13234 6452
rect 15010 6400 15016 6452
rect 15068 6440 15074 6452
rect 15930 6440 15936 6452
rect 15068 6412 15936 6440
rect 15068 6400 15074 6412
rect 15930 6400 15936 6412
rect 15988 6400 15994 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6440 17279 6443
rect 17310 6440 17316 6452
rect 17267 6412 17316 6440
rect 17267 6409 17279 6412
rect 17221 6403 17279 6409
rect 17310 6400 17316 6412
rect 17368 6400 17374 6452
rect 18414 6400 18420 6452
rect 18472 6400 18478 6452
rect 19058 6400 19064 6452
rect 19116 6400 19122 6452
rect 20714 6400 20720 6452
rect 20772 6400 20778 6452
rect 24670 6400 24676 6452
rect 24728 6400 24734 6452
rect 28258 6400 28264 6452
rect 28316 6440 28322 6452
rect 28445 6443 28503 6449
rect 28445 6440 28457 6443
rect 28316 6412 28457 6440
rect 28316 6400 28322 6412
rect 28445 6409 28457 6412
rect 28491 6409 28503 6443
rect 28445 6403 28503 6409
rect 28800 6443 28858 6449
rect 28800 6409 28812 6443
rect 28846 6440 28858 6443
rect 30098 6440 30104 6452
rect 28846 6412 30104 6440
rect 28846 6409 28858 6412
rect 28800 6403 28858 6409
rect 30098 6400 30104 6412
rect 30156 6400 30162 6452
rect 30466 6400 30472 6452
rect 30524 6400 30530 6452
rect 6932 6304 6960 6400
rect 7193 6307 7251 6313
rect 7193 6304 7205 6307
rect 6932 6276 7205 6304
rect 7193 6273 7205 6276
rect 7239 6273 7251 6307
rect 13188 6304 13216 6400
rect 13262 6332 13268 6384
rect 13320 6372 13326 6384
rect 16850 6372 16856 6384
rect 13320 6344 16856 6372
rect 13320 6332 13326 6344
rect 16850 6332 16856 6344
rect 16908 6372 16914 6384
rect 17678 6372 17684 6384
rect 16908 6344 17684 6372
rect 16908 6332 16914 6344
rect 17678 6332 17684 6344
rect 17736 6332 17742 6384
rect 18230 6332 18236 6384
rect 18288 6372 18294 6384
rect 18288 6344 18552 6372
rect 18288 6332 18294 6344
rect 13449 6307 13507 6313
rect 13449 6304 13461 6307
rect 7193 6267 7251 6273
rect 7300 6276 12434 6304
rect 13188 6276 13461 6304
rect 1302 6196 1308 6248
rect 1360 6236 1366 6248
rect 3053 6239 3111 6245
rect 3053 6236 3065 6239
rect 1360 6208 3065 6236
rect 1360 6196 1366 6208
rect 3053 6205 3065 6208
rect 3099 6205 3111 6239
rect 3053 6199 3111 6205
rect 5350 6196 5356 6248
rect 5408 6236 5414 6248
rect 7300 6236 7328 6276
rect 5408 6208 7328 6236
rect 5408 6196 5414 6208
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8113 6239 8171 6245
rect 8113 6236 8125 6239
rect 7892 6208 8125 6236
rect 7892 6196 7898 6208
rect 8113 6205 8125 6208
rect 8159 6205 8171 6239
rect 8113 6199 8171 6205
rect 9766 6196 9772 6248
rect 9824 6196 9830 6248
rect 11606 6196 11612 6248
rect 11664 6196 11670 6248
rect 11624 6168 11652 6196
rect 3252 6140 11652 6168
rect 3252 6109 3280 6140
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6069 3295 6103
rect 3237 6063 3295 6069
rect 6638 6060 6644 6112
rect 6696 6060 6702 6112
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7558 6100 7564 6112
rect 7248 6072 7564 6100
rect 7248 6060 7254 6072
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 9030 6060 9036 6112
rect 9088 6100 9094 6112
rect 9217 6103 9275 6109
rect 9217 6100 9229 6103
rect 9088 6072 9229 6100
rect 9088 6060 9094 6072
rect 9217 6069 9229 6072
rect 9263 6069 9275 6103
rect 12406 6100 12434 6276
rect 13449 6273 13461 6276
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 17911 6276 18368 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 14182 6196 14188 6248
rect 14240 6236 14246 6248
rect 14369 6239 14427 6245
rect 14369 6236 14381 6239
rect 14240 6208 14381 6236
rect 14240 6196 14246 6208
rect 14369 6205 14381 6208
rect 14415 6205 14427 6239
rect 14369 6199 14427 6205
rect 15197 6239 15255 6245
rect 15197 6205 15209 6239
rect 15243 6236 15255 6239
rect 15286 6236 15292 6248
rect 15243 6208 15292 6236
rect 15243 6205 15255 6208
rect 15197 6199 15255 6205
rect 15286 6196 15292 6208
rect 15344 6196 15350 6248
rect 16390 6196 16396 6248
rect 16448 6196 16454 6248
rect 17129 6239 17187 6245
rect 17129 6205 17141 6239
rect 17175 6236 17187 6239
rect 17310 6236 17316 6248
rect 17175 6208 17316 6236
rect 17175 6205 17187 6208
rect 17129 6199 17187 6205
rect 17310 6196 17316 6208
rect 17368 6196 17374 6248
rect 17589 6239 17647 6245
rect 17589 6205 17601 6239
rect 17635 6236 17647 6239
rect 17954 6236 17960 6248
rect 17635 6208 17960 6236
rect 17635 6205 17647 6208
rect 17589 6199 17647 6205
rect 17954 6196 17960 6208
rect 18012 6196 18018 6248
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 14274 6168 14280 6180
rect 13964 6140 14280 6168
rect 13964 6128 13970 6140
rect 14274 6128 14280 6140
rect 14332 6168 14338 6180
rect 15565 6171 15623 6177
rect 15565 6168 15577 6171
rect 14332 6140 15577 6168
rect 14332 6128 14338 6140
rect 15565 6137 15577 6140
rect 15611 6168 15623 6171
rect 16485 6171 16543 6177
rect 15611 6140 15884 6168
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 12802 6100 12808 6112
rect 12406 6072 12808 6100
rect 9217 6063 9275 6069
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 12894 6060 12900 6112
rect 12952 6060 12958 6112
rect 13538 6060 13544 6112
rect 13596 6100 13602 6112
rect 13817 6103 13875 6109
rect 13817 6100 13829 6103
rect 13596 6072 13829 6100
rect 13596 6060 13602 6072
rect 13817 6069 13829 6072
rect 13863 6069 13875 6103
rect 13817 6063 13875 6069
rect 14553 6103 14611 6109
rect 14553 6069 14565 6103
rect 14599 6100 14611 6103
rect 14642 6100 14648 6112
rect 14599 6072 14648 6100
rect 14599 6069 14611 6072
rect 14553 6063 14611 6069
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 15746 6060 15752 6112
rect 15804 6060 15810 6112
rect 15856 6100 15884 6140
rect 16485 6137 16497 6171
rect 16531 6168 16543 6171
rect 16850 6168 16856 6180
rect 16531 6140 16856 6168
rect 16531 6137 16543 6140
rect 16485 6131 16543 6137
rect 16850 6128 16856 6140
rect 16908 6168 16914 6180
rect 17681 6171 17739 6177
rect 17681 6168 17693 6171
rect 16908 6140 17693 6168
rect 16908 6128 16914 6140
rect 17681 6137 17693 6140
rect 17727 6137 17739 6171
rect 17681 6131 17739 6137
rect 16574 6100 16580 6112
rect 15856 6072 16580 6100
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 18340 6100 18368 6276
rect 18524 6245 18552 6344
rect 19076 6304 19104 6400
rect 19245 6307 19303 6313
rect 19245 6304 19257 6307
rect 19076 6276 19257 6304
rect 19245 6273 19257 6276
rect 19291 6273 19303 6307
rect 21542 6304 21548 6316
rect 19245 6267 19303 6273
rect 21100 6276 21548 6304
rect 18509 6239 18567 6245
rect 18509 6205 18521 6239
rect 18555 6205 18567 6239
rect 18509 6199 18567 6205
rect 18782 6196 18788 6248
rect 18840 6236 18846 6248
rect 21100 6245 21128 6276
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 22094 6264 22100 6316
rect 22152 6304 22158 6316
rect 22189 6307 22247 6313
rect 22189 6304 22201 6307
rect 22152 6276 22201 6304
rect 22152 6264 22158 6276
rect 22189 6273 22201 6276
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 22465 6307 22523 6313
rect 22465 6273 22477 6307
rect 22511 6304 22523 6307
rect 24029 6307 24087 6313
rect 24029 6304 24041 6307
rect 22511 6276 24041 6304
rect 22511 6273 22523 6276
rect 22465 6267 22523 6273
rect 24029 6273 24041 6276
rect 24075 6273 24087 6307
rect 24688 6304 24716 6400
rect 29822 6332 29828 6384
rect 29880 6372 29886 6384
rect 30285 6375 30343 6381
rect 30285 6372 30297 6375
rect 29880 6344 30297 6372
rect 29880 6332 29886 6344
rect 30285 6341 30297 6344
rect 30331 6341 30343 6375
rect 30285 6335 30343 6341
rect 31665 6375 31723 6381
rect 31665 6341 31677 6375
rect 31711 6341 31723 6375
rect 31665 6335 31723 6341
rect 25317 6307 25375 6313
rect 25317 6304 25329 6307
rect 24688 6276 25329 6304
rect 24029 6267 24087 6273
rect 25317 6273 25329 6276
rect 25363 6273 25375 6307
rect 25317 6267 25375 6273
rect 26234 6264 26240 6316
rect 26292 6304 26298 6316
rect 26697 6307 26755 6313
rect 26697 6304 26709 6307
rect 26292 6276 26709 6304
rect 26292 6264 26298 6276
rect 26697 6273 26709 6276
rect 26743 6304 26755 6307
rect 27614 6304 27620 6316
rect 26743 6276 27620 6304
rect 26743 6273 26755 6276
rect 26697 6267 26755 6273
rect 27614 6264 27620 6276
rect 27672 6304 27678 6316
rect 28537 6307 28595 6313
rect 28537 6304 28549 6307
rect 27672 6276 28549 6304
rect 27672 6264 27678 6276
rect 28537 6273 28549 6276
rect 28583 6304 28595 6307
rect 28902 6304 28908 6316
rect 28583 6276 28908 6304
rect 28583 6273 28595 6276
rect 28537 6267 28595 6273
rect 28902 6264 28908 6276
rect 28960 6264 28966 6316
rect 30006 6264 30012 6316
rect 30064 6304 30070 6316
rect 31680 6304 31708 6335
rect 30064 6276 31708 6304
rect 30064 6264 30070 6276
rect 18969 6239 19027 6245
rect 18969 6236 18981 6239
rect 18840 6208 18981 6236
rect 18840 6196 18846 6208
rect 18969 6205 18981 6208
rect 19015 6205 19027 6239
rect 18969 6199 19027 6205
rect 21085 6239 21143 6245
rect 21085 6205 21097 6239
rect 21131 6205 21143 6239
rect 21085 6199 21143 6205
rect 23566 6196 23572 6248
rect 23624 6196 23630 6248
rect 24578 6196 24584 6248
rect 24636 6196 24642 6248
rect 30561 6239 30619 6245
rect 30561 6205 30573 6239
rect 30607 6236 30619 6239
rect 31202 6236 31208 6248
rect 30607 6208 31208 6236
rect 30607 6205 30619 6208
rect 30561 6199 30619 6205
rect 20993 6171 21051 6177
rect 20993 6168 21005 6171
rect 20470 6140 21005 6168
rect 20993 6137 21005 6140
rect 21039 6137 21051 6171
rect 20993 6131 21051 6137
rect 26973 6171 27031 6177
rect 26973 6137 26985 6171
rect 27019 6168 27031 6171
rect 27246 6168 27252 6180
rect 27019 6140 27252 6168
rect 27019 6137 27031 6140
rect 26973 6131 27031 6137
rect 27246 6128 27252 6140
rect 27304 6128 27310 6180
rect 27706 6128 27712 6180
rect 27764 6128 27770 6180
rect 29546 6128 29552 6180
rect 29604 6128 29610 6180
rect 18877 6103 18935 6109
rect 18877 6100 18889 6103
rect 18340 6072 18889 6100
rect 18877 6069 18889 6072
rect 18923 6100 18935 6103
rect 20254 6100 20260 6112
rect 18923 6072 20260 6100
rect 18923 6069 18935 6072
rect 18877 6063 18935 6069
rect 20254 6060 20260 6072
rect 20312 6060 20318 6112
rect 23934 6060 23940 6112
rect 23992 6060 23998 6112
rect 24026 6060 24032 6112
rect 24084 6100 24090 6112
rect 24765 6103 24823 6109
rect 24765 6100 24777 6103
rect 24084 6072 24777 6100
rect 24084 6060 24090 6072
rect 24765 6069 24777 6072
rect 24811 6069 24823 6103
rect 24765 6063 24823 6069
rect 29454 6060 29460 6112
rect 29512 6100 29518 6112
rect 30576 6100 30604 6199
rect 31202 6196 31208 6208
rect 31260 6196 31266 6248
rect 31849 6239 31907 6245
rect 31849 6205 31861 6239
rect 31895 6236 31907 6239
rect 33134 6236 33140 6248
rect 31895 6208 33140 6236
rect 31895 6205 31907 6208
rect 31849 6199 31907 6205
rect 33134 6196 33140 6208
rect 33192 6196 33198 6248
rect 29512 6072 30604 6100
rect 29512 6060 29518 6072
rect 2760 6010 32200 6032
rect 2760 5958 6946 6010
rect 6998 5958 7010 6010
rect 7062 5958 7074 6010
rect 7126 5958 7138 6010
rect 7190 5958 7202 6010
rect 7254 5958 14306 6010
rect 14358 5958 14370 6010
rect 14422 5958 14434 6010
rect 14486 5958 14498 6010
rect 14550 5958 14562 6010
rect 14614 5958 21666 6010
rect 21718 5958 21730 6010
rect 21782 5958 21794 6010
rect 21846 5958 21858 6010
rect 21910 5958 21922 6010
rect 21974 5958 29026 6010
rect 29078 5958 29090 6010
rect 29142 5958 29154 6010
rect 29206 5958 29218 6010
rect 29270 5958 29282 6010
rect 29334 5958 32200 6010
rect 2760 5936 32200 5958
rect 6638 5856 6644 5908
rect 6696 5856 6702 5908
rect 7834 5856 7840 5908
rect 7892 5856 7898 5908
rect 9401 5899 9459 5905
rect 9401 5865 9413 5899
rect 9447 5896 9459 5899
rect 9766 5896 9772 5908
rect 9447 5868 9772 5896
rect 9447 5865 9459 5868
rect 9401 5859 9459 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 9861 5899 9919 5905
rect 9861 5865 9873 5899
rect 9907 5896 9919 5899
rect 9950 5896 9956 5908
rect 9907 5868 9956 5896
rect 9907 5865 9919 5868
rect 9861 5859 9919 5865
rect 9950 5856 9956 5868
rect 10008 5856 10014 5908
rect 12986 5856 12992 5908
rect 13044 5856 13050 5908
rect 14826 5896 14832 5908
rect 13832 5868 14832 5896
rect 6365 5831 6423 5837
rect 6365 5797 6377 5831
rect 6411 5828 6423 5831
rect 6656 5828 6684 5856
rect 8113 5831 8171 5837
rect 8113 5828 8125 5831
rect 6411 5800 6684 5828
rect 7590 5800 8125 5828
rect 6411 5797 6423 5800
rect 6365 5791 6423 5797
rect 8113 5797 8125 5800
rect 8159 5797 8171 5831
rect 8113 5791 8171 5797
rect 12621 5831 12679 5837
rect 12621 5797 12633 5831
rect 12667 5828 12679 5831
rect 13832 5828 13860 5868
rect 14826 5856 14832 5868
rect 14884 5856 14890 5908
rect 15378 5856 15384 5908
rect 15436 5896 15442 5908
rect 15473 5899 15531 5905
rect 15473 5896 15485 5899
rect 15436 5868 15485 5896
rect 15436 5856 15442 5868
rect 15473 5865 15485 5868
rect 15519 5865 15531 5899
rect 15473 5859 15531 5865
rect 15746 5856 15752 5908
rect 15804 5896 15810 5908
rect 15804 5868 15884 5896
rect 15804 5856 15810 5868
rect 15856 5837 15884 5868
rect 17310 5856 17316 5908
rect 17368 5856 17374 5908
rect 17678 5856 17684 5908
rect 17736 5856 17742 5908
rect 18598 5856 18604 5908
rect 18656 5896 18662 5908
rect 19058 5896 19064 5908
rect 18656 5868 19064 5896
rect 18656 5856 18662 5868
rect 19058 5856 19064 5868
rect 19116 5856 19122 5908
rect 20622 5856 20628 5908
rect 20680 5856 20686 5908
rect 21542 5856 21548 5908
rect 21600 5856 21606 5908
rect 22373 5899 22431 5905
rect 22373 5865 22385 5899
rect 22419 5896 22431 5899
rect 23750 5896 23756 5908
rect 22419 5868 23756 5896
rect 22419 5865 22431 5868
rect 22373 5859 22431 5865
rect 23750 5856 23756 5868
rect 23808 5856 23814 5908
rect 23842 5856 23848 5908
rect 23900 5856 23906 5908
rect 23934 5856 23940 5908
rect 23992 5856 23998 5908
rect 24213 5899 24271 5905
rect 24213 5865 24225 5899
rect 24259 5896 24271 5899
rect 24578 5896 24584 5908
rect 24259 5868 24584 5896
rect 24259 5865 24271 5868
rect 24213 5859 24271 5865
rect 24578 5856 24584 5868
rect 24636 5856 24642 5908
rect 25038 5856 25044 5908
rect 25096 5856 25102 5908
rect 27706 5856 27712 5908
rect 27764 5896 27770 5908
rect 27801 5899 27859 5905
rect 27801 5896 27813 5899
rect 27764 5868 27813 5896
rect 27764 5856 27770 5868
rect 27801 5865 27813 5868
rect 27847 5865 27859 5899
rect 27801 5859 27859 5865
rect 28810 5856 28816 5908
rect 28868 5856 28874 5908
rect 28905 5899 28963 5905
rect 28905 5865 28917 5899
rect 28951 5865 28963 5899
rect 28905 5859 28963 5865
rect 12667 5800 13860 5828
rect 15841 5831 15899 5837
rect 12667 5797 12679 5800
rect 12621 5791 12679 5797
rect 15841 5797 15853 5831
rect 15887 5797 15899 5831
rect 17126 5828 17132 5840
rect 17066 5800 17132 5828
rect 15841 5791 15899 5797
rect 17126 5788 17132 5800
rect 17184 5788 17190 5840
rect 17696 5828 17724 5856
rect 18690 5828 18696 5840
rect 17696 5800 18696 5828
rect 18690 5788 18696 5800
rect 18748 5788 18754 5840
rect 21453 5831 21511 5837
rect 21453 5828 21465 5831
rect 20286 5800 21465 5828
rect 21453 5797 21465 5800
rect 21499 5797 21511 5831
rect 21453 5791 21511 5797
rect 8202 5720 8208 5772
rect 8260 5720 8266 5772
rect 9769 5763 9827 5769
rect 9769 5729 9781 5763
rect 9815 5760 9827 5763
rect 10410 5760 10416 5772
rect 9815 5732 10416 5760
rect 9815 5729 9827 5732
rect 9769 5723 9827 5729
rect 10410 5720 10416 5732
rect 10468 5720 10474 5772
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 13817 5763 13875 5769
rect 13817 5760 13829 5763
rect 12860 5732 13829 5760
rect 12860 5720 12866 5732
rect 13817 5729 13829 5732
rect 13863 5729 13875 5763
rect 13817 5723 13875 5729
rect 14826 5720 14832 5772
rect 14884 5720 14890 5772
rect 21560 5769 21588 5856
rect 22554 5828 22560 5840
rect 22204 5800 22560 5828
rect 22204 5769 22232 5800
rect 22554 5788 22560 5800
rect 22612 5788 22618 5840
rect 22738 5788 22744 5840
rect 22796 5788 22802 5840
rect 21545 5763 21603 5769
rect 21545 5729 21557 5763
rect 21591 5729 21603 5763
rect 21545 5723 21603 5729
rect 22189 5763 22247 5769
rect 22189 5729 22201 5763
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 22465 5763 22523 5769
rect 22465 5729 22477 5763
rect 22511 5760 22523 5763
rect 23109 5763 23167 5769
rect 23109 5760 23121 5763
rect 22511 5732 23121 5760
rect 22511 5729 22523 5732
rect 22465 5723 22523 5729
rect 23109 5729 23121 5732
rect 23155 5729 23167 5763
rect 23109 5723 23167 5729
rect 5350 5652 5356 5704
rect 5408 5652 5414 5704
rect 6086 5652 6092 5704
rect 6144 5652 6150 5704
rect 9582 5692 9588 5704
rect 9232 5664 9588 5692
rect 5994 5516 6000 5568
rect 6052 5516 6058 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 9232 5565 9260 5664
rect 9582 5652 9588 5664
rect 9640 5692 9646 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9640 5664 9965 5692
rect 9640 5652 9646 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13633 5695 13691 5701
rect 13633 5692 13645 5695
rect 13044 5664 13645 5692
rect 13044 5652 13050 5664
rect 13633 5661 13645 5664
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13964 5664 14289 5692
rect 13964 5652 13970 5664
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14277 5655 14335 5661
rect 14384 5664 14565 5692
rect 13541 5627 13599 5633
rect 13541 5593 13553 5627
rect 13587 5624 13599 5627
rect 13924 5624 13952 5652
rect 13587 5596 13952 5624
rect 13587 5593 13599 5596
rect 13541 5587 13599 5593
rect 9217 5559 9275 5565
rect 9217 5556 9229 5559
rect 8352 5528 9229 5556
rect 8352 5516 8358 5528
rect 9217 5525 9229 5528
rect 9263 5525 9275 5559
rect 14384 5556 14412 5664
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 14691 5695 14749 5701
rect 14691 5661 14703 5695
rect 14737 5692 14749 5695
rect 15010 5692 15016 5704
rect 14737 5664 15016 5692
rect 14737 5661 14749 5664
rect 14691 5655 14749 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15565 5695 15623 5701
rect 15565 5692 15577 5695
rect 15252 5664 15577 5692
rect 15252 5652 15258 5664
rect 15565 5661 15577 5664
rect 15611 5661 15623 5695
rect 15565 5655 15623 5661
rect 18782 5652 18788 5704
rect 18840 5652 18846 5704
rect 19061 5695 19119 5701
rect 19061 5661 19073 5695
rect 19107 5692 19119 5695
rect 19518 5692 19524 5704
rect 19107 5664 19524 5692
rect 19107 5661 19119 5664
rect 19061 5655 19119 5661
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5692 20591 5695
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 20579 5664 21189 5692
rect 20579 5661 20591 5664
rect 20533 5655 20591 5661
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 21634 5652 21640 5704
rect 21692 5692 21698 5704
rect 22480 5692 22508 5723
rect 21692 5664 22508 5692
rect 23661 5695 23719 5701
rect 21692 5652 21698 5664
rect 23661 5661 23673 5695
rect 23707 5661 23719 5695
rect 23860 5692 23888 5856
rect 23952 5760 23980 5856
rect 24946 5788 24952 5840
rect 25004 5828 25010 5840
rect 26053 5831 26111 5837
rect 26053 5828 26065 5831
rect 25004 5800 26065 5828
rect 25004 5788 25010 5800
rect 26053 5797 26065 5800
rect 26099 5828 26111 5831
rect 28629 5831 28687 5837
rect 28629 5828 28641 5831
rect 26099 5800 28641 5828
rect 26099 5797 26111 5800
rect 26053 5791 26111 5797
rect 28629 5797 28641 5800
rect 28675 5828 28687 5831
rect 28675 5800 28764 5828
rect 28675 5797 28687 5800
rect 28629 5791 28687 5797
rect 24857 5763 24915 5769
rect 24857 5760 24869 5763
rect 23952 5732 24869 5760
rect 24857 5729 24869 5732
rect 24903 5729 24915 5763
rect 24857 5723 24915 5729
rect 24305 5695 24363 5701
rect 24305 5692 24317 5695
rect 23860 5664 24317 5692
rect 23661 5655 23719 5661
rect 24305 5661 24317 5664
rect 24351 5661 24363 5695
rect 24305 5655 24363 5661
rect 15470 5584 15476 5636
rect 15528 5584 15534 5636
rect 21358 5584 21364 5636
rect 21416 5624 21422 5636
rect 23676 5624 23704 5655
rect 24964 5624 24992 5788
rect 28736 5772 28764 5800
rect 27709 5763 27767 5769
rect 27709 5729 27721 5763
rect 27755 5760 27767 5763
rect 28166 5760 28172 5772
rect 27755 5732 28172 5760
rect 27755 5729 27767 5732
rect 27709 5723 27767 5729
rect 28166 5720 28172 5732
rect 28224 5720 28230 5772
rect 28718 5720 28724 5772
rect 28776 5720 28782 5772
rect 28828 5760 28856 5856
rect 28920 5828 28948 5859
rect 29546 5856 29552 5908
rect 29604 5856 29610 5908
rect 30650 5856 30656 5908
rect 30708 5856 30714 5908
rect 30668 5828 30696 5856
rect 28920 5800 30696 5828
rect 28905 5763 28963 5769
rect 28905 5760 28917 5763
rect 28828 5732 28917 5760
rect 28905 5729 28917 5732
rect 28951 5729 28963 5763
rect 28905 5723 28963 5729
rect 29454 5720 29460 5772
rect 29512 5720 29518 5772
rect 25590 5652 25596 5704
rect 25648 5652 25654 5704
rect 21416 5596 22784 5624
rect 23676 5596 24992 5624
rect 28184 5624 28212 5720
rect 28813 5695 28871 5701
rect 28813 5661 28825 5695
rect 28859 5692 28871 5695
rect 29362 5692 29368 5704
rect 28859 5664 29368 5692
rect 28859 5661 28871 5664
rect 28813 5655 28871 5661
rect 29362 5652 29368 5664
rect 29420 5652 29426 5704
rect 29472 5624 29500 5720
rect 28184 5596 29500 5624
rect 21416 5584 21422 5596
rect 14826 5556 14832 5568
rect 14384 5528 14832 5556
rect 9217 5519 9275 5525
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 15488 5556 15516 5584
rect 16022 5556 16028 5568
rect 15488 5528 16028 5556
rect 16022 5516 16028 5528
rect 16080 5556 16086 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 16080 5528 18061 5556
rect 16080 5516 16086 5528
rect 18049 5525 18061 5528
rect 18095 5556 18107 5559
rect 18414 5556 18420 5568
rect 18095 5528 18420 5556
rect 18095 5525 18107 5528
rect 18049 5519 18107 5525
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 22005 5559 22063 5565
rect 22005 5525 22017 5559
rect 22051 5556 22063 5559
rect 22370 5556 22376 5568
rect 22051 5528 22376 5556
rect 22051 5525 22063 5528
rect 22005 5519 22063 5525
rect 22370 5516 22376 5528
rect 22428 5516 22434 5568
rect 22554 5516 22560 5568
rect 22612 5516 22618 5568
rect 22756 5565 22784 5596
rect 22741 5559 22799 5565
rect 22741 5525 22753 5559
rect 22787 5525 22799 5559
rect 22741 5519 22799 5525
rect 23658 5516 23664 5568
rect 23716 5556 23722 5568
rect 24486 5556 24492 5568
rect 23716 5528 24492 5556
rect 23716 5516 23722 5528
rect 24486 5516 24492 5528
rect 24544 5516 24550 5568
rect 28718 5516 28724 5568
rect 28776 5556 28782 5568
rect 29273 5559 29331 5565
rect 29273 5556 29285 5559
rect 28776 5528 29285 5556
rect 28776 5516 28782 5528
rect 29273 5525 29285 5528
rect 29319 5556 29331 5559
rect 29914 5556 29920 5568
rect 29319 5528 29920 5556
rect 29319 5525 29331 5528
rect 29273 5519 29331 5525
rect 29914 5516 29920 5528
rect 29972 5516 29978 5568
rect 2760 5466 32200 5488
rect 2760 5414 6286 5466
rect 6338 5414 6350 5466
rect 6402 5414 6414 5466
rect 6466 5414 6478 5466
rect 6530 5414 6542 5466
rect 6594 5414 13646 5466
rect 13698 5414 13710 5466
rect 13762 5414 13774 5466
rect 13826 5414 13838 5466
rect 13890 5414 13902 5466
rect 13954 5414 21006 5466
rect 21058 5414 21070 5466
rect 21122 5414 21134 5466
rect 21186 5414 21198 5466
rect 21250 5414 21262 5466
rect 21314 5414 28366 5466
rect 28418 5414 28430 5466
rect 28482 5414 28494 5466
rect 28546 5414 28558 5466
rect 28610 5414 28622 5466
rect 28674 5414 32200 5466
rect 2760 5392 32200 5414
rect 6730 5352 6736 5364
rect 5828 5324 6736 5352
rect 5828 5225 5856 5324
rect 6730 5312 6736 5324
rect 6788 5352 6794 5364
rect 6917 5355 6975 5361
rect 6917 5352 6929 5355
rect 6788 5324 6929 5352
rect 6788 5312 6794 5324
rect 6917 5321 6929 5324
rect 6963 5352 6975 5355
rect 8294 5352 8300 5364
rect 6963 5324 8300 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 8294 5312 8300 5324
rect 8352 5312 8358 5364
rect 12986 5312 12992 5364
rect 13044 5352 13050 5364
rect 13044 5324 14136 5352
rect 13044 5312 13050 5324
rect 7558 5284 7564 5296
rect 5920 5256 7564 5284
rect 5920 5225 5948 5256
rect 7558 5244 7564 5256
rect 7616 5244 7622 5296
rect 5813 5219 5871 5225
rect 5813 5185 5825 5219
rect 5859 5185 5871 5219
rect 5813 5179 5871 5185
rect 5905 5219 5963 5225
rect 5905 5185 5917 5219
rect 5951 5185 5963 5219
rect 5905 5179 5963 5185
rect 6086 5176 6092 5228
rect 6144 5216 6150 5228
rect 8665 5219 8723 5225
rect 8665 5216 8677 5219
rect 6144 5188 8677 5216
rect 6144 5176 6150 5188
rect 8665 5185 8677 5188
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8941 5219 8999 5225
rect 8941 5185 8953 5219
rect 8987 5216 8999 5219
rect 9030 5216 9036 5228
rect 8987 5188 9036 5216
rect 8987 5185 8999 5188
rect 8941 5179 8999 5185
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 9582 5176 9588 5228
rect 9640 5216 9646 5228
rect 12250 5216 12256 5228
rect 9640 5188 12256 5216
rect 9640 5176 9646 5188
rect 12250 5176 12256 5188
rect 12308 5216 12314 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 12308 5188 12357 5216
rect 12308 5176 12314 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12526 5176 12532 5228
rect 12584 5176 12590 5228
rect 12805 5219 12863 5225
rect 12805 5185 12817 5219
rect 12851 5216 12863 5219
rect 12894 5216 12900 5228
rect 12851 5188 12900 5216
rect 12851 5185 12863 5188
rect 12805 5179 12863 5185
rect 12894 5176 12900 5188
rect 12952 5176 12958 5228
rect 14108 5216 14136 5324
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 14240 5324 14289 5352
rect 14240 5312 14246 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 16390 5312 16396 5364
rect 16448 5352 16454 5364
rect 16485 5355 16543 5361
rect 16485 5352 16497 5355
rect 16448 5324 16497 5352
rect 16448 5312 16454 5324
rect 16485 5321 16497 5324
rect 16531 5321 16543 5355
rect 16485 5315 16543 5321
rect 17126 5312 17132 5364
rect 17184 5312 17190 5364
rect 17954 5352 17960 5364
rect 17696 5324 17960 5352
rect 17696 5284 17724 5324
rect 17954 5312 17960 5324
rect 18012 5312 18018 5364
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 18104 5324 19334 5352
rect 18104 5312 18110 5324
rect 19306 5284 19334 5324
rect 19518 5312 19524 5364
rect 19576 5312 19582 5364
rect 21085 5355 21143 5361
rect 20180 5324 21036 5352
rect 20070 5284 20076 5296
rect 14844 5256 17724 5284
rect 18616 5256 19012 5284
rect 19306 5256 20076 5284
rect 14844 5225 14872 5256
rect 14829 5219 14887 5225
rect 14829 5216 14841 5219
rect 14108 5188 14841 5216
rect 14829 5185 14841 5188
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 15013 5219 15071 5225
rect 15013 5185 15025 5219
rect 15059 5216 15071 5219
rect 15194 5216 15200 5228
rect 15059 5188 15200 5216
rect 15059 5185 15071 5188
rect 15013 5179 15071 5185
rect 15194 5176 15200 5188
rect 15252 5176 15258 5228
rect 15565 5219 15623 5225
rect 15565 5185 15577 5219
rect 15611 5216 15623 5219
rect 15746 5216 15752 5228
rect 15611 5188 15752 5216
rect 15611 5185 15623 5188
rect 15565 5179 15623 5185
rect 4338 5108 4344 5160
rect 4396 5108 4402 5160
rect 5994 5108 6000 5160
rect 6052 5108 6058 5160
rect 6457 5151 6515 5157
rect 6457 5117 6469 5151
rect 6503 5148 6515 5151
rect 6914 5148 6920 5160
rect 6503 5120 6920 5148
rect 6503 5117 6515 5120
rect 6457 5111 6515 5117
rect 6914 5108 6920 5120
rect 6972 5148 6978 5160
rect 6972 5120 7604 5148
rect 6972 5108 6978 5120
rect 1302 5040 1308 5092
rect 1360 5080 1366 5092
rect 3237 5083 3295 5089
rect 3237 5080 3249 5083
rect 1360 5052 3249 5080
rect 1360 5040 1366 5052
rect 3237 5049 3249 5052
rect 3283 5049 3295 5083
rect 3237 5043 3295 5049
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 7101 5083 7159 5089
rect 7101 5080 7113 5083
rect 6880 5052 7113 5080
rect 6880 5040 6886 5052
rect 7101 5049 7113 5052
rect 7147 5049 7159 5083
rect 7576 5080 7604 5120
rect 7650 5108 7656 5160
rect 7708 5108 7714 5160
rect 8202 5108 8208 5160
rect 8260 5108 8266 5160
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 15580 5148 15608 5179
rect 15746 5176 15752 5188
rect 15804 5176 15810 5228
rect 15930 5176 15936 5228
rect 15988 5216 15994 5228
rect 18506 5216 18512 5228
rect 15988 5188 18512 5216
rect 15988 5176 15994 5188
rect 14976 5120 15608 5148
rect 14976 5108 14982 5120
rect 16298 5108 16304 5160
rect 16356 5108 16362 5160
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 16850 5108 16856 5160
rect 16908 5108 16914 5160
rect 16960 5157 16988 5188
rect 18506 5176 18512 5188
rect 18564 5176 18570 5228
rect 18616 5225 18644 5256
rect 18601 5219 18659 5225
rect 18601 5185 18613 5219
rect 18647 5185 18659 5219
rect 18601 5179 18659 5185
rect 16945 5151 17003 5157
rect 16945 5117 16957 5151
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17034 5108 17040 5160
rect 17092 5148 17098 5160
rect 17221 5151 17279 5157
rect 17221 5148 17233 5151
rect 17092 5120 17233 5148
rect 17092 5108 17098 5120
rect 17221 5117 17233 5120
rect 17267 5117 17279 5151
rect 17221 5111 17279 5117
rect 18046 5108 18052 5160
rect 18104 5108 18110 5160
rect 18138 5108 18144 5160
rect 18196 5157 18202 5160
rect 18196 5151 18245 5157
rect 18196 5117 18199 5151
rect 18233 5117 18245 5151
rect 18196 5111 18245 5117
rect 18196 5108 18202 5111
rect 18322 5108 18328 5160
rect 18380 5108 18386 5160
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 18984 5148 19012 5256
rect 20070 5244 20076 5256
rect 20128 5244 20134 5296
rect 19058 5176 19064 5228
rect 19116 5176 19122 5228
rect 19242 5176 19248 5228
rect 19300 5176 19306 5228
rect 20180 5216 20208 5324
rect 20901 5287 20959 5293
rect 20901 5253 20913 5287
rect 20947 5253 20959 5287
rect 21008 5284 21036 5324
rect 21085 5321 21097 5355
rect 21131 5352 21143 5355
rect 21266 5352 21272 5364
rect 21131 5324 21272 5352
rect 21131 5321 21143 5324
rect 21085 5315 21143 5321
rect 21266 5312 21272 5324
rect 21324 5312 21330 5364
rect 23934 5352 23940 5364
rect 21376 5324 23940 5352
rect 21376 5284 21404 5324
rect 23934 5312 23940 5324
rect 23992 5312 23998 5364
rect 24026 5312 24032 5364
rect 24084 5312 24090 5364
rect 24305 5355 24363 5361
rect 24305 5321 24317 5355
rect 24351 5352 24363 5355
rect 25590 5352 25596 5364
rect 24351 5324 25596 5352
rect 24351 5321 24363 5324
rect 24305 5315 24363 5321
rect 25590 5312 25596 5324
rect 25648 5312 25654 5364
rect 21008 5256 21404 5284
rect 21453 5287 21511 5293
rect 20901 5247 20959 5253
rect 21453 5253 21465 5287
rect 21499 5284 21511 5287
rect 21634 5284 21640 5296
rect 21499 5256 21640 5284
rect 21499 5253 21511 5256
rect 21453 5247 21511 5253
rect 20916 5216 20944 5247
rect 19352 5188 20208 5216
rect 20456 5188 20944 5216
rect 19352 5148 19380 5188
rect 20456 5157 20484 5188
rect 18932 5120 19380 5148
rect 20165 5151 20223 5157
rect 18932 5108 18938 5120
rect 20165 5117 20177 5151
rect 20211 5148 20223 5151
rect 20257 5151 20315 5157
rect 20257 5148 20269 5151
rect 20211 5120 20269 5148
rect 20211 5117 20223 5120
rect 20165 5111 20223 5117
rect 20257 5117 20269 5120
rect 20303 5117 20315 5151
rect 20257 5111 20315 5117
rect 20441 5151 20499 5157
rect 20441 5117 20453 5151
rect 20487 5117 20499 5151
rect 20441 5111 20499 5117
rect 20622 5108 20628 5160
rect 20680 5108 20686 5160
rect 20714 5108 20720 5160
rect 20772 5148 20778 5160
rect 21468 5148 21496 5247
rect 21634 5244 21640 5256
rect 21692 5244 21698 5296
rect 21542 5176 21548 5228
rect 21600 5216 21606 5228
rect 22094 5216 22100 5228
rect 21600 5188 22100 5216
rect 21600 5176 21606 5188
rect 22094 5176 22100 5188
rect 22152 5216 22158 5228
rect 22557 5219 22615 5225
rect 22557 5216 22569 5219
rect 22152 5188 22569 5216
rect 22152 5176 22158 5188
rect 22557 5185 22569 5188
rect 22603 5185 22615 5219
rect 22557 5179 22615 5185
rect 22833 5219 22891 5225
rect 22833 5185 22845 5219
rect 22879 5216 22891 5219
rect 24044 5216 24072 5312
rect 24762 5244 24768 5296
rect 24820 5244 24826 5296
rect 22879 5188 24072 5216
rect 22879 5185 22891 5188
rect 22833 5179 22891 5185
rect 24210 5176 24216 5228
rect 24268 5216 24274 5228
rect 24780 5216 24808 5244
rect 24268 5188 25176 5216
rect 24268 5176 24274 5188
rect 20772 5120 21496 5148
rect 21821 5151 21879 5157
rect 20772 5108 20778 5120
rect 21821 5117 21833 5151
rect 21867 5148 21879 5151
rect 22002 5148 22008 5160
rect 21867 5120 22008 5148
rect 21867 5117 21879 5120
rect 21821 5111 21879 5117
rect 22002 5108 22008 5120
rect 22060 5108 22066 5160
rect 22370 5108 22376 5160
rect 22428 5108 22434 5160
rect 24118 5108 24124 5160
rect 24176 5148 24182 5160
rect 24176 5120 24808 5148
rect 24176 5108 24182 5120
rect 8220 5080 8248 5108
rect 7576 5052 8248 5080
rect 7101 5043 7159 5049
rect 9674 5040 9680 5092
rect 9732 5040 9738 5092
rect 13538 5040 13544 5092
rect 13596 5040 13602 5092
rect 14737 5083 14795 5089
rect 14737 5049 14749 5083
rect 14783 5080 14795 5083
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 14783 5052 15761 5080
rect 14783 5049 14795 5052
rect 14737 5043 14795 5049
rect 15749 5049 15761 5052
rect 15795 5049 15807 5083
rect 21085 5083 21143 5089
rect 21085 5080 21097 5083
rect 15749 5043 15807 5049
rect 19260 5052 21097 5080
rect 5994 4972 6000 5024
rect 6052 5012 6058 5024
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 6052 4984 6377 5012
rect 6052 4972 6058 4984
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 6365 4975 6423 4981
rect 6549 5015 6607 5021
rect 6549 4981 6561 5015
rect 6595 5012 6607 5015
rect 6638 5012 6644 5024
rect 6595 4984 6644 5012
rect 6595 4981 6607 4984
rect 6549 4975 6607 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 10410 4972 10416 5024
rect 10468 4972 10474 5024
rect 13446 4972 13452 5024
rect 13504 5012 13510 5024
rect 14369 5015 14427 5021
rect 14369 5012 14381 5015
rect 13504 4984 14381 5012
rect 13504 4972 13510 4984
rect 14369 4981 14381 4984
rect 14415 4981 14427 5015
rect 14369 4975 14427 4981
rect 17405 5015 17463 5021
rect 17405 4981 17417 5015
rect 17451 5012 17463 5015
rect 19260 5012 19288 5052
rect 21085 5049 21097 5052
rect 21131 5049 21143 5083
rect 21085 5043 21143 5049
rect 21174 5040 21180 5092
rect 21232 5080 21238 5092
rect 24670 5080 24676 5092
rect 21232 5052 22094 5080
rect 24058 5052 24676 5080
rect 21232 5040 21238 5052
rect 17451 4984 19288 5012
rect 22066 5012 22094 5052
rect 24670 5040 24676 5052
rect 24728 5040 24734 5092
rect 23658 5012 23664 5024
rect 22066 4984 23664 5012
rect 17451 4981 17463 4984
rect 17405 4975 17463 4981
rect 23658 4972 23664 4984
rect 23716 4972 23722 5024
rect 23750 4972 23756 5024
rect 23808 5012 23814 5024
rect 24397 5015 24455 5021
rect 24397 5012 24409 5015
rect 23808 4984 24409 5012
rect 23808 4972 23814 4984
rect 24397 4981 24409 4984
rect 24443 4981 24455 5015
rect 24780 5012 24808 5120
rect 24946 5108 24952 5160
rect 25004 5108 25010 5160
rect 25148 5157 25176 5188
rect 25133 5151 25191 5157
rect 25133 5117 25145 5151
rect 25179 5117 25191 5151
rect 25133 5111 25191 5117
rect 30006 5108 30012 5160
rect 30064 5108 30070 5160
rect 24854 5040 24860 5092
rect 24912 5080 24918 5092
rect 25225 5083 25283 5089
rect 25225 5080 25237 5083
rect 24912 5052 25237 5080
rect 24912 5040 24918 5052
rect 25225 5049 25237 5052
rect 25271 5049 25283 5083
rect 25225 5043 25283 5049
rect 28534 5012 28540 5024
rect 24780 4984 28540 5012
rect 24397 4975 24455 4981
rect 28534 4972 28540 4984
rect 28592 4972 28598 5024
rect 29454 4972 29460 5024
rect 29512 4972 29518 5024
rect 2760 4922 32200 4944
rect 2760 4870 6946 4922
rect 6998 4870 7010 4922
rect 7062 4870 7074 4922
rect 7126 4870 7138 4922
rect 7190 4870 7202 4922
rect 7254 4870 14306 4922
rect 14358 4870 14370 4922
rect 14422 4870 14434 4922
rect 14486 4870 14498 4922
rect 14550 4870 14562 4922
rect 14614 4870 21666 4922
rect 21718 4870 21730 4922
rect 21782 4870 21794 4922
rect 21846 4870 21858 4922
rect 21910 4870 21922 4922
rect 21974 4870 29026 4922
rect 29078 4870 29090 4922
rect 29142 4870 29154 4922
rect 29206 4870 29218 4922
rect 29270 4870 29282 4922
rect 29334 4870 32200 4922
rect 2760 4848 32200 4870
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4488 4780 4629 4808
rect 4488 4768 4494 4780
rect 4617 4777 4629 4780
rect 4663 4808 4675 4811
rect 5350 4808 5356 4820
rect 4663 4780 5356 4808
rect 4663 4777 4675 4780
rect 4617 4771 4675 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 6822 4768 6828 4820
rect 6880 4768 6886 4820
rect 6917 4811 6975 4817
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 6963 4780 7880 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 7852 4749 7880 4780
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 9769 4811 9827 4817
rect 9769 4808 9781 4811
rect 9732 4780 9781 4808
rect 9732 4768 9738 4780
rect 9769 4777 9781 4780
rect 9815 4777 9827 4811
rect 9769 4771 9827 4777
rect 10226 4768 10232 4820
rect 10284 4768 10290 4820
rect 12250 4768 12256 4820
rect 12308 4808 12314 4820
rect 12529 4811 12587 4817
rect 12529 4808 12541 4811
rect 12308 4780 12541 4808
rect 12308 4768 12314 4780
rect 12529 4777 12541 4780
rect 12575 4777 12587 4811
rect 12529 4771 12587 4777
rect 7377 4743 7435 4749
rect 7377 4740 7389 4743
rect 5658 4712 7389 4740
rect 7377 4709 7389 4712
rect 7423 4709 7435 4743
rect 7377 4703 7435 4709
rect 7837 4743 7895 4749
rect 7837 4709 7849 4743
rect 7883 4740 7895 4743
rect 10244 4740 10272 4768
rect 7883 4712 10272 4740
rect 12544 4740 12572 4771
rect 12986 4768 12992 4820
rect 13044 4768 13050 4820
rect 13538 4768 13544 4820
rect 13596 4768 13602 4820
rect 13630 4768 13636 4820
rect 13688 4808 13694 4820
rect 14277 4811 14335 4817
rect 14277 4808 14289 4811
rect 13688 4780 14289 4808
rect 13688 4768 13694 4780
rect 14277 4777 14289 4780
rect 14323 4777 14335 4811
rect 14277 4771 14335 4777
rect 14645 4811 14703 4817
rect 14645 4777 14657 4811
rect 14691 4808 14703 4811
rect 15286 4808 15292 4820
rect 14691 4780 15292 4808
rect 14691 4777 14703 4780
rect 14645 4771 14703 4777
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 17405 4811 17463 4817
rect 17405 4777 17417 4811
rect 17451 4808 17463 4811
rect 17494 4808 17500 4820
rect 17451 4780 17500 4808
rect 17451 4777 17463 4780
rect 17405 4771 17463 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 19058 4808 19064 4820
rect 18340 4780 19064 4808
rect 14185 4743 14243 4749
rect 12544 4712 14136 4740
rect 7883 4709 7895 4712
rect 7837 4703 7895 4709
rect 7469 4675 7527 4681
rect 7469 4641 7481 4675
rect 7515 4672 7527 4675
rect 8202 4672 8208 4684
rect 7515 4644 8208 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 8202 4632 8208 4644
rect 8260 4672 8266 4684
rect 9677 4675 9735 4681
rect 9677 4672 9689 4675
rect 8260 4644 9689 4672
rect 8260 4632 8266 4644
rect 9677 4641 9689 4644
rect 9723 4672 9735 4675
rect 13449 4675 13507 4681
rect 13449 4672 13461 4675
rect 9723 4644 13461 4672
rect 9723 4641 9735 4644
rect 9677 4635 9735 4641
rect 13449 4641 13461 4644
rect 13495 4641 13507 4675
rect 14108 4672 14136 4712
rect 14185 4709 14197 4743
rect 14231 4740 14243 4743
rect 15473 4743 15531 4749
rect 15473 4740 15485 4743
rect 14231 4712 15485 4740
rect 14231 4709 14243 4712
rect 14185 4703 14243 4709
rect 15473 4709 15485 4712
rect 15519 4709 15531 4743
rect 15473 4703 15531 4709
rect 15013 4675 15071 4681
rect 14108 4644 14412 4672
rect 13449 4635 13507 4641
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 6052 4576 6101 4604
rect 6052 4564 6058 4576
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6089 4567 6147 4573
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 6086 4428 6092 4480
rect 6144 4468 6150 4480
rect 6380 4468 6408 4567
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6788 4576 7021 4604
rect 6788 4564 6794 4576
rect 7009 4573 7021 4576
rect 7055 4573 7067 4607
rect 13464 4604 13492 4635
rect 13538 4604 13544 4616
rect 13464 4576 13544 4604
rect 7009 4567 7067 4573
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 13998 4564 14004 4616
rect 14056 4604 14062 4616
rect 14182 4604 14188 4616
rect 14056 4576 14188 4604
rect 14056 4564 14062 4576
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14384 4613 14412 4644
rect 15013 4641 15025 4675
rect 15059 4672 15071 4675
rect 15562 4672 15568 4684
rect 15059 4644 15568 4672
rect 15059 4641 15071 4644
rect 15013 4635 15071 4641
rect 15562 4632 15568 4644
rect 15620 4632 15626 4684
rect 16390 4672 16396 4684
rect 16040 4644 16396 4672
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14384 4536 14412 4567
rect 15102 4564 15108 4616
rect 15160 4564 15166 4616
rect 15194 4564 15200 4616
rect 15252 4604 15258 4616
rect 16040 4604 16068 4644
rect 16390 4632 16396 4644
rect 16448 4672 16454 4684
rect 17313 4675 17371 4681
rect 16448 4644 17080 4672
rect 16448 4632 16454 4644
rect 15252 4576 16068 4604
rect 15252 4564 15258 4576
rect 16114 4564 16120 4616
rect 16172 4564 16178 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 17052 4604 17080 4644
rect 17313 4641 17325 4675
rect 17359 4672 17371 4675
rect 18046 4672 18052 4684
rect 17359 4644 18052 4672
rect 17359 4641 17371 4644
rect 17313 4635 17371 4641
rect 18046 4632 18052 4644
rect 18104 4632 18110 4684
rect 18141 4675 18199 4681
rect 18141 4641 18153 4675
rect 18187 4672 18199 4675
rect 18230 4672 18236 4684
rect 18187 4644 18236 4672
rect 18187 4641 18199 4644
rect 18141 4635 18199 4641
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 18340 4681 18368 4780
rect 19058 4768 19064 4780
rect 19116 4808 19122 4820
rect 21174 4808 21180 4820
rect 19116 4780 21180 4808
rect 19116 4768 19122 4780
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 21450 4768 21456 4820
rect 21508 4768 21514 4820
rect 22002 4768 22008 4820
rect 22060 4768 22066 4820
rect 23293 4811 23351 4817
rect 23293 4777 23305 4811
rect 23339 4777 23351 4811
rect 23293 4771 23351 4777
rect 18414 4700 18420 4752
rect 18472 4740 18478 4752
rect 18509 4743 18567 4749
rect 18509 4740 18521 4743
rect 18472 4712 18521 4740
rect 18472 4700 18478 4712
rect 18509 4709 18521 4712
rect 18555 4709 18567 4743
rect 18966 4740 18972 4752
rect 18509 4703 18567 4709
rect 18616 4712 18972 4740
rect 18616 4681 18644 4712
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 19794 4700 19800 4752
rect 19852 4740 19858 4752
rect 21269 4743 21327 4749
rect 21269 4740 21281 4743
rect 19852 4712 21281 4740
rect 19852 4700 19858 4712
rect 21269 4709 21281 4712
rect 21315 4709 21327 4743
rect 21269 4703 21327 4709
rect 18325 4675 18383 4681
rect 18325 4641 18337 4675
rect 18371 4641 18383 4675
rect 18325 4635 18383 4641
rect 18601 4675 18659 4681
rect 18601 4641 18613 4675
rect 18647 4641 18659 4675
rect 18601 4635 18659 4641
rect 18690 4632 18696 4684
rect 18748 4632 18754 4684
rect 20714 4672 20720 4684
rect 18800 4644 19104 4672
rect 17497 4607 17555 4613
rect 17497 4604 17509 4607
rect 16899 4576 16988 4604
rect 17052 4576 17509 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 15212 4536 15240 4564
rect 16960 4545 16988 4576
rect 17497 4573 17509 4576
rect 17543 4604 17555 4607
rect 18800 4604 18828 4644
rect 18969 4607 19027 4613
rect 18969 4604 18981 4607
rect 17543 4576 18828 4604
rect 18892 4576 18981 4604
rect 17543 4573 17555 4576
rect 17497 4567 17555 4573
rect 18892 4545 18920 4576
rect 18969 4573 18981 4576
rect 19015 4573 19027 4607
rect 19076 4604 19104 4644
rect 19306 4644 20720 4672
rect 19306 4604 19334 4644
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 21361 4675 21419 4681
rect 21361 4641 21373 4675
rect 21407 4672 21419 4675
rect 21468 4672 21496 4768
rect 21821 4743 21879 4749
rect 21821 4709 21833 4743
rect 21867 4740 21879 4743
rect 22020 4740 22048 4768
rect 23106 4740 23112 4752
rect 21867 4712 22048 4740
rect 23046 4712 23112 4740
rect 21867 4709 21879 4712
rect 21821 4703 21879 4709
rect 23106 4700 23112 4712
rect 23164 4700 23170 4752
rect 23308 4740 23336 4771
rect 23566 4768 23572 4820
rect 23624 4768 23630 4820
rect 23934 4768 23940 4820
rect 23992 4808 23998 4820
rect 28997 4811 29055 4817
rect 23992 4780 27660 4808
rect 23992 4768 23998 4780
rect 24946 4740 24952 4752
rect 23308 4712 24952 4740
rect 24946 4700 24952 4712
rect 25004 4700 25010 4752
rect 27632 4740 27660 4780
rect 28997 4777 29009 4811
rect 29043 4808 29055 4811
rect 29454 4808 29460 4820
rect 29043 4780 29460 4808
rect 29043 4777 29055 4780
rect 28997 4771 29055 4777
rect 29454 4768 29460 4780
rect 29512 4768 29518 4820
rect 29730 4768 29736 4820
rect 29788 4808 29794 4820
rect 30009 4811 30067 4817
rect 30009 4808 30021 4811
rect 29788 4780 30021 4808
rect 29788 4768 29794 4780
rect 30009 4777 30021 4780
rect 30055 4777 30067 4811
rect 30009 4771 30067 4777
rect 29641 4743 29699 4749
rect 29641 4740 29653 4743
rect 27632 4712 29653 4740
rect 29641 4709 29653 4712
rect 29687 4709 29699 4743
rect 29641 4703 29699 4709
rect 21407 4644 21496 4672
rect 21407 4641 21419 4644
rect 21361 4635 21419 4641
rect 21542 4632 21548 4684
rect 21600 4632 21606 4684
rect 23474 4632 23480 4684
rect 23532 4672 23538 4684
rect 23661 4675 23719 4681
rect 23661 4672 23673 4675
rect 23532 4644 23673 4672
rect 23532 4632 23538 4644
rect 23661 4641 23673 4644
rect 23707 4672 23719 4675
rect 24118 4672 24124 4684
rect 23707 4644 24124 4672
rect 23707 4641 23719 4644
rect 23661 4635 23719 4641
rect 24118 4632 24124 4644
rect 24176 4632 24182 4684
rect 24305 4675 24363 4681
rect 24305 4641 24317 4675
rect 24351 4641 24363 4675
rect 24305 4635 24363 4641
rect 19076 4576 19334 4604
rect 18969 4567 19027 4573
rect 19426 4564 19432 4616
rect 19484 4604 19490 4616
rect 19705 4607 19763 4613
rect 19705 4604 19717 4607
rect 19484 4576 19717 4604
rect 19484 4564 19490 4576
rect 19705 4573 19717 4576
rect 19751 4573 19763 4607
rect 19705 4567 19763 4573
rect 20346 4564 20352 4616
rect 20404 4604 20410 4616
rect 20993 4607 21051 4613
rect 20993 4604 21005 4607
rect 20404 4576 21005 4604
rect 20404 4564 20410 4576
rect 20993 4573 21005 4576
rect 21039 4573 21051 4607
rect 20993 4567 21051 4573
rect 24026 4564 24032 4616
rect 24084 4564 24090 4616
rect 24213 4607 24271 4613
rect 24213 4573 24225 4607
rect 24259 4573 24271 4607
rect 24213 4567 24271 4573
rect 14384 4508 15240 4536
rect 16945 4539 17003 4545
rect 16945 4505 16957 4539
rect 16991 4505 17003 4539
rect 16945 4499 17003 4505
rect 18877 4539 18935 4545
rect 18877 4505 18889 4539
rect 18923 4505 18935 4539
rect 18877 4499 18935 4505
rect 19242 4496 19248 4548
rect 19300 4536 19306 4548
rect 24228 4536 24256 4567
rect 19300 4508 21680 4536
rect 19300 4496 19306 4508
rect 6144 4440 6408 4468
rect 6457 4471 6515 4477
rect 6144 4428 6150 4440
rect 6457 4437 6469 4471
rect 6503 4468 6515 4471
rect 6730 4468 6736 4480
rect 6503 4440 6736 4468
rect 6503 4437 6515 4440
rect 6457 4431 6515 4437
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 13817 4471 13875 4477
rect 13817 4437 13829 4471
rect 13863 4468 13875 4471
rect 13998 4468 14004 4480
rect 13863 4440 14004 4468
rect 13863 4437 13875 4440
rect 13817 4431 13875 4437
rect 13998 4428 14004 4440
rect 14056 4428 14062 4480
rect 16206 4428 16212 4480
rect 16264 4428 16270 4480
rect 18049 4471 18107 4477
rect 18049 4437 18061 4471
rect 18095 4468 18107 4471
rect 19518 4468 19524 4480
rect 18095 4440 19524 4468
rect 18095 4437 18107 4440
rect 18049 4431 18107 4437
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19610 4428 19616 4480
rect 19668 4428 19674 4480
rect 20254 4428 20260 4480
rect 20312 4468 20318 4480
rect 20349 4471 20407 4477
rect 20349 4468 20361 4471
rect 20312 4440 20361 4468
rect 20312 4428 20318 4440
rect 20349 4437 20361 4440
rect 20395 4437 20407 4471
rect 20349 4431 20407 4437
rect 20438 4428 20444 4480
rect 20496 4428 20502 4480
rect 21652 4468 21680 4508
rect 23400 4508 24256 4536
rect 23400 4480 23428 4508
rect 23382 4468 23388 4480
rect 21652 4440 23388 4468
rect 23382 4428 23388 4440
rect 23440 4428 23446 4480
rect 23566 4428 23572 4480
rect 23624 4468 23630 4480
rect 24320 4468 24348 4635
rect 24486 4632 24492 4684
rect 24544 4672 24550 4684
rect 28261 4675 28319 4681
rect 28261 4672 28273 4675
rect 24544 4644 28273 4672
rect 24544 4632 24550 4644
rect 28261 4641 28273 4644
rect 28307 4641 28319 4675
rect 28261 4635 28319 4641
rect 24765 4607 24823 4613
rect 24765 4604 24777 4607
rect 24688 4576 24777 4604
rect 24688 4545 24716 4576
rect 24765 4573 24777 4576
rect 24811 4573 24823 4607
rect 28276 4604 28304 4635
rect 28534 4632 28540 4684
rect 28592 4672 28598 4684
rect 28592 4644 29224 4672
rect 28592 4632 28598 4644
rect 29196 4613 29224 4644
rect 29089 4607 29147 4613
rect 29089 4604 29101 4607
rect 28276 4576 29101 4604
rect 24765 4567 24823 4573
rect 29089 4573 29101 4576
rect 29135 4573 29147 4607
rect 29089 4567 29147 4573
rect 29181 4607 29239 4613
rect 29181 4573 29193 4607
rect 29227 4573 29239 4607
rect 29656 4604 29684 4703
rect 30834 4681 30840 4684
rect 30812 4675 30840 4681
rect 30812 4641 30824 4675
rect 30812 4635 30840 4641
rect 30834 4632 30840 4635
rect 30892 4632 30898 4684
rect 29656 4576 30236 4604
rect 29181 4567 29239 4573
rect 24673 4539 24731 4545
rect 24673 4505 24685 4539
rect 24719 4505 24731 4539
rect 24673 4499 24731 4505
rect 23624 4440 24348 4468
rect 23624 4428 23630 4440
rect 25406 4428 25412 4480
rect 25464 4428 25470 4480
rect 28258 4428 28264 4480
rect 28316 4468 28322 4480
rect 28629 4471 28687 4477
rect 28629 4468 28641 4471
rect 28316 4440 28641 4468
rect 28316 4428 28322 4440
rect 28629 4437 28641 4440
rect 28675 4437 28687 4471
rect 30208 4468 30236 4576
rect 30466 4564 30472 4616
rect 30524 4604 30530 4616
rect 30653 4607 30711 4613
rect 30653 4604 30665 4607
rect 30524 4576 30665 4604
rect 30524 4564 30530 4576
rect 30653 4573 30665 4576
rect 30699 4573 30711 4607
rect 30653 4567 30711 4573
rect 30926 4564 30932 4616
rect 30984 4564 30990 4616
rect 31662 4564 31668 4616
rect 31720 4564 31726 4616
rect 31846 4564 31852 4616
rect 31904 4564 31910 4616
rect 31205 4539 31263 4545
rect 31205 4505 31217 4539
rect 31251 4505 31263 4539
rect 31205 4499 31263 4505
rect 31220 4468 31248 4499
rect 30208 4440 31248 4468
rect 28629 4431 28687 4437
rect 2760 4378 32200 4400
rect 2760 4326 6286 4378
rect 6338 4326 6350 4378
rect 6402 4326 6414 4378
rect 6466 4326 6478 4378
rect 6530 4326 6542 4378
rect 6594 4326 13646 4378
rect 13698 4326 13710 4378
rect 13762 4326 13774 4378
rect 13826 4326 13838 4378
rect 13890 4326 13902 4378
rect 13954 4326 21006 4378
rect 21058 4326 21070 4378
rect 21122 4326 21134 4378
rect 21186 4326 21198 4378
rect 21250 4326 21262 4378
rect 21314 4326 28366 4378
rect 28418 4326 28430 4378
rect 28482 4326 28494 4378
rect 28546 4326 28558 4378
rect 28610 4326 28622 4378
rect 28674 4326 32200 4378
rect 2760 4304 32200 4326
rect 5708 4267 5766 4273
rect 5708 4233 5720 4267
rect 5754 4264 5766 4267
rect 6730 4264 6736 4276
rect 5754 4236 6736 4264
rect 5754 4233 5766 4236
rect 5708 4227 5766 4233
rect 6730 4224 6736 4236
rect 6788 4224 6794 4276
rect 7193 4267 7251 4273
rect 7193 4233 7205 4267
rect 7239 4264 7251 4267
rect 7650 4264 7656 4276
rect 7239 4236 7656 4264
rect 7239 4233 7251 4236
rect 7193 4227 7251 4233
rect 7650 4224 7656 4236
rect 7708 4224 7714 4276
rect 12240 4267 12298 4273
rect 12240 4233 12252 4267
rect 12286 4264 12298 4267
rect 13446 4264 13452 4276
rect 12286 4236 13452 4264
rect 12286 4233 12298 4236
rect 12240 4227 12298 4233
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 14080 4267 14138 4273
rect 14080 4233 14092 4267
rect 14126 4264 14138 4267
rect 14642 4264 14648 4276
rect 14126 4236 14648 4264
rect 14126 4233 14138 4236
rect 14080 4227 14138 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 15212 4236 15424 4264
rect 5445 4131 5503 4137
rect 5445 4097 5457 4131
rect 5491 4128 5503 4131
rect 6086 4128 6092 4140
rect 5491 4100 6092 4128
rect 5491 4097 5503 4100
rect 5445 4091 5503 4097
rect 6086 4088 6092 4100
rect 6144 4088 6150 4140
rect 11977 4131 12035 4137
rect 11977 4097 11989 4131
rect 12023 4128 12035 4131
rect 12618 4128 12624 4140
rect 12023 4100 12624 4128
rect 12023 4097 12035 4100
rect 11977 4091 12035 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 13817 4131 13875 4137
rect 13817 4097 13829 4131
rect 13863 4128 13875 4131
rect 14090 4128 14096 4140
rect 13863 4100 14096 4128
rect 13863 4097 13875 4100
rect 13817 4091 13875 4097
rect 14090 4088 14096 4100
rect 14148 4128 14154 4140
rect 15212 4128 15240 4236
rect 14148 4100 15240 4128
rect 15396 4128 15424 4236
rect 16206 4224 16212 4276
rect 16264 4264 16270 4276
rect 16558 4267 16616 4273
rect 16558 4264 16570 4267
rect 16264 4236 16570 4264
rect 16264 4224 16270 4236
rect 16558 4233 16570 4236
rect 16604 4233 16616 4267
rect 16558 4227 16616 4233
rect 18046 4224 18052 4276
rect 18104 4224 18110 4276
rect 18874 4264 18880 4276
rect 18156 4236 18880 4264
rect 17586 4156 17592 4208
rect 17644 4196 17650 4208
rect 18156 4196 18184 4236
rect 18874 4224 18880 4236
rect 18932 4224 18938 4276
rect 19048 4267 19106 4273
rect 19048 4233 19060 4267
rect 19094 4264 19106 4267
rect 19610 4264 19616 4276
rect 19094 4236 19616 4264
rect 19094 4233 19106 4236
rect 19048 4227 19106 4233
rect 19610 4224 19616 4236
rect 19668 4224 19674 4276
rect 20070 4224 20076 4276
rect 20128 4264 20134 4276
rect 20128 4236 23336 4264
rect 20128 4224 20134 4236
rect 18414 4196 18420 4208
rect 17644 4168 18184 4196
rect 18340 4168 18420 4196
rect 17644 4156 17650 4168
rect 16301 4131 16359 4137
rect 16301 4128 16313 4131
rect 15396 4100 16313 4128
rect 14148 4088 14154 4100
rect 16301 4097 16313 4100
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 3050 4020 3056 4072
rect 3108 4020 3114 4072
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 2590 3952 2596 4004
rect 2648 3992 2654 4004
rect 3344 3992 3372 4023
rect 15470 4020 15476 4072
rect 15528 4060 15534 4072
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15528 4032 15945 4060
rect 15528 4020 15534 4032
rect 15933 4029 15945 4032
rect 15979 4060 15991 4063
rect 16209 4063 16267 4069
rect 16209 4060 16221 4063
rect 15979 4032 16221 4060
rect 15979 4029 15991 4032
rect 15933 4023 15991 4029
rect 16209 4029 16221 4032
rect 16255 4029 16267 4063
rect 16209 4023 16267 4029
rect 2648 3964 3372 3992
rect 3436 3964 6132 3992
rect 2648 3952 2654 3964
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3436 3924 3464 3964
rect 3283 3896 3464 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3510 3884 3516 3936
rect 3568 3884 3574 3936
rect 6104 3924 6132 3964
rect 6730 3952 6736 4004
rect 6788 3952 6794 4004
rect 13538 3992 13544 4004
rect 13478 3964 13544 3992
rect 13538 3952 13544 3964
rect 13596 3952 13602 4004
rect 16117 3995 16175 4001
rect 16117 3992 16129 3995
rect 15318 3964 16129 3992
rect 16117 3961 16129 3964
rect 16163 3961 16175 3995
rect 16224 3992 16252 4023
rect 17954 4020 17960 4072
rect 18012 4060 18018 4072
rect 18141 4063 18199 4069
rect 18141 4060 18153 4063
rect 18012 4032 18153 4060
rect 18012 4020 18018 4032
rect 18141 4029 18153 4032
rect 18187 4060 18199 4063
rect 18230 4060 18236 4072
rect 18187 4032 18236 4060
rect 18187 4029 18199 4032
rect 18141 4023 18199 4029
rect 18230 4020 18236 4032
rect 18288 4020 18294 4072
rect 18340 4069 18368 4168
rect 18414 4156 18420 4168
rect 18472 4156 18478 4208
rect 23308 4196 23336 4236
rect 23382 4224 23388 4276
rect 23440 4224 23446 4276
rect 25059 4267 25117 4273
rect 25059 4233 25071 4267
rect 25105 4264 25117 4267
rect 25406 4264 25412 4276
rect 25105 4236 25412 4264
rect 25105 4233 25117 4236
rect 25059 4227 25117 4233
rect 25406 4224 25412 4236
rect 25464 4224 25470 4276
rect 29825 4267 29883 4273
rect 29825 4233 29837 4267
rect 29871 4264 29883 4267
rect 30006 4264 30012 4276
rect 29871 4236 30012 4264
rect 29871 4233 29883 4236
rect 29825 4227 29883 4233
rect 30006 4224 30012 4236
rect 30064 4224 30070 4276
rect 31573 4267 31631 4273
rect 31573 4233 31585 4267
rect 31619 4264 31631 4267
rect 31662 4264 31668 4276
rect 31619 4236 31668 4264
rect 31619 4233 31631 4236
rect 31573 4227 31631 4233
rect 31662 4224 31668 4236
rect 31720 4224 31726 4276
rect 30377 4199 30435 4205
rect 30377 4196 30389 4199
rect 18708 4168 18920 4196
rect 23308 4168 24072 4196
rect 18708 4128 18736 4168
rect 18432 4100 18736 4128
rect 18432 4069 18460 4100
rect 18782 4088 18788 4140
rect 18840 4088 18846 4140
rect 18892 4128 18920 4168
rect 20254 4128 20260 4140
rect 18892 4100 20260 4128
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 20898 4088 20904 4140
rect 20956 4128 20962 4140
rect 21542 4128 21548 4140
rect 20956 4100 21548 4128
rect 20956 4088 20962 4100
rect 21542 4088 21548 4100
rect 21600 4088 21606 4140
rect 21818 4088 21824 4140
rect 21876 4128 21882 4140
rect 22741 4131 22799 4137
rect 22741 4128 22753 4131
rect 21876 4100 22753 4128
rect 21876 4088 21882 4100
rect 22741 4097 22753 4100
rect 22787 4097 22799 4131
rect 24044 4128 24072 4168
rect 25240 4168 28212 4196
rect 25240 4128 25268 4168
rect 24044 4100 25268 4128
rect 25317 4131 25375 4137
rect 22741 4091 22799 4097
rect 25317 4097 25329 4131
rect 25363 4128 25375 4131
rect 27614 4128 27620 4140
rect 25363 4100 27620 4128
rect 25363 4097 25375 4100
rect 25317 4091 25375 4097
rect 27614 4088 27620 4100
rect 27672 4128 27678 4140
rect 28077 4131 28135 4137
rect 28077 4128 28089 4131
rect 27672 4100 28089 4128
rect 27672 4088 27678 4100
rect 28077 4097 28089 4100
rect 28123 4097 28135 4131
rect 28184 4128 28212 4168
rect 29380 4168 30389 4196
rect 29380 4128 29408 4168
rect 30377 4165 30389 4168
rect 30423 4196 30435 4199
rect 30466 4196 30472 4208
rect 30423 4168 30472 4196
rect 30423 4165 30435 4168
rect 30377 4159 30435 4165
rect 30466 4156 30472 4168
rect 30524 4156 30530 4208
rect 33042 4128 33048 4140
rect 28184 4100 29408 4128
rect 31864 4100 33048 4128
rect 28077 4091 28135 4097
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4029 18383 4063
rect 18325 4023 18383 4029
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4029 18475 4063
rect 18417 4023 18475 4029
rect 18509 4063 18567 4069
rect 18509 4029 18521 4063
rect 18555 4060 18567 4063
rect 18690 4060 18696 4072
rect 18555 4032 18696 4060
rect 18555 4029 18567 4032
rect 18509 4023 18567 4029
rect 18690 4020 18696 4032
rect 18748 4020 18754 4072
rect 31864 4069 31892 4100
rect 33042 4088 33048 4100
rect 33100 4088 33106 4140
rect 25593 4063 25651 4069
rect 17862 3992 17868 4004
rect 16224 3964 16988 3992
rect 17802 3964 17868 3992
rect 16117 3955 16175 3961
rect 16960 3936 16988 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 19518 3952 19524 4004
rect 19576 3952 19582 4004
rect 20346 3952 20352 4004
rect 20404 3952 20410 4004
rect 21174 3952 21180 4004
rect 21232 3952 21238 4004
rect 11698 3924 11704 3936
rect 6104 3896 11704 3924
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 13725 3927 13783 3933
rect 13725 3893 13737 3927
rect 13771 3924 13783 3927
rect 15378 3924 15384 3936
rect 13771 3896 15384 3924
rect 13771 3893 13783 3896
rect 13725 3887 13783 3893
rect 15378 3884 15384 3896
rect 15436 3884 15442 3936
rect 15562 3884 15568 3936
rect 15620 3884 15626 3936
rect 15838 3884 15844 3936
rect 15896 3884 15902 3936
rect 16942 3884 16948 3936
rect 17000 3884 17006 3936
rect 18693 3927 18751 3933
rect 18693 3893 18705 3927
rect 18739 3924 18751 3927
rect 20364 3924 20392 3952
rect 18739 3896 20392 3924
rect 20533 3927 20591 3933
rect 18739 3893 18751 3896
rect 18693 3887 18751 3893
rect 20533 3893 20545 3927
rect 20579 3924 20591 3927
rect 21818 3924 21824 3936
rect 20579 3896 21824 3924
rect 20579 3893 20591 3896
rect 20533 3887 20591 3893
rect 21818 3884 21824 3896
rect 21876 3884 21882 3936
rect 22186 3884 22192 3936
rect 22244 3924 22250 3936
rect 22296 3924 22324 4046
rect 25593 4029 25605 4063
rect 25639 4029 25651 4063
rect 25593 4023 25651 4029
rect 30101 4063 30159 4069
rect 30101 4029 30113 4063
rect 30147 4029 30159 4063
rect 30101 4023 30159 4029
rect 31389 4063 31447 4069
rect 31389 4029 31401 4063
rect 31435 4060 31447 4063
rect 31849 4063 31907 4069
rect 31435 4032 31754 4060
rect 31435 4029 31447 4032
rect 31389 4023 31447 4029
rect 25501 3995 25559 4001
rect 24610 3964 24716 3992
rect 22244 3896 22324 3924
rect 22649 3927 22707 3933
rect 22244 3884 22250 3896
rect 22649 3893 22661 3927
rect 22695 3924 22707 3927
rect 23474 3924 23480 3936
rect 22695 3896 23480 3924
rect 22695 3893 22707 3896
rect 22649 3887 22707 3893
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 23566 3884 23572 3936
rect 23624 3884 23630 3936
rect 24688 3924 24716 3964
rect 25501 3961 25513 3995
rect 25547 3961 25559 3995
rect 25608 3992 25636 4023
rect 25608 3964 28212 3992
rect 25501 3955 25559 3961
rect 25516 3924 25544 3955
rect 28184 3936 28212 3964
rect 28258 3952 28264 4004
rect 28316 3992 28322 4004
rect 28353 3995 28411 4001
rect 28353 3992 28365 3995
rect 28316 3964 28365 3992
rect 28316 3952 28322 3964
rect 28353 3961 28365 3964
rect 28399 3961 28411 3995
rect 30009 3995 30067 4001
rect 30009 3992 30021 3995
rect 29578 3964 30021 3992
rect 28353 3955 28411 3961
rect 30009 3961 30021 3964
rect 30055 3961 30067 3995
rect 30009 3955 30067 3961
rect 24688 3896 25544 3924
rect 28166 3884 28172 3936
rect 28224 3924 28230 3936
rect 30116 3924 30144 4023
rect 31726 3992 31754 4032
rect 31849 4029 31861 4063
rect 31895 4029 31907 4063
rect 31849 4023 31907 4029
rect 33502 3992 33508 4004
rect 31726 3964 33508 3992
rect 33502 3952 33508 3964
rect 33560 3952 33566 4004
rect 28224 3896 30144 3924
rect 28224 3884 28230 3896
rect 31294 3884 31300 3936
rect 31352 3924 31358 3936
rect 31665 3927 31723 3933
rect 31665 3924 31677 3927
rect 31352 3896 31677 3924
rect 31352 3884 31358 3896
rect 31665 3893 31677 3896
rect 31711 3893 31723 3927
rect 31665 3887 31723 3893
rect 2760 3834 32200 3856
rect 2760 3782 6946 3834
rect 6998 3782 7010 3834
rect 7062 3782 7074 3834
rect 7126 3782 7138 3834
rect 7190 3782 7202 3834
rect 7254 3782 14306 3834
rect 14358 3782 14370 3834
rect 14422 3782 14434 3834
rect 14486 3782 14498 3834
rect 14550 3782 14562 3834
rect 14614 3782 21666 3834
rect 21718 3782 21730 3834
rect 21782 3782 21794 3834
rect 21846 3782 21858 3834
rect 21910 3782 21922 3834
rect 21974 3782 29026 3834
rect 29078 3782 29090 3834
rect 29142 3782 29154 3834
rect 29206 3782 29218 3834
rect 29270 3782 29282 3834
rect 29334 3782 32200 3834
rect 2760 3760 32200 3782
rect 3510 3680 3516 3732
rect 3568 3720 3574 3732
rect 13354 3720 13360 3732
rect 3568 3692 13360 3720
rect 3568 3680 3574 3692
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13538 3680 13544 3732
rect 13596 3720 13602 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13596 3692 13737 3720
rect 13596 3680 13602 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 13998 3680 14004 3732
rect 14056 3720 14062 3732
rect 14056 3692 14228 3720
rect 14056 3680 14062 3692
rect 6365 3655 6423 3661
rect 6365 3621 6377 3655
rect 6411 3652 6423 3655
rect 6822 3652 6828 3664
rect 6411 3624 6828 3652
rect 6411 3621 6423 3624
rect 6365 3615 6423 3621
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 14200 3661 14228 3692
rect 16022 3680 16028 3732
rect 16080 3720 16086 3732
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 16080 3692 16221 3720
rect 16080 3680 16086 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 16669 3723 16727 3729
rect 16669 3720 16681 3723
rect 16632 3692 16681 3720
rect 16632 3680 16638 3692
rect 16669 3689 16681 3692
rect 16715 3720 16727 3723
rect 17586 3720 17592 3732
rect 16715 3692 17592 3720
rect 16715 3689 16727 3692
rect 16669 3683 16727 3689
rect 17586 3680 17592 3692
rect 17644 3680 17650 3732
rect 17862 3680 17868 3732
rect 17920 3720 17926 3732
rect 18417 3723 18475 3729
rect 18417 3720 18429 3723
rect 17920 3692 18429 3720
rect 17920 3680 17926 3692
rect 18417 3689 18429 3692
rect 18463 3689 18475 3723
rect 18417 3683 18475 3689
rect 18785 3723 18843 3729
rect 18785 3689 18797 3723
rect 18831 3720 18843 3723
rect 19426 3720 19432 3732
rect 18831 3692 19432 3720
rect 18831 3689 18843 3692
rect 18785 3683 18843 3689
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 20438 3720 20444 3732
rect 20272 3692 20444 3720
rect 14185 3655 14243 3661
rect 12636 3624 13952 3652
rect 12636 3596 12664 3624
rect 4246 3544 4252 3596
rect 4304 3544 4310 3596
rect 5718 3544 5724 3596
rect 5776 3584 5782 3596
rect 5813 3587 5871 3593
rect 5813 3584 5825 3587
rect 5776 3556 5825 3584
rect 5776 3544 5782 3556
rect 5813 3553 5825 3556
rect 5859 3553 5871 3587
rect 5813 3547 5871 3553
rect 10410 3544 10416 3596
rect 10468 3544 10474 3596
rect 12618 3544 12624 3596
rect 12676 3544 12682 3596
rect 13630 3544 13636 3596
rect 13688 3584 13694 3596
rect 13817 3587 13875 3593
rect 13817 3584 13829 3587
rect 13688 3556 13829 3584
rect 13688 3544 13694 3556
rect 13817 3553 13829 3556
rect 13863 3553 13875 3587
rect 13817 3547 13875 3553
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 1360 3488 3249 3516
rect 1360 3476 1366 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4801 3519 4859 3525
rect 4801 3516 4813 3519
rect 4580 3488 4813 3516
rect 4580 3476 4586 3488
rect 4801 3485 4813 3488
rect 4847 3485 4859 3519
rect 4801 3479 4859 3485
rect 10318 3476 10324 3528
rect 10376 3516 10382 3528
rect 10873 3519 10931 3525
rect 10873 3516 10885 3519
rect 10376 3488 10885 3516
rect 10376 3476 10382 3488
rect 10873 3485 10885 3488
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 13832 3448 13860 3547
rect 13924 3525 13952 3624
rect 14185 3621 14197 3655
rect 14231 3621 14243 3655
rect 15838 3652 15844 3664
rect 15410 3624 15844 3652
rect 14185 3615 14243 3621
rect 15838 3612 15844 3624
rect 15896 3612 15902 3664
rect 19794 3612 19800 3664
rect 19852 3612 19858 3664
rect 20272 3661 20300 3692
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 20993 3723 21051 3729
rect 20993 3689 21005 3723
rect 21039 3720 21051 3723
rect 21174 3720 21180 3732
rect 21039 3692 21180 3720
rect 21039 3689 21051 3692
rect 20993 3683 21051 3689
rect 21174 3680 21180 3692
rect 21232 3680 21238 3732
rect 21913 3723 21971 3729
rect 21913 3689 21925 3723
rect 21959 3720 21971 3723
rect 22186 3720 22192 3732
rect 21959 3692 22192 3720
rect 21959 3689 21971 3692
rect 21913 3683 21971 3689
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 23106 3680 23112 3732
rect 23164 3680 23170 3732
rect 23382 3680 23388 3732
rect 23440 3680 23446 3732
rect 23845 3723 23903 3729
rect 23845 3689 23857 3723
rect 23891 3720 23903 3723
rect 24026 3720 24032 3732
rect 23891 3692 24032 3720
rect 23891 3689 23903 3692
rect 23845 3683 23903 3689
rect 20257 3655 20315 3661
rect 20257 3621 20269 3655
rect 20303 3621 20315 3655
rect 20257 3615 20315 3621
rect 21361 3655 21419 3661
rect 21361 3621 21373 3655
rect 21407 3652 21419 3655
rect 22097 3655 22155 3661
rect 22097 3652 22109 3655
rect 21407 3624 22109 3652
rect 21407 3621 21419 3624
rect 21361 3615 21419 3621
rect 22097 3621 22109 3624
rect 22143 3621 22155 3655
rect 22097 3615 22155 3621
rect 15470 3544 15476 3596
rect 15528 3544 15534 3596
rect 16114 3584 16120 3596
rect 15672 3556 16120 3584
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 15488 3516 15516 3544
rect 15672 3525 15700 3556
rect 16114 3544 16120 3556
rect 16172 3584 16178 3596
rect 16761 3587 16819 3593
rect 16761 3584 16773 3587
rect 16172 3556 16773 3584
rect 16172 3544 16178 3556
rect 16761 3553 16773 3556
rect 16807 3553 16819 3587
rect 16761 3547 16819 3553
rect 17034 3544 17040 3596
rect 17092 3584 17098 3596
rect 18325 3587 18383 3593
rect 18325 3584 18337 3587
rect 17092 3556 18337 3584
rect 17092 3544 17098 3556
rect 18325 3553 18337 3556
rect 18371 3553 18383 3587
rect 18325 3547 18383 3553
rect 20533 3587 20591 3593
rect 20533 3553 20545 3587
rect 20579 3584 20591 3587
rect 20898 3584 20904 3596
rect 20579 3556 20904 3584
rect 20579 3553 20591 3556
rect 20533 3547 20591 3553
rect 20898 3544 20904 3556
rect 20956 3544 20962 3596
rect 21821 3587 21879 3593
rect 21821 3553 21833 3587
rect 21867 3584 21879 3587
rect 23201 3587 23259 3593
rect 23201 3584 23213 3587
rect 21867 3556 23213 3584
rect 21867 3553 21879 3556
rect 21821 3547 21879 3553
rect 23201 3553 23213 3556
rect 23247 3584 23259 3587
rect 23400 3584 23428 3680
rect 23247 3556 23428 3584
rect 23247 3553 23259 3556
rect 23201 3547 23259 3553
rect 13909 3479 13967 3485
rect 14016 3488 15516 3516
rect 15657 3519 15715 3525
rect 14016 3448 14044 3488
rect 15657 3485 15669 3519
rect 15703 3485 15715 3519
rect 15657 3479 15715 3485
rect 16942 3476 16948 3528
rect 17000 3516 17006 3528
rect 17221 3519 17279 3525
rect 17221 3516 17233 3519
rect 17000 3488 17233 3516
rect 17000 3476 17006 3488
rect 17221 3485 17233 3488
rect 17267 3485 17279 3519
rect 17221 3479 17279 3485
rect 20254 3476 20260 3528
rect 20312 3516 20318 3528
rect 21453 3519 21511 3525
rect 21453 3516 21465 3519
rect 20312 3488 21465 3516
rect 20312 3476 20318 3488
rect 21453 3485 21465 3488
rect 21499 3485 21511 3519
rect 21453 3479 21511 3485
rect 21637 3519 21695 3525
rect 21637 3485 21649 3519
rect 21683 3485 21695 3519
rect 21637 3479 21695 3485
rect 22741 3519 22799 3525
rect 22741 3485 22753 3519
rect 22787 3516 22799 3519
rect 23474 3516 23480 3528
rect 22787 3488 23480 3516
rect 22787 3485 22799 3488
rect 22741 3479 22799 3485
rect 13832 3420 14044 3448
rect 20714 3408 20720 3460
rect 20772 3448 20778 3460
rect 20901 3451 20959 3457
rect 20901 3448 20913 3451
rect 20772 3420 20913 3448
rect 20772 3408 20778 3420
rect 20901 3417 20913 3420
rect 20947 3448 20959 3451
rect 21652 3448 21680 3479
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 23860 3448 23888 3683
rect 24026 3680 24032 3692
rect 24084 3680 24090 3732
rect 30101 3655 30159 3661
rect 30101 3621 30113 3655
rect 30147 3652 30159 3655
rect 31662 3652 31668 3664
rect 30147 3624 31668 3652
rect 30147 3621 30159 3624
rect 30101 3615 30159 3621
rect 31662 3612 31668 3624
rect 31720 3612 31726 3664
rect 25774 3544 25780 3596
rect 25832 3544 25838 3596
rect 29089 3587 29147 3593
rect 29089 3553 29101 3587
rect 29135 3584 29147 3587
rect 30006 3584 30012 3596
rect 29135 3556 30012 3584
rect 29135 3553 29147 3556
rect 29089 3547 29147 3553
rect 30006 3544 30012 3556
rect 30064 3544 30070 3596
rect 30377 3587 30435 3593
rect 30377 3584 30389 3587
rect 30116 3556 30389 3584
rect 24486 3476 24492 3528
rect 24544 3516 24550 3528
rect 24765 3519 24823 3525
rect 24765 3516 24777 3519
rect 24544 3488 24777 3516
rect 24544 3476 24550 3488
rect 24765 3485 24777 3488
rect 24811 3485 24823 3519
rect 24765 3479 24823 3485
rect 20947 3420 23888 3448
rect 20947 3417 20959 3420
rect 20901 3411 20959 3417
rect 20622 3340 20628 3392
rect 20680 3380 20686 3392
rect 30116 3380 30144 3556
rect 30377 3553 30389 3556
rect 30423 3553 30435 3587
rect 30377 3547 30435 3553
rect 30282 3476 30288 3528
rect 30340 3516 30346 3528
rect 30837 3519 30895 3525
rect 30837 3516 30849 3519
rect 30340 3488 30849 3516
rect 30340 3476 30346 3488
rect 30837 3485 30849 3488
rect 30883 3485 30895 3519
rect 30837 3479 30895 3485
rect 20680 3352 30144 3380
rect 20680 3340 20686 3352
rect 2760 3290 32200 3312
rect 2760 3238 6286 3290
rect 6338 3238 6350 3290
rect 6402 3238 6414 3290
rect 6466 3238 6478 3290
rect 6530 3238 6542 3290
rect 6594 3238 13646 3290
rect 13698 3238 13710 3290
rect 13762 3238 13774 3290
rect 13826 3238 13838 3290
rect 13890 3238 13902 3290
rect 13954 3238 21006 3290
rect 21058 3238 21070 3290
rect 21122 3238 21134 3290
rect 21186 3238 21198 3290
rect 21250 3238 21262 3290
rect 21314 3238 28366 3290
rect 28418 3238 28430 3290
rect 28482 3238 28494 3290
rect 28546 3238 28558 3290
rect 28610 3238 28622 3290
rect 28674 3238 32200 3290
rect 2760 3216 32200 3238
rect 13817 3179 13875 3185
rect 13817 3145 13829 3179
rect 13863 3176 13875 3179
rect 14182 3176 14188 3188
rect 13863 3148 14188 3176
rect 13863 3145 13875 3148
rect 13817 3139 13875 3145
rect 14182 3136 14188 3148
rect 14240 3136 14246 3188
rect 14826 3136 14832 3188
rect 14884 3136 14890 3188
rect 15010 3136 15016 3188
rect 15068 3176 15074 3188
rect 15068 3148 19472 3176
rect 15068 3136 15074 3148
rect 9677 3111 9735 3117
rect 9677 3077 9689 3111
rect 9723 3108 9735 3111
rect 14844 3108 14872 3136
rect 9723 3080 14872 3108
rect 9723 3077 9735 3080
rect 9677 3071 9735 3077
rect 15562 3068 15568 3120
rect 15620 3108 15626 3120
rect 19444 3108 19472 3148
rect 20898 3136 20904 3188
rect 20956 3176 20962 3188
rect 28997 3179 29055 3185
rect 28997 3176 29009 3179
rect 20956 3148 29009 3176
rect 20956 3136 20962 3148
rect 28997 3145 29009 3148
rect 29043 3145 29055 3179
rect 28997 3139 29055 3145
rect 29273 3179 29331 3185
rect 29273 3145 29285 3179
rect 29319 3176 29331 3179
rect 30926 3176 30932 3188
rect 29319 3148 30932 3176
rect 29319 3145 29331 3148
rect 29273 3139 29331 3145
rect 15620 3080 19380 3108
rect 19444 3080 26740 3108
rect 15620 3068 15626 3080
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 16209 3043 16267 3049
rect 16209 3009 16221 3043
rect 16255 3040 16267 3043
rect 16390 3040 16396 3052
rect 16255 3012 16396 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 16390 3000 16396 3012
rect 16448 3000 16454 3052
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3040 17739 3043
rect 18046 3040 18052 3052
rect 17727 3012 18052 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18230 3000 18236 3052
rect 18288 3040 18294 3052
rect 18601 3043 18659 3049
rect 18601 3040 18613 3043
rect 18288 3012 18613 3040
rect 18288 3000 18294 3012
rect 18601 3009 18613 3012
rect 18647 3009 18659 3043
rect 18601 3003 18659 3009
rect 19058 3000 19064 3052
rect 19116 3000 19122 3052
rect 4430 2932 4436 2984
rect 4488 2932 4494 2984
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2941 4583 2975
rect 4525 2935 4583 2941
rect 7193 2975 7251 2981
rect 7193 2941 7205 2975
rect 7239 2972 7251 2975
rect 7650 2972 7656 2984
rect 7239 2944 7656 2972
rect 7239 2941 7251 2944
rect 7193 2935 7251 2941
rect 14 2864 20 2916
rect 72 2904 78 2916
rect 3237 2907 3295 2913
rect 3237 2904 3249 2907
rect 72 2876 3249 2904
rect 72 2864 78 2876
rect 3237 2873 3249 2876
rect 3283 2873 3295 2907
rect 3237 2867 3295 2873
rect 3602 2864 3608 2916
rect 3660 2904 3666 2916
rect 4540 2904 4568 2935
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 9214 2932 9220 2984
rect 9272 2932 9278 2984
rect 9493 2975 9551 2981
rect 9493 2941 9505 2975
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 3660 2876 4568 2904
rect 3660 2864 3666 2876
rect 5810 2864 5816 2916
rect 5868 2904 5874 2916
rect 6089 2907 6147 2913
rect 6089 2904 6101 2907
rect 5868 2876 6101 2904
rect 5868 2864 5874 2876
rect 6089 2873 6101 2876
rect 6135 2873 6147 2907
rect 6089 2867 6147 2873
rect 7282 2864 7288 2916
rect 7340 2904 7346 2916
rect 8205 2907 8263 2913
rect 8205 2904 8217 2907
rect 7340 2876 8217 2904
rect 7340 2864 7346 2876
rect 8205 2873 8217 2876
rect 8251 2873 8263 2907
rect 8205 2867 8263 2873
rect 9030 2864 9036 2916
rect 9088 2904 9094 2916
rect 9508 2904 9536 2935
rect 11514 2932 11520 2984
rect 11572 2972 11578 2984
rect 11609 2975 11667 2981
rect 11609 2972 11621 2975
rect 11572 2944 11621 2972
rect 11572 2932 11578 2944
rect 11609 2941 11621 2944
rect 11655 2941 11667 2975
rect 11609 2935 11667 2941
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 15378 2932 15384 2984
rect 15436 2972 15442 2984
rect 15565 2975 15623 2981
rect 15565 2972 15577 2975
rect 15436 2944 15577 2972
rect 15436 2932 15442 2944
rect 15565 2941 15577 2944
rect 15611 2972 15623 2975
rect 16298 2972 16304 2984
rect 15611 2944 16304 2972
rect 15611 2941 15623 2944
rect 15565 2935 15623 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 17954 2932 17960 2984
rect 18012 2932 18018 2984
rect 19352 2981 19380 3080
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19484 3012 19809 3040
rect 19484 3000 19490 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 23937 3043 23995 3049
rect 23937 3040 23949 3043
rect 22612 3012 23949 3040
rect 22612 3000 22618 3012
rect 23937 3009 23949 3012
rect 23983 3009 23995 3043
rect 23937 3003 23995 3009
rect 25774 3000 25780 3052
rect 25832 3040 25838 3052
rect 26513 3043 26571 3049
rect 26513 3040 26525 3043
rect 25832 3012 26525 3040
rect 25832 3000 25838 3012
rect 26513 3009 26525 3012
rect 26559 3009 26571 3043
rect 26513 3003 26571 3009
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 21266 2932 21272 2984
rect 21324 2972 21330 2984
rect 21545 2975 21603 2981
rect 21545 2972 21557 2975
rect 21324 2944 21557 2972
rect 21324 2932 21330 2944
rect 21545 2941 21557 2944
rect 21591 2941 21603 2975
rect 21545 2935 21603 2941
rect 23474 2932 23480 2984
rect 23532 2932 23538 2984
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 26053 2975 26111 2981
rect 26053 2972 26065 2975
rect 23624 2944 26065 2972
rect 23624 2932 23630 2944
rect 26053 2941 26065 2944
rect 26099 2941 26111 2975
rect 26053 2935 26111 2941
rect 18138 2904 18144 2916
rect 9088 2876 9536 2904
rect 9600 2876 18144 2904
rect 9088 2864 9094 2876
rect 4709 2839 4767 2845
rect 4709 2805 4721 2839
rect 4755 2836 4767 2839
rect 9600 2836 9628 2876
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 18322 2864 18328 2916
rect 18380 2904 18386 2916
rect 26712 2904 26740 3080
rect 29012 3040 29040 3139
rect 30926 3136 30932 3148
rect 30984 3136 30990 3188
rect 31665 3179 31723 3185
rect 31665 3145 31677 3179
rect 31711 3176 31723 3179
rect 31846 3176 31852 3188
rect 31711 3148 31852 3176
rect 31711 3145 31723 3148
rect 31665 3139 31723 3145
rect 31846 3136 31852 3148
rect 31904 3136 31910 3188
rect 30837 3043 30895 3049
rect 29012 3012 29684 3040
rect 27062 2932 27068 2984
rect 27120 2972 27126 2984
rect 27709 2975 27767 2981
rect 27709 2972 27721 2975
rect 27120 2944 27721 2972
rect 27120 2932 27126 2944
rect 27709 2941 27721 2944
rect 27755 2941 27767 2975
rect 27709 2935 27767 2941
rect 29089 2975 29147 2981
rect 29089 2941 29101 2975
rect 29135 2972 29147 2975
rect 29362 2972 29368 2984
rect 29135 2944 29368 2972
rect 29135 2941 29147 2944
rect 29089 2935 29147 2941
rect 29362 2932 29368 2944
rect 29420 2932 29426 2984
rect 29656 2981 29684 3012
rect 30837 3009 30849 3043
rect 30883 3040 30895 3043
rect 32214 3040 32220 3052
rect 30883 3012 32220 3040
rect 30883 3009 30895 3012
rect 30837 3003 30895 3009
rect 32214 3000 32220 3012
rect 32272 3000 32278 3052
rect 29641 2975 29699 2981
rect 29641 2941 29653 2975
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 31573 2975 31631 2981
rect 31573 2941 31585 2975
rect 31619 2972 31631 2975
rect 31849 2975 31907 2981
rect 31619 2944 31754 2972
rect 31619 2941 31631 2944
rect 31573 2935 31631 2941
rect 18380 2876 22094 2904
rect 26712 2876 31432 2904
rect 18380 2864 18386 2876
rect 4755 2808 9628 2836
rect 16669 2839 16727 2845
rect 4755 2805 4767 2808
rect 4709 2799 4767 2805
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 18690 2836 18696 2848
rect 16715 2808 18696 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 19702 2796 19708 2848
rect 19760 2836 19766 2848
rect 21361 2839 21419 2845
rect 21361 2836 21373 2839
rect 19760 2808 21373 2836
rect 19760 2796 19766 2808
rect 21361 2805 21373 2808
rect 21407 2805 21419 2839
rect 22066 2836 22094 2876
rect 31404 2845 31432 2876
rect 27525 2839 27583 2845
rect 27525 2836 27537 2839
rect 22066 2808 27537 2836
rect 21361 2799 21419 2805
rect 27525 2805 27537 2808
rect 27571 2805 27583 2839
rect 27525 2799 27583 2805
rect 31389 2839 31447 2845
rect 31389 2805 31401 2839
rect 31435 2805 31447 2839
rect 31726 2836 31754 2944
rect 31849 2941 31861 2975
rect 31895 2941 31907 2975
rect 31849 2935 31907 2941
rect 31864 2904 31892 2935
rect 33134 2904 33140 2916
rect 31864 2876 33140 2904
rect 33134 2864 33140 2876
rect 33192 2864 33198 2916
rect 34790 2836 34796 2848
rect 31726 2808 34796 2836
rect 31389 2799 31447 2805
rect 34790 2796 34796 2808
rect 34848 2796 34854 2848
rect 2760 2746 32200 2768
rect 2760 2694 6946 2746
rect 6998 2694 7010 2746
rect 7062 2694 7074 2746
rect 7126 2694 7138 2746
rect 7190 2694 7202 2746
rect 7254 2694 14306 2746
rect 14358 2694 14370 2746
rect 14422 2694 14434 2746
rect 14486 2694 14498 2746
rect 14550 2694 14562 2746
rect 14614 2694 21666 2746
rect 21718 2694 21730 2746
rect 21782 2694 21794 2746
rect 21846 2694 21858 2746
rect 21910 2694 21922 2746
rect 21974 2694 29026 2746
rect 29078 2694 29090 2746
rect 29142 2694 29154 2746
rect 29206 2694 29218 2746
rect 29270 2694 29282 2746
rect 29334 2694 32200 2746
rect 2760 2672 32200 2694
<< via1 >>
rect 21456 32308 21508 32360
rect 17776 32240 17828 32292
rect 25964 32240 26016 32292
rect 25780 32172 25832 32224
rect 28264 32172 28316 32224
rect 28632 32172 28684 32224
rect 6946 32070 6998 32122
rect 7010 32070 7062 32122
rect 7074 32070 7126 32122
rect 7138 32070 7190 32122
rect 7202 32070 7254 32122
rect 14306 32070 14358 32122
rect 14370 32070 14422 32122
rect 14434 32070 14486 32122
rect 14498 32070 14550 32122
rect 14562 32070 14614 32122
rect 21666 32070 21718 32122
rect 21730 32070 21782 32122
rect 21794 32070 21846 32122
rect 21858 32070 21910 32122
rect 21922 32070 21974 32122
rect 29026 32070 29078 32122
rect 29090 32070 29142 32122
rect 29154 32070 29206 32122
rect 29218 32070 29270 32122
rect 29282 32070 29334 32122
rect 7564 31968 7616 32020
rect 9680 31968 9732 32020
rect 1032 31900 1084 31952
rect 4160 31900 4212 31952
rect 5172 31900 5224 31952
rect 6460 31900 6512 31952
rect 3884 31875 3936 31884
rect 3884 31841 3893 31875
rect 3893 31841 3927 31875
rect 3927 31841 3936 31875
rect 3884 31832 3936 31841
rect 6644 31875 6696 31884
rect 6644 31841 6653 31875
rect 6653 31841 6687 31875
rect 6687 31841 6696 31875
rect 6644 31832 6696 31841
rect 8668 31943 8720 31952
rect 8668 31909 8677 31943
rect 8677 31909 8711 31943
rect 8711 31909 8720 31943
rect 8668 31900 8720 31909
rect 11612 31968 11664 32020
rect 9680 31875 9732 31884
rect 9680 31841 9689 31875
rect 9689 31841 9723 31875
rect 9723 31841 9732 31875
rect 9680 31832 9732 31841
rect 12348 31832 12400 31884
rect 14372 31943 14424 31952
rect 14372 31909 14381 31943
rect 14381 31909 14415 31943
rect 14415 31909 14424 31943
rect 14372 31900 14424 31909
rect 16120 31900 16172 31952
rect 15384 31875 15436 31884
rect 15384 31841 15393 31875
rect 15393 31841 15427 31875
rect 15427 31841 15436 31875
rect 15384 31832 15436 31841
rect 16580 31832 16632 31884
rect 14096 31807 14148 31816
rect 14096 31773 14105 31807
rect 14105 31773 14139 31807
rect 14139 31773 14148 31807
rect 14096 31764 14148 31773
rect 17408 31968 17460 32020
rect 17868 32011 17920 32020
rect 17868 31977 17877 32011
rect 17877 31977 17911 32011
rect 17911 31977 17920 32011
rect 17868 31968 17920 31977
rect 18696 31968 18748 32020
rect 18788 32011 18840 32020
rect 18788 31977 18797 32011
rect 18797 31977 18831 32011
rect 18831 31977 18840 32011
rect 18788 31968 18840 31977
rect 18972 31968 19024 32020
rect 20628 31900 20680 31952
rect 22008 31968 22060 32020
rect 25780 31968 25832 32020
rect 31024 31968 31076 32020
rect 33140 31968 33192 32020
rect 23848 31900 23900 31952
rect 24032 31875 24084 31884
rect 24032 31841 24041 31875
rect 24041 31841 24075 31875
rect 24075 31841 24084 31875
rect 24032 31832 24084 31841
rect 25136 31900 25188 31952
rect 25504 31875 25556 31884
rect 25504 31841 25513 31875
rect 25513 31841 25547 31875
rect 25547 31841 25556 31875
rect 25504 31832 25556 31841
rect 26424 31900 26476 31952
rect 25964 31764 26016 31816
rect 28080 31900 28132 31952
rect 28632 31875 28684 31884
rect 28632 31841 28641 31875
rect 28641 31841 28675 31875
rect 28675 31841 28684 31875
rect 28632 31832 28684 31841
rect 28724 31832 28776 31884
rect 28356 31764 28408 31816
rect 19524 31696 19576 31748
rect 11888 31628 11940 31680
rect 18420 31628 18472 31680
rect 22376 31671 22428 31680
rect 22376 31637 22385 31671
rect 22385 31637 22419 31671
rect 22419 31637 22428 31671
rect 22376 31628 22428 31637
rect 25964 31628 26016 31680
rect 6286 31526 6338 31578
rect 6350 31526 6402 31578
rect 6414 31526 6466 31578
rect 6478 31526 6530 31578
rect 6542 31526 6594 31578
rect 13646 31526 13698 31578
rect 13710 31526 13762 31578
rect 13774 31526 13826 31578
rect 13838 31526 13890 31578
rect 13902 31526 13954 31578
rect 21006 31526 21058 31578
rect 21070 31526 21122 31578
rect 21134 31526 21186 31578
rect 21198 31526 21250 31578
rect 21262 31526 21314 31578
rect 28366 31526 28418 31578
rect 28430 31526 28482 31578
rect 28494 31526 28546 31578
rect 28558 31526 28610 31578
rect 28622 31526 28674 31578
rect 15016 31424 15068 31476
rect 2320 31288 2372 31340
rect 23664 31356 23716 31408
rect 24584 31356 24636 31408
rect 24952 31356 25004 31408
rect 4160 31220 4212 31272
rect 12900 31288 12952 31340
rect 14188 31288 14240 31340
rect 14556 31331 14608 31340
rect 14556 31297 14565 31331
rect 14565 31297 14599 31331
rect 14599 31297 14608 31331
rect 14556 31288 14608 31297
rect 12440 31220 12492 31272
rect 16580 31263 16632 31272
rect 16580 31229 16589 31263
rect 16589 31229 16623 31263
rect 16623 31229 16632 31263
rect 16580 31220 16632 31229
rect 18052 31263 18104 31272
rect 18052 31229 18061 31263
rect 18061 31229 18095 31263
rect 18095 31229 18104 31263
rect 18052 31220 18104 31229
rect 22100 31220 22152 31272
rect 23112 31220 23164 31272
rect 24492 31288 24544 31340
rect 23756 31263 23808 31272
rect 23756 31229 23765 31263
rect 23765 31229 23799 31263
rect 23799 31229 23808 31263
rect 23756 31220 23808 31229
rect 24032 31220 24084 31272
rect 24584 31263 24636 31272
rect 24584 31229 24593 31263
rect 24593 31229 24627 31263
rect 24627 31229 24636 31263
rect 24584 31220 24636 31229
rect 24676 31220 24728 31272
rect 25872 31356 25924 31408
rect 26332 31356 26384 31408
rect 25136 31220 25188 31272
rect 24308 31195 24360 31204
rect 24308 31161 24325 31195
rect 24325 31161 24360 31195
rect 24308 31152 24360 31161
rect 24400 31195 24452 31204
rect 24400 31161 24409 31195
rect 24409 31161 24443 31195
rect 24443 31161 24452 31195
rect 24400 31152 24452 31161
rect 24492 31195 24544 31204
rect 24492 31161 24501 31195
rect 24501 31161 24535 31195
rect 24535 31161 24544 31195
rect 24492 31152 24544 31161
rect 10784 31127 10836 31136
rect 10784 31093 10793 31127
rect 10793 31093 10827 31127
rect 10827 31093 10836 31127
rect 10784 31084 10836 31093
rect 11336 31084 11388 31136
rect 11796 31127 11848 31136
rect 11796 31093 11805 31127
rect 11805 31093 11839 31127
rect 11839 31093 11848 31127
rect 11796 31084 11848 31093
rect 15108 31127 15160 31136
rect 15108 31093 15117 31127
rect 15117 31093 15151 31127
rect 15151 31093 15160 31127
rect 15108 31084 15160 31093
rect 15292 31127 15344 31136
rect 15292 31093 15301 31127
rect 15301 31093 15335 31127
rect 15335 31093 15344 31127
rect 15292 31084 15344 31093
rect 15936 31084 15988 31136
rect 16028 31127 16080 31136
rect 16028 31093 16037 31127
rect 16037 31093 16071 31127
rect 16071 31093 16080 31127
rect 16028 31084 16080 31093
rect 17500 31127 17552 31136
rect 17500 31093 17509 31127
rect 17509 31093 17543 31127
rect 17543 31093 17552 31127
rect 17500 31084 17552 31093
rect 18604 31084 18656 31136
rect 21364 31127 21416 31136
rect 21364 31093 21373 31127
rect 21373 31093 21407 31127
rect 21407 31093 21416 31127
rect 21364 31084 21416 31093
rect 23664 31084 23716 31136
rect 23940 31127 23992 31136
rect 23940 31093 23949 31127
rect 23949 31093 23983 31127
rect 23983 31093 23992 31127
rect 23940 31084 23992 31093
rect 24768 31127 24820 31136
rect 24768 31093 24777 31127
rect 24777 31093 24811 31127
rect 24811 31093 24820 31127
rect 24768 31084 24820 31093
rect 25228 31084 25280 31136
rect 25320 31084 25372 31136
rect 25688 31263 25740 31272
rect 25688 31229 25697 31263
rect 25697 31229 25731 31263
rect 25731 31229 25740 31263
rect 25688 31220 25740 31229
rect 26056 31331 26108 31340
rect 26056 31297 26065 31331
rect 26065 31297 26099 31331
rect 26099 31297 26108 31331
rect 26056 31288 26108 31297
rect 26332 31263 26384 31272
rect 26332 31229 26341 31263
rect 26341 31229 26375 31263
rect 26375 31229 26384 31263
rect 26332 31220 26384 31229
rect 26424 31263 26476 31272
rect 26424 31229 26433 31263
rect 26433 31229 26467 31263
rect 26467 31229 26476 31263
rect 26424 31220 26476 31229
rect 25596 31195 25648 31204
rect 25596 31161 25605 31195
rect 25605 31161 25639 31195
rect 25639 31161 25648 31195
rect 25596 31152 25648 31161
rect 26884 31263 26936 31272
rect 26884 31229 26893 31263
rect 26893 31229 26927 31263
rect 26927 31229 26936 31263
rect 26884 31220 26936 31229
rect 30104 31331 30156 31340
rect 30104 31297 30113 31331
rect 30113 31297 30147 31331
rect 30147 31297 30156 31331
rect 30104 31288 30156 31297
rect 34152 31288 34204 31340
rect 29644 31263 29696 31272
rect 29644 31229 29653 31263
rect 29653 31229 29687 31263
rect 29687 31229 29696 31263
rect 29644 31220 29696 31229
rect 25780 31084 25832 31136
rect 26516 31084 26568 31136
rect 26608 31084 26660 31136
rect 27160 31084 27212 31136
rect 6946 30982 6998 31034
rect 7010 30982 7062 31034
rect 7074 30982 7126 31034
rect 7138 30982 7190 31034
rect 7202 30982 7254 31034
rect 14306 30982 14358 31034
rect 14370 30982 14422 31034
rect 14434 30982 14486 31034
rect 14498 30982 14550 31034
rect 14562 30982 14614 31034
rect 21666 30982 21718 31034
rect 21730 30982 21782 31034
rect 21794 30982 21846 31034
rect 21858 30982 21910 31034
rect 21922 30982 21974 31034
rect 29026 30982 29078 31034
rect 29090 30982 29142 31034
rect 29154 30982 29206 31034
rect 29218 30982 29270 31034
rect 29282 30982 29334 31034
rect 11796 30880 11848 30932
rect 11888 30880 11940 30932
rect 15292 30812 15344 30864
rect 16028 30812 16080 30864
rect 16948 30812 17000 30864
rect 4436 30787 4488 30796
rect 4436 30753 4445 30787
rect 4445 30753 4479 30787
rect 4479 30753 4488 30787
rect 4436 30744 4488 30753
rect 4528 30787 4580 30796
rect 4528 30753 4537 30787
rect 4537 30753 4571 30787
rect 4571 30753 4580 30787
rect 4528 30744 4580 30753
rect 1308 30676 1360 30728
rect 5356 30676 5408 30728
rect 10876 30676 10928 30728
rect 12440 30744 12492 30796
rect 12624 30787 12676 30796
rect 12624 30753 12633 30787
rect 12633 30753 12667 30787
rect 12667 30753 12676 30787
rect 12624 30744 12676 30753
rect 12900 30583 12952 30592
rect 12900 30549 12909 30583
rect 12909 30549 12943 30583
rect 12943 30549 12952 30583
rect 12900 30540 12952 30549
rect 13544 30719 13596 30728
rect 13544 30685 13553 30719
rect 13553 30685 13587 30719
rect 13587 30685 13596 30719
rect 13544 30676 13596 30685
rect 14280 30540 14332 30592
rect 15016 30651 15068 30660
rect 15016 30617 15025 30651
rect 15025 30617 15059 30651
rect 15059 30617 15068 30651
rect 15016 30608 15068 30617
rect 18420 30719 18472 30728
rect 18420 30685 18429 30719
rect 18429 30685 18463 30719
rect 18463 30685 18472 30719
rect 18420 30676 18472 30685
rect 22376 30880 22428 30932
rect 23756 30880 23808 30932
rect 24584 30880 24636 30932
rect 24952 30880 25004 30932
rect 25136 30880 25188 30932
rect 25688 30880 25740 30932
rect 26424 30923 26476 30932
rect 26424 30889 26433 30923
rect 26433 30889 26467 30923
rect 26467 30889 26476 30923
rect 26424 30880 26476 30889
rect 21364 30812 21416 30864
rect 24308 30812 24360 30864
rect 24676 30812 24728 30864
rect 25044 30812 25096 30864
rect 19524 30744 19576 30796
rect 23848 30787 23900 30796
rect 23848 30753 23857 30787
rect 23857 30753 23891 30787
rect 23891 30753 23900 30787
rect 23848 30744 23900 30753
rect 24032 30744 24084 30796
rect 24768 30744 24820 30796
rect 25320 30787 25372 30796
rect 25320 30753 25329 30787
rect 25329 30753 25363 30787
rect 25363 30753 25372 30787
rect 25320 30744 25372 30753
rect 17316 30608 17368 30660
rect 17776 30608 17828 30660
rect 18788 30608 18840 30660
rect 15200 30540 15252 30592
rect 17040 30540 17092 30592
rect 18604 30540 18656 30592
rect 20352 30719 20404 30728
rect 20352 30685 20361 30719
rect 20361 30685 20395 30719
rect 20395 30685 20404 30719
rect 20352 30676 20404 30685
rect 20720 30676 20772 30728
rect 22928 30719 22980 30728
rect 22928 30685 22937 30719
rect 22937 30685 22971 30719
rect 22971 30685 22980 30719
rect 22928 30676 22980 30685
rect 25228 30676 25280 30728
rect 26240 30855 26292 30864
rect 26240 30821 26247 30855
rect 26247 30821 26281 30855
rect 26281 30821 26292 30855
rect 26240 30812 26292 30821
rect 25872 30744 25924 30796
rect 27620 30880 27672 30932
rect 28172 30880 28224 30932
rect 28724 30880 28776 30932
rect 32588 30880 32640 30932
rect 28264 30744 28316 30796
rect 28816 30787 28868 30796
rect 28816 30753 28825 30787
rect 28825 30753 28859 30787
rect 28859 30753 28868 30787
rect 28816 30744 28868 30753
rect 29828 30744 29880 30796
rect 31576 30855 31628 30864
rect 31576 30821 31585 30855
rect 31585 30821 31619 30855
rect 31619 30821 31628 30855
rect 31576 30812 31628 30821
rect 30380 30744 30432 30796
rect 26424 30608 26476 30660
rect 20260 30583 20312 30592
rect 20260 30549 20269 30583
rect 20269 30549 20303 30583
rect 20303 30549 20312 30583
rect 20260 30540 20312 30549
rect 22284 30583 22336 30592
rect 22284 30549 22293 30583
rect 22293 30549 22327 30583
rect 22327 30549 22336 30583
rect 22284 30540 22336 30549
rect 24584 30583 24636 30592
rect 24584 30549 24593 30583
rect 24593 30549 24627 30583
rect 24627 30549 24636 30583
rect 24584 30540 24636 30549
rect 26240 30540 26292 30592
rect 26792 30719 26844 30728
rect 26792 30685 26801 30719
rect 26801 30685 26835 30719
rect 26835 30685 26844 30719
rect 26792 30676 26844 30685
rect 29736 30676 29788 30728
rect 28724 30583 28776 30592
rect 28724 30549 28733 30583
rect 28733 30549 28767 30583
rect 28767 30549 28776 30583
rect 28724 30540 28776 30549
rect 6286 30438 6338 30490
rect 6350 30438 6402 30490
rect 6414 30438 6466 30490
rect 6478 30438 6530 30490
rect 6542 30438 6594 30490
rect 13646 30438 13698 30490
rect 13710 30438 13762 30490
rect 13774 30438 13826 30490
rect 13838 30438 13890 30490
rect 13902 30438 13954 30490
rect 21006 30438 21058 30490
rect 21070 30438 21122 30490
rect 21134 30438 21186 30490
rect 21198 30438 21250 30490
rect 21262 30438 21314 30490
rect 28366 30438 28418 30490
rect 28430 30438 28482 30490
rect 28494 30438 28546 30490
rect 28558 30438 28610 30490
rect 28622 30438 28674 30490
rect 12348 30311 12400 30320
rect 12348 30277 12357 30311
rect 12357 30277 12391 30311
rect 12391 30277 12400 30311
rect 12348 30268 12400 30277
rect 2780 30200 2832 30252
rect 9680 30243 9732 30252
rect 9680 30209 9689 30243
rect 9689 30209 9723 30243
rect 9723 30209 9732 30243
rect 9680 30200 9732 30209
rect 10876 30200 10928 30252
rect 14188 30200 14240 30252
rect 14280 30200 14332 30252
rect 4528 30132 4580 30184
rect 11980 30132 12032 30184
rect 10324 30064 10376 30116
rect 12900 30064 12952 30116
rect 16580 30336 16632 30388
rect 16948 30379 17000 30388
rect 16948 30345 16957 30379
rect 16957 30345 16991 30379
rect 16991 30345 17000 30379
rect 16948 30336 17000 30345
rect 17316 30336 17368 30388
rect 20720 30336 20772 30388
rect 14740 30200 14792 30252
rect 15200 30243 15252 30252
rect 15200 30209 15209 30243
rect 15209 30209 15243 30243
rect 15243 30209 15252 30243
rect 15200 30200 15252 30209
rect 18972 30311 19024 30320
rect 18972 30277 18981 30311
rect 18981 30277 19015 30311
rect 19015 30277 19024 30311
rect 18972 30268 19024 30277
rect 15108 30132 15160 30184
rect 17500 30243 17552 30252
rect 17500 30209 17509 30243
rect 17509 30209 17543 30243
rect 17543 30209 17552 30243
rect 17500 30200 17552 30209
rect 16304 30064 16356 30116
rect 7656 29996 7708 30048
rect 8300 30039 8352 30048
rect 8300 30005 8309 30039
rect 8309 30005 8343 30039
rect 8343 30005 8352 30039
rect 8300 29996 8352 30005
rect 8760 29996 8812 30048
rect 11888 29996 11940 30048
rect 15936 29996 15988 30048
rect 17040 30132 17092 30184
rect 19340 30200 19392 30252
rect 22100 30336 22152 30388
rect 22560 30336 22612 30388
rect 23848 30336 23900 30388
rect 23940 30336 23992 30388
rect 24400 30336 24452 30388
rect 24952 30336 25004 30388
rect 25320 30379 25372 30388
rect 25320 30345 25329 30379
rect 25329 30345 25363 30379
rect 25363 30345 25372 30379
rect 25320 30336 25372 30345
rect 26884 30336 26936 30388
rect 27528 30336 27580 30388
rect 28816 30336 28868 30388
rect 20260 30175 20312 30184
rect 20260 30141 20269 30175
rect 20269 30141 20303 30175
rect 20303 30141 20312 30175
rect 20260 30132 20312 30141
rect 22100 30200 22152 30252
rect 23480 30200 23532 30252
rect 24584 30200 24636 30252
rect 25228 30200 25280 30252
rect 21548 30132 21600 30184
rect 25504 30132 25556 30184
rect 25872 30175 25924 30184
rect 25872 30141 25881 30175
rect 25881 30141 25915 30175
rect 25915 30141 25924 30175
rect 27068 30200 27120 30252
rect 27160 30200 27212 30252
rect 30380 30336 30432 30388
rect 25872 30132 25924 30141
rect 27896 30175 27948 30184
rect 27896 30141 27905 30175
rect 27905 30141 27939 30175
rect 27939 30141 27948 30175
rect 27896 30132 27948 30141
rect 28264 30132 28316 30184
rect 28908 30132 28960 30184
rect 29920 30175 29972 30184
rect 29920 30141 29929 30175
rect 29929 30141 29963 30175
rect 29963 30141 29972 30175
rect 29920 30132 29972 30141
rect 30012 30132 30064 30184
rect 30656 30175 30708 30184
rect 30656 30141 30665 30175
rect 30665 30141 30699 30175
rect 30699 30141 30708 30175
rect 30656 30132 30708 30141
rect 30932 30132 30984 30184
rect 33048 30200 33100 30252
rect 19708 30039 19760 30048
rect 19708 30005 19717 30039
rect 19717 30005 19751 30039
rect 19751 30005 19760 30039
rect 19708 29996 19760 30005
rect 19892 29996 19944 30048
rect 20444 29996 20496 30048
rect 22008 30107 22060 30116
rect 22008 30073 22017 30107
rect 22017 30073 22051 30107
rect 22051 30073 22060 30107
rect 22008 30064 22060 30073
rect 22744 30064 22796 30116
rect 25964 30064 26016 30116
rect 28356 30064 28408 30116
rect 22284 29996 22336 30048
rect 22928 29996 22980 30048
rect 27160 29996 27212 30048
rect 27252 29996 27304 30048
rect 29368 30039 29420 30048
rect 29368 30005 29377 30039
rect 29377 30005 29411 30039
rect 29411 30005 29420 30039
rect 29368 29996 29420 30005
rect 29552 29996 29604 30048
rect 31300 30039 31352 30048
rect 31300 30005 31309 30039
rect 31309 30005 31343 30039
rect 31343 30005 31352 30039
rect 31300 29996 31352 30005
rect 31484 29996 31536 30048
rect 6946 29894 6998 29946
rect 7010 29894 7062 29946
rect 7074 29894 7126 29946
rect 7138 29894 7190 29946
rect 7202 29894 7254 29946
rect 14306 29894 14358 29946
rect 14370 29894 14422 29946
rect 14434 29894 14486 29946
rect 14498 29894 14550 29946
rect 14562 29894 14614 29946
rect 21666 29894 21718 29946
rect 21730 29894 21782 29946
rect 21794 29894 21846 29946
rect 21858 29894 21910 29946
rect 21922 29894 21974 29946
rect 29026 29894 29078 29946
rect 29090 29894 29142 29946
rect 29154 29894 29206 29946
rect 29218 29894 29270 29946
rect 29282 29894 29334 29946
rect 4436 29792 4488 29844
rect 9680 29792 9732 29844
rect 10324 29835 10376 29844
rect 10324 29801 10333 29835
rect 10333 29801 10367 29835
rect 10367 29801 10376 29835
rect 10324 29792 10376 29801
rect 11980 29835 12032 29844
rect 11980 29801 11989 29835
rect 11989 29801 12023 29835
rect 12023 29801 12032 29835
rect 11980 29792 12032 29801
rect 12348 29792 12400 29844
rect 13544 29792 13596 29844
rect 15016 29792 15068 29844
rect 15200 29792 15252 29844
rect 8300 29724 8352 29776
rect 3148 29699 3200 29708
rect 3148 29665 3157 29699
rect 3157 29665 3191 29699
rect 3191 29665 3200 29699
rect 3148 29656 3200 29665
rect 3516 29631 3568 29640
rect 3516 29597 3525 29631
rect 3525 29597 3559 29631
rect 3559 29597 3568 29631
rect 3516 29588 3568 29597
rect 15108 29724 15160 29776
rect 18052 29792 18104 29844
rect 18972 29792 19024 29844
rect 7380 29588 7432 29640
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 8300 29588 8352 29597
rect 11244 29588 11296 29640
rect 11612 29631 11664 29640
rect 11612 29597 11621 29631
rect 11621 29597 11655 29631
rect 11655 29597 11664 29631
rect 11612 29588 11664 29597
rect 12072 29520 12124 29572
rect 14832 29656 14884 29708
rect 16304 29656 16356 29708
rect 13636 29588 13688 29640
rect 14096 29631 14148 29640
rect 14096 29597 14105 29631
rect 14105 29597 14139 29631
rect 14139 29597 14148 29631
rect 14096 29588 14148 29597
rect 14740 29588 14792 29640
rect 15752 29631 15804 29640
rect 15752 29597 15761 29631
rect 15761 29597 15795 29631
rect 15795 29597 15804 29631
rect 15752 29588 15804 29597
rect 19340 29724 19392 29776
rect 16580 29631 16632 29640
rect 16580 29597 16589 29631
rect 16589 29597 16623 29631
rect 16623 29597 16632 29631
rect 16580 29588 16632 29597
rect 18512 29656 18564 29708
rect 20352 29792 20404 29844
rect 20720 29792 20772 29844
rect 21456 29792 21508 29844
rect 22008 29792 22060 29844
rect 22744 29835 22796 29844
rect 22744 29801 22753 29835
rect 22753 29801 22787 29835
rect 22787 29801 22796 29835
rect 22744 29792 22796 29801
rect 23756 29792 23808 29844
rect 24492 29792 24544 29844
rect 24768 29792 24820 29844
rect 25688 29792 25740 29844
rect 26332 29792 26384 29844
rect 27896 29792 27948 29844
rect 19708 29767 19760 29776
rect 19708 29733 19717 29767
rect 19717 29733 19751 29767
rect 19751 29733 19760 29767
rect 19708 29724 19760 29733
rect 20444 29724 20496 29776
rect 22560 29656 22612 29708
rect 23112 29656 23164 29708
rect 13452 29495 13504 29504
rect 13452 29461 13461 29495
rect 13461 29461 13495 29495
rect 13495 29461 13504 29495
rect 17776 29588 17828 29640
rect 18696 29588 18748 29640
rect 23664 29588 23716 29640
rect 24400 29699 24452 29708
rect 24400 29665 24409 29699
rect 24409 29665 24443 29699
rect 24443 29665 24452 29699
rect 24400 29656 24452 29665
rect 24676 29699 24728 29708
rect 24676 29665 24711 29699
rect 24711 29665 24728 29699
rect 24676 29656 24728 29665
rect 25228 29699 25280 29708
rect 25228 29665 25237 29699
rect 25237 29665 25271 29699
rect 25271 29665 25280 29699
rect 25228 29656 25280 29665
rect 26056 29724 26108 29776
rect 28724 29724 28776 29776
rect 29000 29835 29052 29844
rect 29000 29801 29009 29835
rect 29009 29801 29043 29835
rect 29043 29801 29052 29835
rect 29000 29792 29052 29801
rect 29276 29792 29328 29844
rect 29736 29792 29788 29844
rect 29920 29792 29972 29844
rect 30196 29835 30248 29844
rect 30196 29801 30205 29835
rect 30205 29801 30239 29835
rect 30239 29801 30248 29835
rect 30196 29792 30248 29801
rect 31668 29767 31720 29776
rect 31668 29733 31677 29767
rect 31677 29733 31711 29767
rect 31711 29733 31720 29767
rect 31668 29724 31720 29733
rect 29184 29656 29236 29708
rect 30380 29656 30432 29708
rect 24768 29520 24820 29572
rect 13452 29452 13504 29461
rect 14372 29495 14424 29504
rect 14372 29461 14381 29495
rect 14381 29461 14415 29495
rect 14415 29461 14424 29495
rect 14372 29452 14424 29461
rect 16856 29452 16908 29504
rect 18328 29495 18380 29504
rect 18328 29461 18337 29495
rect 18337 29461 18371 29495
rect 18371 29461 18380 29495
rect 18328 29452 18380 29461
rect 19156 29495 19208 29504
rect 19156 29461 19165 29495
rect 19165 29461 19199 29495
rect 19199 29461 19208 29495
rect 19156 29452 19208 29461
rect 21548 29495 21600 29504
rect 21548 29461 21557 29495
rect 21557 29461 21591 29495
rect 21591 29461 21600 29495
rect 21548 29452 21600 29461
rect 23756 29452 23808 29504
rect 24952 29452 25004 29504
rect 27988 29588 28040 29640
rect 28356 29631 28408 29640
rect 28356 29597 28365 29631
rect 28365 29597 28399 29631
rect 28399 29597 28408 29631
rect 28356 29588 28408 29597
rect 27160 29520 27212 29572
rect 26148 29452 26200 29504
rect 26240 29452 26292 29504
rect 29276 29452 29328 29504
rect 29552 29452 29604 29504
rect 31392 29452 31444 29504
rect 6286 29350 6338 29402
rect 6350 29350 6402 29402
rect 6414 29350 6466 29402
rect 6478 29350 6530 29402
rect 6542 29350 6594 29402
rect 13646 29350 13698 29402
rect 13710 29350 13762 29402
rect 13774 29350 13826 29402
rect 13838 29350 13890 29402
rect 13902 29350 13954 29402
rect 21006 29350 21058 29402
rect 21070 29350 21122 29402
rect 21134 29350 21186 29402
rect 21198 29350 21250 29402
rect 21262 29350 21314 29402
rect 28366 29350 28418 29402
rect 28430 29350 28482 29402
rect 28494 29350 28546 29402
rect 28558 29350 28610 29402
rect 28622 29350 28674 29402
rect 3884 29248 3936 29300
rect 8300 29248 8352 29300
rect 14372 29248 14424 29300
rect 18328 29248 18380 29300
rect 20260 29248 20312 29300
rect 8392 29180 8444 29232
rect 4988 29019 5040 29028
rect 4988 28985 4997 29019
rect 4997 28985 5031 29019
rect 5031 28985 5040 29019
rect 4988 28976 5040 28985
rect 4252 28908 4304 28960
rect 7656 29087 7708 29096
rect 7656 29053 7665 29087
rect 7665 29053 7699 29087
rect 7699 29053 7708 29087
rect 7656 29044 7708 29053
rect 6184 28976 6236 29028
rect 6828 28908 6880 28960
rect 10784 29112 10836 29164
rect 11612 29180 11664 29232
rect 11152 29112 11204 29164
rect 11888 29155 11940 29164
rect 11888 29121 11897 29155
rect 11897 29121 11931 29155
rect 11931 29121 11940 29155
rect 11888 29112 11940 29121
rect 14096 29112 14148 29164
rect 18696 29180 18748 29232
rect 18512 29112 18564 29164
rect 21548 29180 21600 29232
rect 8760 29044 8812 29096
rect 8852 29087 8904 29096
rect 8852 29053 8861 29087
rect 8861 29053 8895 29087
rect 8895 29053 8904 29087
rect 8852 29044 8904 29053
rect 11796 29087 11848 29096
rect 11796 29053 11805 29087
rect 11805 29053 11839 29087
rect 11839 29053 11848 29087
rect 11796 29044 11848 29053
rect 12532 29087 12584 29096
rect 12532 29053 12541 29087
rect 12541 29053 12575 29087
rect 12575 29053 12584 29087
rect 12532 29044 12584 29053
rect 13360 29087 13412 29096
rect 13360 29053 13369 29087
rect 13369 29053 13403 29087
rect 13403 29053 13412 29087
rect 13360 29044 13412 29053
rect 14188 29044 14240 29096
rect 9956 28976 10008 29028
rect 11244 28976 11296 29028
rect 12440 28976 12492 29028
rect 13544 28976 13596 29028
rect 16120 29044 16172 29096
rect 17040 29087 17092 29096
rect 17040 29053 17049 29087
rect 17049 29053 17083 29087
rect 17083 29053 17092 29087
rect 17040 29044 17092 29053
rect 19156 29044 19208 29096
rect 22100 29112 22152 29164
rect 23756 29112 23808 29164
rect 26240 29248 26292 29300
rect 24952 29180 25004 29232
rect 26792 29248 26844 29300
rect 27528 29248 27580 29300
rect 27620 29248 27672 29300
rect 28264 29291 28316 29300
rect 28264 29257 28273 29291
rect 28273 29257 28307 29291
rect 28307 29257 28316 29291
rect 28264 29248 28316 29257
rect 29000 29248 29052 29300
rect 29368 29248 29420 29300
rect 30656 29291 30708 29300
rect 30656 29257 30665 29291
rect 30665 29257 30699 29291
rect 30699 29257 30708 29291
rect 30656 29248 30708 29257
rect 31300 29248 31352 29300
rect 25136 29112 25188 29164
rect 25228 29155 25280 29164
rect 25228 29121 25237 29155
rect 25237 29121 25271 29155
rect 25271 29121 25280 29155
rect 25228 29112 25280 29121
rect 26056 29112 26108 29164
rect 16856 29019 16908 29028
rect 16856 28985 16865 29019
rect 16865 28985 16899 29019
rect 16899 28985 16908 29019
rect 16856 28976 16908 28985
rect 20720 28976 20772 29028
rect 14096 28951 14148 28960
rect 14096 28917 14105 28951
rect 14105 28917 14139 28951
rect 14139 28917 14148 28951
rect 14096 28908 14148 28917
rect 14648 28908 14700 28960
rect 15844 28951 15896 28960
rect 15844 28917 15853 28951
rect 15853 28917 15887 28951
rect 15887 28917 15896 28951
rect 15844 28908 15896 28917
rect 15936 28908 15988 28960
rect 20444 28908 20496 28960
rect 22652 28976 22704 29028
rect 26516 29112 26568 29164
rect 28172 29112 28224 29164
rect 25136 28976 25188 29028
rect 27620 29044 27672 29096
rect 27988 29087 28040 29096
rect 27988 29053 27997 29087
rect 27997 29053 28031 29087
rect 28031 29053 28040 29087
rect 27988 29044 28040 29053
rect 28632 29044 28684 29096
rect 28908 29087 28960 29096
rect 28908 29053 28917 29087
rect 28917 29053 28951 29087
rect 28951 29053 28960 29087
rect 28908 29044 28960 29053
rect 31392 29112 31444 29164
rect 30932 29087 30984 29096
rect 30932 29053 30941 29087
rect 30941 29053 30975 29087
rect 30975 29053 30984 29087
rect 30932 29044 30984 29053
rect 23572 28908 23624 28960
rect 23940 28951 23992 28960
rect 23940 28917 23949 28951
rect 23949 28917 23983 28951
rect 23983 28917 23992 28951
rect 23940 28908 23992 28917
rect 26056 28951 26108 28960
rect 26056 28917 26065 28951
rect 26065 28917 26099 28951
rect 26099 28917 26108 28951
rect 26056 28908 26108 28917
rect 26424 28908 26476 28960
rect 27896 28976 27948 29028
rect 26884 28908 26936 28960
rect 30012 28908 30064 28960
rect 30840 28951 30892 28960
rect 30840 28917 30849 28951
rect 30849 28917 30883 28951
rect 30883 28917 30892 28951
rect 30840 28908 30892 28917
rect 31300 28976 31352 29028
rect 31668 28908 31720 28960
rect 6946 28806 6998 28858
rect 7010 28806 7062 28858
rect 7074 28806 7126 28858
rect 7138 28806 7190 28858
rect 7202 28806 7254 28858
rect 14306 28806 14358 28858
rect 14370 28806 14422 28858
rect 14434 28806 14486 28858
rect 14498 28806 14550 28858
rect 14562 28806 14614 28858
rect 21666 28806 21718 28858
rect 21730 28806 21782 28858
rect 21794 28806 21846 28858
rect 21858 28806 21910 28858
rect 21922 28806 21974 28858
rect 29026 28806 29078 28858
rect 29090 28806 29142 28858
rect 29154 28806 29206 28858
rect 29218 28806 29270 28858
rect 29282 28806 29334 28858
rect 8852 28704 8904 28756
rect 12532 28704 12584 28756
rect 14648 28704 14700 28756
rect 15752 28747 15804 28756
rect 15752 28713 15761 28747
rect 15761 28713 15795 28747
rect 15795 28713 15804 28747
rect 15752 28704 15804 28713
rect 22652 28747 22704 28756
rect 22652 28713 22661 28747
rect 22661 28713 22695 28747
rect 22695 28713 22704 28747
rect 22652 28704 22704 28713
rect 23572 28747 23624 28756
rect 23572 28713 23581 28747
rect 23581 28713 23615 28747
rect 23615 28713 23624 28747
rect 23572 28704 23624 28713
rect 23940 28704 23992 28756
rect 27068 28704 27120 28756
rect 5264 28636 5316 28688
rect 15844 28636 15896 28688
rect 20352 28636 20404 28688
rect 21364 28636 21416 28688
rect 23480 28636 23532 28688
rect 5448 28500 5500 28552
rect 6644 28568 6696 28620
rect 8392 28568 8444 28620
rect 10876 28611 10928 28620
rect 6644 28432 6696 28484
rect 9496 28543 9548 28552
rect 9496 28509 9505 28543
rect 9505 28509 9539 28543
rect 9539 28509 9548 28543
rect 9496 28500 9548 28509
rect 10876 28577 10885 28611
rect 10885 28577 10919 28611
rect 10919 28577 10928 28611
rect 10876 28568 10928 28577
rect 12900 28611 12952 28620
rect 12900 28577 12909 28611
rect 12909 28577 12943 28611
rect 12943 28577 12952 28611
rect 12900 28568 12952 28577
rect 15936 28568 15988 28620
rect 22100 28568 22152 28620
rect 22560 28611 22612 28620
rect 22560 28577 22569 28611
rect 22569 28577 22603 28611
rect 22603 28577 22612 28611
rect 22560 28568 22612 28577
rect 10232 28543 10284 28552
rect 10232 28509 10241 28543
rect 10241 28509 10275 28543
rect 10275 28509 10284 28543
rect 10232 28500 10284 28509
rect 14004 28543 14056 28552
rect 14004 28509 14013 28543
rect 14013 28509 14047 28543
rect 14047 28509 14056 28543
rect 14004 28500 14056 28509
rect 17132 28543 17184 28552
rect 17132 28509 17141 28543
rect 17141 28509 17175 28543
rect 17175 28509 17184 28543
rect 17132 28500 17184 28509
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 24032 28636 24084 28688
rect 27528 28704 27580 28756
rect 28632 28747 28684 28756
rect 28632 28713 28641 28747
rect 28641 28713 28675 28747
rect 28675 28713 28684 28747
rect 28632 28704 28684 28713
rect 31116 28704 31168 28756
rect 23756 28611 23808 28620
rect 23756 28577 23765 28611
rect 23765 28577 23799 28611
rect 23799 28577 23808 28611
rect 23756 28568 23808 28577
rect 25136 28568 25188 28620
rect 26976 28500 27028 28552
rect 27528 28568 27580 28620
rect 27712 28568 27764 28620
rect 4252 28364 4304 28416
rect 5816 28407 5868 28416
rect 5816 28373 5825 28407
rect 5825 28373 5859 28407
rect 5859 28373 5868 28407
rect 5816 28364 5868 28373
rect 7840 28407 7892 28416
rect 7840 28373 7849 28407
rect 7849 28373 7883 28407
rect 7883 28373 7892 28407
rect 7840 28364 7892 28373
rect 9680 28364 9732 28416
rect 14648 28364 14700 28416
rect 16028 28364 16080 28416
rect 16212 28407 16264 28416
rect 16212 28373 16221 28407
rect 16221 28373 16255 28407
rect 16255 28373 16264 28407
rect 16212 28364 16264 28373
rect 16580 28407 16632 28416
rect 16580 28373 16589 28407
rect 16589 28373 16623 28407
rect 16623 28373 16632 28407
rect 16580 28364 16632 28373
rect 17776 28407 17828 28416
rect 17776 28373 17785 28407
rect 17785 28373 17819 28407
rect 17819 28373 17828 28407
rect 17776 28364 17828 28373
rect 20444 28407 20496 28416
rect 20444 28373 20453 28407
rect 20453 28373 20487 28407
rect 20487 28373 20496 28407
rect 20444 28364 20496 28373
rect 26424 28364 26476 28416
rect 27436 28432 27488 28484
rect 27896 28611 27948 28620
rect 27896 28577 27905 28611
rect 27905 28577 27939 28611
rect 27939 28577 27948 28611
rect 27896 28568 27948 28577
rect 28172 28500 28224 28552
rect 29552 28636 29604 28688
rect 30840 28636 30892 28688
rect 31668 28679 31720 28688
rect 31668 28645 31677 28679
rect 31677 28645 31711 28679
rect 31711 28645 31720 28679
rect 31668 28636 31720 28645
rect 28816 28611 28868 28620
rect 28816 28577 28825 28611
rect 28825 28577 28859 28611
rect 28859 28577 28868 28611
rect 28816 28568 28868 28577
rect 28908 28500 28960 28552
rect 29184 28432 29236 28484
rect 31208 28500 31260 28552
rect 30196 28364 30248 28416
rect 6286 28262 6338 28314
rect 6350 28262 6402 28314
rect 6414 28262 6466 28314
rect 6478 28262 6530 28314
rect 6542 28262 6594 28314
rect 13646 28262 13698 28314
rect 13710 28262 13762 28314
rect 13774 28262 13826 28314
rect 13838 28262 13890 28314
rect 13902 28262 13954 28314
rect 21006 28262 21058 28314
rect 21070 28262 21122 28314
rect 21134 28262 21186 28314
rect 21198 28262 21250 28314
rect 21262 28262 21314 28314
rect 28366 28262 28418 28314
rect 28430 28262 28482 28314
rect 28494 28262 28546 28314
rect 28558 28262 28610 28314
rect 28622 28262 28674 28314
rect 4988 28160 5040 28212
rect 5448 28203 5500 28212
rect 5448 28169 5457 28203
rect 5457 28169 5491 28203
rect 5491 28169 5500 28203
rect 5448 28160 5500 28169
rect 5816 28160 5868 28212
rect 9496 28160 9548 28212
rect 10232 28160 10284 28212
rect 3884 28067 3936 28076
rect 3884 28033 3893 28067
rect 3893 28033 3927 28067
rect 3927 28033 3936 28067
rect 3884 28024 3936 28033
rect 12072 28160 12124 28212
rect 12900 28160 12952 28212
rect 5540 27888 5592 27940
rect 6828 27888 6880 27940
rect 9864 27999 9916 28008
rect 9864 27965 9873 27999
rect 9873 27965 9907 27999
rect 9907 27965 9916 27999
rect 9864 27956 9916 27965
rect 7840 27888 7892 27940
rect 9772 27888 9824 27940
rect 10876 28092 10928 28144
rect 10600 27956 10652 28008
rect 11152 27956 11204 28008
rect 13360 28160 13412 28212
rect 14096 28067 14148 28076
rect 14096 28033 14105 28067
rect 14105 28033 14139 28067
rect 14139 28033 14148 28067
rect 14096 28024 14148 28033
rect 16120 28160 16172 28212
rect 19800 28160 19852 28212
rect 23848 28160 23900 28212
rect 24032 28160 24084 28212
rect 26608 28160 26660 28212
rect 28540 28160 28592 28212
rect 28724 28160 28776 28212
rect 28816 28160 28868 28212
rect 29460 28160 29512 28212
rect 30196 28160 30248 28212
rect 30380 28160 30432 28212
rect 15936 28024 15988 28076
rect 17040 28024 17092 28076
rect 10508 27888 10560 27940
rect 11060 27931 11112 27940
rect 11060 27897 11069 27931
rect 11069 27897 11103 27931
rect 11103 27897 11112 27931
rect 11060 27888 11112 27897
rect 6552 27820 6604 27872
rect 7288 27820 7340 27872
rect 7380 27820 7432 27872
rect 9036 27863 9088 27872
rect 9036 27829 9045 27863
rect 9045 27829 9079 27863
rect 9079 27829 9088 27863
rect 9036 27820 9088 27829
rect 10324 27863 10376 27872
rect 10324 27829 10333 27863
rect 10333 27829 10367 27863
rect 10367 27829 10376 27863
rect 10324 27820 10376 27829
rect 13544 27956 13596 28008
rect 11612 27931 11664 27940
rect 11612 27897 11621 27931
rect 11621 27897 11655 27931
rect 11655 27897 11664 27931
rect 11612 27888 11664 27897
rect 16212 27956 16264 28008
rect 19708 27999 19760 28008
rect 19708 27965 19717 27999
rect 19717 27965 19751 27999
rect 19751 27965 19760 27999
rect 19708 27956 19760 27965
rect 22100 27956 22152 28008
rect 23112 27956 23164 28008
rect 23572 27999 23624 28008
rect 23572 27965 23597 27999
rect 23597 27965 23624 27999
rect 23572 27956 23624 27965
rect 23664 27999 23716 28008
rect 23664 27965 23673 27999
rect 23673 27965 23707 27999
rect 23707 27965 23716 27999
rect 23664 27956 23716 27965
rect 24492 28092 24544 28144
rect 27620 28092 27672 28144
rect 28264 28135 28316 28144
rect 28264 28101 28273 28135
rect 28273 28101 28307 28135
rect 28307 28101 28316 28135
rect 28264 28092 28316 28101
rect 26056 28067 26108 28076
rect 26056 28033 26065 28067
rect 26065 28033 26099 28067
rect 26099 28033 26108 28067
rect 26056 28024 26108 28033
rect 27896 28024 27948 28076
rect 28724 28067 28776 28076
rect 28724 28033 28733 28067
rect 28733 28033 28767 28067
rect 28767 28033 28776 28067
rect 28724 28024 28776 28033
rect 29184 28135 29236 28144
rect 29184 28101 29193 28135
rect 29193 28101 29227 28135
rect 29227 28101 29236 28135
rect 29184 28092 29236 28101
rect 29644 28092 29696 28144
rect 29920 28092 29972 28144
rect 31116 28092 31168 28144
rect 29368 28024 29420 28076
rect 30196 28024 30248 28076
rect 24400 27956 24452 28008
rect 24584 27999 24636 28008
rect 24584 27965 24593 27999
rect 24593 27965 24627 27999
rect 24627 27965 24636 27999
rect 24584 27956 24636 27965
rect 14004 27888 14056 27940
rect 11428 27820 11480 27872
rect 16304 27820 16356 27872
rect 17960 27931 18012 27940
rect 17960 27897 17969 27931
rect 17969 27897 18003 27931
rect 18003 27897 18012 27931
rect 17960 27888 18012 27897
rect 25136 27956 25188 28008
rect 26700 27999 26752 28008
rect 26700 27965 26709 27999
rect 26709 27965 26743 27999
rect 26743 27965 26752 27999
rect 26700 27956 26752 27965
rect 26884 27999 26936 28008
rect 26884 27965 26893 27999
rect 26893 27965 26927 27999
rect 26927 27965 26936 27999
rect 26884 27956 26936 27965
rect 27620 27956 27672 28008
rect 17592 27820 17644 27872
rect 22744 27863 22796 27872
rect 22744 27829 22753 27863
rect 22753 27829 22787 27863
rect 22787 27829 22796 27863
rect 22744 27820 22796 27829
rect 26424 27931 26476 27940
rect 26424 27897 26433 27931
rect 26433 27897 26467 27931
rect 26467 27897 26476 27931
rect 26424 27888 26476 27897
rect 27252 27888 27304 27940
rect 27528 27888 27580 27940
rect 28172 27888 28224 27940
rect 28632 27999 28684 28008
rect 28632 27965 28641 27999
rect 28641 27965 28675 27999
rect 28675 27965 28684 27999
rect 28632 27956 28684 27965
rect 30104 27956 30156 28008
rect 29460 27931 29512 27940
rect 24308 27863 24360 27872
rect 24308 27829 24317 27863
rect 24317 27829 24351 27863
rect 24351 27829 24360 27863
rect 24308 27820 24360 27829
rect 25596 27820 25648 27872
rect 25872 27820 25924 27872
rect 26976 27863 27028 27872
rect 26976 27829 26985 27863
rect 26985 27829 27019 27863
rect 27019 27829 27028 27863
rect 26976 27820 27028 27829
rect 27804 27820 27856 27872
rect 29460 27897 29469 27931
rect 29469 27897 29503 27931
rect 29503 27897 29512 27931
rect 29460 27888 29512 27897
rect 28816 27820 28868 27872
rect 29920 27820 29972 27872
rect 30748 27820 30800 27872
rect 30840 27863 30892 27872
rect 30840 27829 30865 27863
rect 30865 27829 30892 27863
rect 30840 27820 30892 27829
rect 31208 27820 31260 27872
rect 31852 27863 31904 27872
rect 31852 27829 31861 27863
rect 31861 27829 31895 27863
rect 31895 27829 31904 27863
rect 31852 27820 31904 27829
rect 6946 27718 6998 27770
rect 7010 27718 7062 27770
rect 7074 27718 7126 27770
rect 7138 27718 7190 27770
rect 7202 27718 7254 27770
rect 14306 27718 14358 27770
rect 14370 27718 14422 27770
rect 14434 27718 14486 27770
rect 14498 27718 14550 27770
rect 14562 27718 14614 27770
rect 21666 27718 21718 27770
rect 21730 27718 21782 27770
rect 21794 27718 21846 27770
rect 21858 27718 21910 27770
rect 21922 27718 21974 27770
rect 29026 27718 29078 27770
rect 29090 27718 29142 27770
rect 29154 27718 29206 27770
rect 29218 27718 29270 27770
rect 29282 27718 29334 27770
rect 5264 27616 5316 27668
rect 6644 27616 6696 27668
rect 6552 27548 6604 27600
rect 6920 27548 6972 27600
rect 1308 27412 1360 27464
rect 6184 27480 6236 27532
rect 5540 27319 5592 27328
rect 5540 27285 5549 27319
rect 5549 27285 5583 27319
rect 5583 27285 5592 27319
rect 5540 27276 5592 27285
rect 6828 27523 6880 27532
rect 6828 27489 6837 27523
rect 6837 27489 6871 27523
rect 6871 27489 6880 27523
rect 6828 27480 6880 27489
rect 7288 27616 7340 27668
rect 8944 27616 8996 27668
rect 10324 27616 10376 27668
rect 7196 27548 7248 27600
rect 9680 27548 9732 27600
rect 11612 27616 11664 27668
rect 14004 27616 14056 27668
rect 14740 27616 14792 27668
rect 17960 27616 18012 27668
rect 9036 27480 9088 27532
rect 12440 27591 12492 27600
rect 12440 27557 12449 27591
rect 12449 27557 12483 27591
rect 12483 27557 12492 27591
rect 12440 27548 12492 27557
rect 13452 27548 13504 27600
rect 14924 27548 14976 27600
rect 16028 27548 16080 27600
rect 20444 27548 20496 27600
rect 23940 27616 23992 27668
rect 24400 27616 24452 27668
rect 24768 27616 24820 27668
rect 25688 27616 25740 27668
rect 26884 27616 26936 27668
rect 28172 27616 28224 27668
rect 30380 27616 30432 27668
rect 30748 27659 30800 27668
rect 30748 27625 30757 27659
rect 30757 27625 30791 27659
rect 30791 27625 30800 27659
rect 30748 27616 30800 27625
rect 6644 27276 6696 27328
rect 6828 27344 6880 27396
rect 8116 27455 8168 27464
rect 8116 27421 8125 27455
rect 8125 27421 8159 27455
rect 8159 27421 8168 27455
rect 8116 27412 8168 27421
rect 12164 27523 12216 27532
rect 12164 27489 12173 27523
rect 12173 27489 12207 27523
rect 12207 27489 12216 27523
rect 12164 27480 12216 27489
rect 14464 27480 14516 27532
rect 16304 27480 16356 27532
rect 16764 27480 16816 27532
rect 9772 27344 9824 27396
rect 10324 27455 10376 27464
rect 10324 27421 10333 27455
rect 10333 27421 10367 27455
rect 10367 27421 10376 27455
rect 10324 27412 10376 27421
rect 11796 27387 11848 27396
rect 11796 27353 11805 27387
rect 11805 27353 11839 27387
rect 11839 27353 11848 27387
rect 11796 27344 11848 27353
rect 12532 27455 12584 27464
rect 12532 27421 12541 27455
rect 12541 27421 12575 27455
rect 12575 27421 12584 27455
rect 12532 27412 12584 27421
rect 12348 27344 12400 27396
rect 14372 27412 14424 27464
rect 7656 27276 7708 27328
rect 8392 27276 8444 27328
rect 8760 27319 8812 27328
rect 8760 27285 8769 27319
rect 8769 27285 8803 27319
rect 8803 27285 8812 27319
rect 8760 27276 8812 27285
rect 10048 27276 10100 27328
rect 14188 27276 14240 27328
rect 14740 27455 14792 27464
rect 14740 27421 14749 27455
rect 14749 27421 14783 27455
rect 14783 27421 14792 27455
rect 14740 27412 14792 27421
rect 15016 27455 15068 27464
rect 15016 27421 15025 27455
rect 15025 27421 15059 27455
rect 15059 27421 15068 27455
rect 15016 27412 15068 27421
rect 17132 27412 17184 27464
rect 17500 27523 17552 27532
rect 17500 27489 17509 27523
rect 17509 27489 17543 27523
rect 17543 27489 17552 27523
rect 17500 27480 17552 27489
rect 17684 27523 17736 27532
rect 17684 27489 17693 27523
rect 17693 27489 17727 27523
rect 17727 27489 17736 27523
rect 17684 27480 17736 27489
rect 18972 27480 19024 27532
rect 19708 27480 19760 27532
rect 23572 27548 23624 27600
rect 24032 27548 24084 27600
rect 24308 27548 24360 27600
rect 26424 27548 26476 27600
rect 27344 27548 27396 27600
rect 19248 27455 19300 27464
rect 19248 27421 19257 27455
rect 19257 27421 19291 27455
rect 19291 27421 19300 27455
rect 19248 27412 19300 27421
rect 19800 27412 19852 27464
rect 22008 27523 22060 27532
rect 22008 27489 22017 27523
rect 22017 27489 22051 27523
rect 22051 27489 22060 27523
rect 22008 27480 22060 27489
rect 22744 27412 22796 27464
rect 23112 27412 23164 27464
rect 16856 27276 16908 27328
rect 17132 27319 17184 27328
rect 17132 27285 17141 27319
rect 17141 27285 17175 27319
rect 17175 27285 17184 27319
rect 17132 27276 17184 27285
rect 17684 27276 17736 27328
rect 19064 27319 19116 27328
rect 19064 27285 19073 27319
rect 19073 27285 19107 27319
rect 19107 27285 19116 27319
rect 19064 27276 19116 27285
rect 19156 27276 19208 27328
rect 19984 27319 20036 27328
rect 19984 27285 19993 27319
rect 19993 27285 20027 27319
rect 20027 27285 20036 27319
rect 19984 27276 20036 27285
rect 22100 27319 22152 27328
rect 22100 27285 22109 27319
rect 22109 27285 22143 27319
rect 22143 27285 22152 27319
rect 22100 27276 22152 27285
rect 22192 27276 22244 27328
rect 23112 27276 23164 27328
rect 23388 27480 23440 27532
rect 23664 27412 23716 27464
rect 24584 27412 24636 27464
rect 26056 27480 26108 27532
rect 27620 27480 27672 27532
rect 30564 27548 30616 27600
rect 31116 27591 31168 27600
rect 31116 27557 31125 27591
rect 31125 27557 31159 27591
rect 31159 27557 31168 27591
rect 31116 27548 31168 27557
rect 31852 27548 31904 27600
rect 28172 27480 28224 27532
rect 28540 27480 28592 27532
rect 29000 27480 29052 27532
rect 29552 27480 29604 27532
rect 29736 27523 29788 27532
rect 29736 27489 29745 27523
rect 29745 27489 29779 27523
rect 29779 27489 29788 27523
rect 29736 27480 29788 27489
rect 30840 27480 30892 27532
rect 31300 27480 31352 27532
rect 26884 27455 26936 27464
rect 26884 27421 26893 27455
rect 26893 27421 26927 27455
rect 26927 27421 26936 27455
rect 26884 27412 26936 27421
rect 24032 27344 24084 27396
rect 24952 27387 25004 27396
rect 24952 27353 24961 27387
rect 24961 27353 24995 27387
rect 24995 27353 25004 27387
rect 24952 27344 25004 27353
rect 23572 27276 23624 27328
rect 24216 27319 24268 27328
rect 24216 27285 24225 27319
rect 24225 27285 24259 27319
rect 24259 27285 24268 27319
rect 24216 27276 24268 27285
rect 24492 27276 24544 27328
rect 24584 27276 24636 27328
rect 26792 27344 26844 27396
rect 27436 27344 27488 27396
rect 27988 27455 28040 27464
rect 27988 27421 27997 27455
rect 27997 27421 28031 27455
rect 28031 27421 28040 27455
rect 27988 27412 28040 27421
rect 28632 27412 28684 27464
rect 29552 27344 29604 27396
rect 25504 27319 25556 27328
rect 25504 27285 25513 27319
rect 25513 27285 25547 27319
rect 25547 27285 25556 27319
rect 25504 27276 25556 27285
rect 25596 27319 25648 27328
rect 25596 27285 25605 27319
rect 25605 27285 25639 27319
rect 25639 27285 25648 27319
rect 25596 27276 25648 27285
rect 26056 27319 26108 27328
rect 26056 27285 26065 27319
rect 26065 27285 26099 27319
rect 26099 27285 26108 27319
rect 26056 27276 26108 27285
rect 26332 27319 26384 27328
rect 26332 27285 26341 27319
rect 26341 27285 26375 27319
rect 26375 27285 26384 27319
rect 26332 27276 26384 27285
rect 26608 27276 26660 27328
rect 28908 27276 28960 27328
rect 30380 27412 30432 27464
rect 30656 27455 30708 27464
rect 30656 27421 30665 27455
rect 30665 27421 30699 27455
rect 30699 27421 30708 27455
rect 30656 27412 30708 27421
rect 30932 27412 30984 27464
rect 30472 27276 30524 27328
rect 6286 27174 6338 27226
rect 6350 27174 6402 27226
rect 6414 27174 6466 27226
rect 6478 27174 6530 27226
rect 6542 27174 6594 27226
rect 13646 27174 13698 27226
rect 13710 27174 13762 27226
rect 13774 27174 13826 27226
rect 13838 27174 13890 27226
rect 13902 27174 13954 27226
rect 21006 27174 21058 27226
rect 21070 27174 21122 27226
rect 21134 27174 21186 27226
rect 21198 27174 21250 27226
rect 21262 27174 21314 27226
rect 28366 27174 28418 27226
rect 28430 27174 28482 27226
rect 28494 27174 28546 27226
rect 28558 27174 28610 27226
rect 28622 27174 28674 27226
rect 8116 27072 8168 27124
rect 9864 27072 9916 27124
rect 10324 27072 10376 27124
rect 11152 27072 11204 27124
rect 11428 27072 11480 27124
rect 15016 27072 15068 27124
rect 8944 27004 8996 27056
rect 9956 26936 10008 26988
rect 6184 26868 6236 26920
rect 6644 26732 6696 26784
rect 7748 26800 7800 26852
rect 8484 26800 8536 26852
rect 9404 26911 9456 26920
rect 9404 26877 9413 26911
rect 9413 26877 9447 26911
rect 9447 26877 9456 26911
rect 9404 26868 9456 26877
rect 9680 26868 9732 26920
rect 10600 27004 10652 27056
rect 9588 26800 9640 26852
rect 10968 26911 11020 26920
rect 10968 26877 10977 26911
rect 10977 26877 11011 26911
rect 11011 26877 11020 26911
rect 10968 26868 11020 26877
rect 11244 26979 11296 26988
rect 11244 26945 11253 26979
rect 11253 26945 11287 26979
rect 11287 26945 11296 26979
rect 11244 26936 11296 26945
rect 17500 27072 17552 27124
rect 19984 27072 20036 27124
rect 23112 27115 23164 27124
rect 23112 27081 23121 27115
rect 23121 27081 23155 27115
rect 23155 27081 23164 27115
rect 23112 27072 23164 27081
rect 23664 27072 23716 27124
rect 24216 27072 24268 27124
rect 26332 27115 26384 27124
rect 26332 27081 26362 27115
rect 26362 27081 26384 27115
rect 26332 27072 26384 27081
rect 27988 27072 28040 27124
rect 11152 26800 11204 26852
rect 14372 26936 14424 26988
rect 14096 26911 14148 26920
rect 14096 26877 14105 26911
rect 14105 26877 14139 26911
rect 14139 26877 14148 26911
rect 14096 26868 14148 26877
rect 14924 26868 14976 26920
rect 15200 26911 15252 26920
rect 15200 26877 15209 26911
rect 15209 26877 15243 26911
rect 15243 26877 15252 26911
rect 15200 26868 15252 26877
rect 17776 26936 17828 26988
rect 20536 26936 20588 26988
rect 21364 26979 21416 26988
rect 21364 26945 21373 26979
rect 21373 26945 21407 26979
rect 21407 26945 21416 26979
rect 21364 26936 21416 26945
rect 25780 27047 25832 27056
rect 17316 26911 17368 26920
rect 17316 26877 17325 26911
rect 17325 26877 17359 26911
rect 17359 26877 17368 26911
rect 17316 26868 17368 26877
rect 7840 26732 7892 26784
rect 9864 26732 9916 26784
rect 10048 26732 10100 26784
rect 12348 26800 12400 26852
rect 12440 26843 12492 26852
rect 12440 26809 12449 26843
rect 12449 26809 12483 26843
rect 12483 26809 12492 26843
rect 12440 26800 12492 26809
rect 17132 26800 17184 26852
rect 19064 26800 19116 26852
rect 19524 26800 19576 26852
rect 12624 26732 12676 26784
rect 14924 26732 14976 26784
rect 16672 26775 16724 26784
rect 16672 26741 16681 26775
rect 16681 26741 16715 26775
rect 16715 26741 16724 26775
rect 16672 26732 16724 26741
rect 17500 26732 17552 26784
rect 20076 26732 20128 26784
rect 22100 26800 22152 26852
rect 24124 26868 24176 26920
rect 24492 26911 24544 26920
rect 24492 26877 24501 26911
rect 24501 26877 24535 26911
rect 24535 26877 24544 26911
rect 24492 26868 24544 26877
rect 23572 26843 23624 26852
rect 23572 26809 23581 26843
rect 23581 26809 23615 26843
rect 23615 26809 23624 26843
rect 23572 26800 23624 26809
rect 25780 27013 25789 27047
rect 25789 27013 25823 27047
rect 25823 27013 25832 27047
rect 25780 27004 25832 27013
rect 25872 27004 25924 27056
rect 29828 27072 29880 27124
rect 30840 27072 30892 27124
rect 25688 26936 25740 26988
rect 25412 26911 25464 26920
rect 25412 26877 25421 26911
rect 25421 26877 25455 26911
rect 25455 26877 25464 26911
rect 25412 26868 25464 26877
rect 28908 27004 28960 27056
rect 24860 26843 24912 26852
rect 24860 26809 24869 26843
rect 24869 26809 24903 26843
rect 24903 26809 24912 26843
rect 24860 26800 24912 26809
rect 25044 26800 25096 26852
rect 30472 27047 30524 27056
rect 30472 27013 30481 27047
rect 30481 27013 30515 27047
rect 30515 27013 30524 27047
rect 30472 27004 30524 27013
rect 27896 26868 27948 26920
rect 28448 26911 28500 26920
rect 28448 26877 28457 26911
rect 28457 26877 28491 26911
rect 28491 26877 28500 26911
rect 28448 26868 28500 26877
rect 30564 26868 30616 26920
rect 33140 26868 33192 26920
rect 24492 26732 24544 26784
rect 24952 26732 25004 26784
rect 25596 26775 25648 26784
rect 25596 26741 25605 26775
rect 25605 26741 25639 26775
rect 25639 26741 25648 26775
rect 25596 26732 25648 26741
rect 26148 26732 26200 26784
rect 26332 26732 26384 26784
rect 27344 26732 27396 26784
rect 27896 26775 27948 26784
rect 27896 26741 27905 26775
rect 27905 26741 27939 26775
rect 27939 26741 27948 26775
rect 27896 26732 27948 26741
rect 30104 26800 30156 26852
rect 29368 26732 29420 26784
rect 29460 26732 29512 26784
rect 30380 26732 30432 26784
rect 31392 26732 31444 26784
rect 6946 26630 6998 26682
rect 7010 26630 7062 26682
rect 7074 26630 7126 26682
rect 7138 26630 7190 26682
rect 7202 26630 7254 26682
rect 14306 26630 14358 26682
rect 14370 26630 14422 26682
rect 14434 26630 14486 26682
rect 14498 26630 14550 26682
rect 14562 26630 14614 26682
rect 21666 26630 21718 26682
rect 21730 26630 21782 26682
rect 21794 26630 21846 26682
rect 21858 26630 21910 26682
rect 21922 26630 21974 26682
rect 29026 26630 29078 26682
rect 29090 26630 29142 26682
rect 29154 26630 29206 26682
rect 29218 26630 29270 26682
rect 29282 26630 29334 26682
rect 6828 26528 6880 26580
rect 7748 26571 7800 26580
rect 7748 26537 7757 26571
rect 7757 26537 7791 26571
rect 7791 26537 7800 26571
rect 7748 26528 7800 26537
rect 6644 26460 6696 26512
rect 8392 26571 8444 26580
rect 8392 26537 8401 26571
rect 8401 26537 8435 26571
rect 8435 26537 8444 26571
rect 8392 26528 8444 26537
rect 8760 26528 8812 26580
rect 9404 26528 9456 26580
rect 10324 26528 10376 26580
rect 10600 26528 10652 26580
rect 9312 26460 9364 26512
rect 4528 26435 4580 26444
rect 4528 26401 4537 26435
rect 4537 26401 4571 26435
rect 4571 26401 4580 26435
rect 4528 26392 4580 26401
rect 5816 26392 5868 26444
rect 7840 26435 7892 26444
rect 7840 26401 7849 26435
rect 7849 26401 7883 26435
rect 7883 26401 7892 26435
rect 7840 26392 7892 26401
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 7380 26367 7432 26376
rect 7380 26333 7389 26367
rect 7389 26333 7423 26367
rect 7423 26333 7432 26367
rect 7380 26324 7432 26333
rect 8484 26324 8536 26376
rect 9036 26435 9088 26444
rect 9036 26401 9045 26435
rect 9045 26401 9079 26435
rect 9079 26401 9088 26435
rect 9036 26392 9088 26401
rect 10600 26435 10652 26444
rect 10600 26401 10609 26435
rect 10609 26401 10643 26435
rect 10643 26401 10652 26435
rect 10600 26392 10652 26401
rect 11244 26528 11296 26580
rect 10876 26460 10928 26512
rect 12164 26460 12216 26512
rect 11428 26392 11480 26444
rect 11612 26435 11664 26444
rect 11612 26401 11621 26435
rect 11621 26401 11655 26435
rect 11655 26401 11664 26435
rect 11612 26392 11664 26401
rect 12440 26528 12492 26580
rect 14832 26528 14884 26580
rect 15200 26528 15252 26580
rect 15384 26528 15436 26580
rect 17040 26528 17092 26580
rect 19248 26528 19300 26580
rect 19524 26528 19576 26580
rect 13268 26460 13320 26512
rect 14740 26460 14792 26512
rect 12624 26392 12676 26444
rect 5172 26231 5224 26240
rect 5172 26197 5181 26231
rect 5181 26197 5215 26231
rect 5215 26197 5224 26231
rect 5172 26188 5224 26197
rect 8116 26188 8168 26240
rect 13360 26367 13412 26376
rect 13360 26333 13369 26367
rect 13369 26333 13403 26367
rect 13403 26333 13412 26367
rect 13360 26324 13412 26333
rect 14188 26324 14240 26376
rect 18880 26392 18932 26444
rect 9220 26256 9272 26308
rect 9588 26188 9640 26240
rect 10048 26188 10100 26240
rect 10508 26188 10560 26240
rect 11520 26188 11572 26240
rect 11888 26231 11940 26240
rect 11888 26197 11897 26231
rect 11897 26197 11931 26231
rect 11931 26197 11940 26231
rect 11888 26188 11940 26197
rect 14648 26256 14700 26308
rect 15568 26299 15620 26308
rect 13452 26188 13504 26240
rect 15568 26265 15577 26299
rect 15577 26265 15611 26299
rect 15611 26265 15620 26299
rect 15568 26256 15620 26265
rect 15108 26231 15160 26240
rect 15108 26197 15117 26231
rect 15117 26197 15151 26231
rect 15151 26197 15160 26231
rect 15108 26188 15160 26197
rect 15936 26188 15988 26240
rect 16672 26367 16724 26376
rect 16672 26333 16681 26367
rect 16681 26333 16715 26367
rect 16715 26333 16724 26367
rect 16672 26324 16724 26333
rect 18420 26324 18472 26376
rect 19156 26460 19208 26512
rect 19800 26571 19852 26580
rect 19800 26537 19809 26571
rect 19809 26537 19843 26571
rect 19843 26537 19852 26571
rect 19800 26528 19852 26537
rect 20076 26528 20128 26580
rect 16764 26188 16816 26240
rect 18512 26188 18564 26240
rect 19432 26324 19484 26376
rect 22192 26528 22244 26580
rect 23388 26528 23440 26580
rect 22468 26460 22520 26512
rect 25044 26528 25096 26580
rect 25412 26528 25464 26580
rect 26884 26528 26936 26580
rect 27344 26571 27396 26580
rect 21456 26392 21508 26444
rect 25688 26460 25740 26512
rect 23480 26435 23532 26444
rect 23480 26401 23489 26435
rect 23489 26401 23523 26435
rect 23523 26401 23532 26435
rect 23480 26392 23532 26401
rect 26332 26460 26384 26512
rect 26516 26503 26568 26512
rect 26516 26469 26525 26503
rect 26525 26469 26559 26503
rect 26559 26469 26568 26503
rect 26516 26460 26568 26469
rect 26608 26503 26660 26512
rect 26608 26469 26617 26503
rect 26617 26469 26651 26503
rect 26651 26469 26660 26503
rect 26608 26460 26660 26469
rect 26792 26460 26844 26512
rect 20076 26256 20128 26308
rect 25228 26324 25280 26376
rect 27344 26537 27353 26571
rect 27353 26537 27387 26571
rect 27387 26537 27396 26571
rect 27344 26528 27396 26537
rect 27528 26571 27580 26580
rect 27528 26537 27537 26571
rect 27537 26537 27571 26571
rect 27571 26537 27580 26571
rect 27528 26528 27580 26537
rect 28448 26528 28500 26580
rect 24952 26256 25004 26308
rect 26424 26256 26476 26308
rect 26976 26324 27028 26376
rect 27804 26392 27856 26444
rect 27712 26299 27764 26308
rect 27712 26265 27721 26299
rect 27721 26265 27755 26299
rect 27755 26265 27764 26299
rect 28264 26435 28316 26444
rect 28264 26401 28273 26435
rect 28273 26401 28307 26435
rect 28307 26401 28316 26435
rect 28264 26392 28316 26401
rect 29092 26460 29144 26512
rect 29460 26528 29512 26580
rect 30656 26571 30708 26580
rect 30656 26537 30665 26571
rect 30665 26537 30699 26571
rect 30699 26537 30708 26571
rect 30656 26528 30708 26537
rect 28632 26392 28684 26444
rect 28816 26435 28868 26444
rect 28816 26401 28825 26435
rect 28825 26401 28859 26435
rect 28859 26401 28868 26435
rect 28816 26392 28868 26401
rect 30932 26435 30984 26444
rect 30932 26401 30941 26435
rect 30941 26401 30975 26435
rect 30975 26401 30984 26435
rect 30932 26392 30984 26401
rect 28172 26324 28224 26376
rect 27712 26256 27764 26265
rect 30288 26256 30340 26308
rect 20628 26231 20680 26240
rect 20628 26197 20637 26231
rect 20637 26197 20671 26231
rect 20671 26197 20680 26231
rect 20628 26188 20680 26197
rect 24860 26188 24912 26240
rect 28816 26188 28868 26240
rect 28908 26188 28960 26240
rect 6286 26086 6338 26138
rect 6350 26086 6402 26138
rect 6414 26086 6466 26138
rect 6478 26086 6530 26138
rect 6542 26086 6594 26138
rect 13646 26086 13698 26138
rect 13710 26086 13762 26138
rect 13774 26086 13826 26138
rect 13838 26086 13890 26138
rect 13902 26086 13954 26138
rect 21006 26086 21058 26138
rect 21070 26086 21122 26138
rect 21134 26086 21186 26138
rect 21198 26086 21250 26138
rect 21262 26086 21314 26138
rect 28366 26086 28418 26138
rect 28430 26086 28482 26138
rect 28494 26086 28546 26138
rect 28558 26086 28610 26138
rect 28622 26086 28674 26138
rect 4528 25984 4580 26036
rect 9036 25984 9088 26036
rect 9588 25984 9640 26036
rect 10324 26027 10376 26036
rect 10324 25993 10333 26027
rect 10333 25993 10367 26027
rect 10367 25993 10376 26027
rect 10324 25984 10376 25993
rect 10876 26027 10928 26036
rect 10876 25993 10885 26027
rect 10885 25993 10919 26027
rect 10919 25993 10928 26027
rect 10876 25984 10928 25993
rect 11612 25984 11664 26036
rect 4252 25848 4304 25900
rect 5816 25848 5868 25900
rect 8484 25823 8536 25832
rect 8484 25789 8493 25823
rect 8493 25789 8527 25823
rect 8527 25789 8536 25823
rect 8484 25780 8536 25789
rect 9404 25780 9456 25832
rect 4988 25755 5040 25764
rect 4988 25721 4997 25755
rect 4997 25721 5031 25755
rect 5031 25721 5040 25755
rect 4988 25712 5040 25721
rect 7748 25712 7800 25764
rect 8208 25755 8260 25764
rect 8208 25721 8217 25755
rect 8217 25721 8251 25755
rect 8251 25721 8260 25755
rect 8208 25712 8260 25721
rect 5264 25644 5316 25696
rect 5632 25687 5684 25696
rect 5632 25653 5641 25687
rect 5641 25653 5675 25687
rect 5675 25653 5684 25687
rect 5632 25644 5684 25653
rect 6184 25687 6236 25696
rect 6184 25653 6193 25687
rect 6193 25653 6227 25687
rect 6227 25653 6236 25687
rect 6184 25644 6236 25653
rect 7288 25644 7340 25696
rect 7840 25644 7892 25696
rect 8576 25687 8628 25696
rect 8576 25653 8585 25687
rect 8585 25653 8619 25687
rect 8619 25653 8628 25687
rect 8576 25644 8628 25653
rect 9312 25687 9364 25696
rect 9312 25653 9321 25687
rect 9321 25653 9355 25687
rect 9355 25653 9364 25687
rect 9312 25644 9364 25653
rect 9588 25644 9640 25696
rect 10968 25916 11020 25968
rect 17316 25984 17368 26036
rect 19708 25984 19760 26036
rect 21456 25984 21508 26036
rect 25228 26027 25280 26036
rect 25228 25993 25237 26027
rect 25237 25993 25271 26027
rect 25271 25993 25280 26027
rect 25228 25984 25280 25993
rect 29368 25984 29420 26036
rect 10600 25780 10652 25832
rect 10784 25780 10836 25832
rect 11336 25848 11388 25900
rect 13268 25848 13320 25900
rect 15292 25891 15344 25900
rect 15292 25857 15301 25891
rect 15301 25857 15335 25891
rect 15335 25857 15344 25891
rect 15292 25848 15344 25857
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 10508 25644 10560 25696
rect 12808 25823 12860 25832
rect 12808 25789 12817 25823
rect 12817 25789 12851 25823
rect 12851 25789 12860 25823
rect 12808 25780 12860 25789
rect 14740 25823 14792 25832
rect 14740 25789 14749 25823
rect 14749 25789 14783 25823
rect 14783 25789 14792 25823
rect 14740 25780 14792 25789
rect 16304 25823 16356 25832
rect 16304 25789 16313 25823
rect 16313 25789 16347 25823
rect 16347 25789 16356 25823
rect 16304 25780 16356 25789
rect 17224 25823 17276 25832
rect 17224 25789 17233 25823
rect 17233 25789 17267 25823
rect 17267 25789 17276 25823
rect 17224 25780 17276 25789
rect 18420 25848 18472 25900
rect 19616 25848 19668 25900
rect 19892 25848 19944 25900
rect 28908 25916 28960 25968
rect 13176 25755 13228 25764
rect 13176 25721 13185 25755
rect 13185 25721 13219 25755
rect 13219 25721 13228 25755
rect 13176 25712 13228 25721
rect 15108 25712 15160 25764
rect 11428 25644 11480 25696
rect 14096 25644 14148 25696
rect 15476 25644 15528 25696
rect 16488 25687 16540 25696
rect 16488 25653 16497 25687
rect 16497 25653 16531 25687
rect 16531 25653 16540 25687
rect 16488 25644 16540 25653
rect 17500 25644 17552 25696
rect 20536 25823 20588 25832
rect 20536 25789 20545 25823
rect 20545 25789 20579 25823
rect 20579 25789 20588 25823
rect 20536 25780 20588 25789
rect 21456 25823 21508 25832
rect 21456 25789 21465 25823
rect 21465 25789 21499 25823
rect 21499 25789 21508 25823
rect 21456 25780 21508 25789
rect 18512 25687 18564 25696
rect 18512 25653 18521 25687
rect 18521 25653 18555 25687
rect 18555 25653 18564 25687
rect 18512 25644 18564 25653
rect 19432 25644 19484 25696
rect 19892 25644 19944 25696
rect 20628 25712 20680 25764
rect 22008 25712 22060 25764
rect 23480 25780 23532 25832
rect 22284 25712 22336 25764
rect 22376 25755 22428 25764
rect 22376 25721 22385 25755
rect 22385 25721 22419 25755
rect 22419 25721 22428 25755
rect 22376 25712 22428 25721
rect 28172 25848 28224 25900
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 25320 25780 25372 25832
rect 25872 25780 25924 25832
rect 26332 25780 26384 25832
rect 28816 25780 28868 25832
rect 30380 25823 30432 25832
rect 30380 25789 30389 25823
rect 30389 25789 30423 25823
rect 30423 25789 30432 25823
rect 30380 25780 30432 25789
rect 27896 25712 27948 25764
rect 30104 25712 30156 25764
rect 23848 25687 23900 25696
rect 23848 25653 23857 25687
rect 23857 25653 23891 25687
rect 23891 25653 23900 25687
rect 23848 25644 23900 25653
rect 25504 25644 25556 25696
rect 26608 25644 26660 25696
rect 29092 25644 29144 25696
rect 6946 25542 6998 25594
rect 7010 25542 7062 25594
rect 7074 25542 7126 25594
rect 7138 25542 7190 25594
rect 7202 25542 7254 25594
rect 14306 25542 14358 25594
rect 14370 25542 14422 25594
rect 14434 25542 14486 25594
rect 14498 25542 14550 25594
rect 14562 25542 14614 25594
rect 21666 25542 21718 25594
rect 21730 25542 21782 25594
rect 21794 25542 21846 25594
rect 21858 25542 21910 25594
rect 21922 25542 21974 25594
rect 29026 25542 29078 25594
rect 29090 25542 29142 25594
rect 29154 25542 29206 25594
rect 29218 25542 29270 25594
rect 29282 25542 29334 25594
rect 4988 25440 5040 25492
rect 5172 25440 5224 25492
rect 5264 25440 5316 25492
rect 5816 25415 5868 25424
rect 5816 25381 5825 25415
rect 5825 25381 5859 25415
rect 5859 25381 5868 25415
rect 5816 25372 5868 25381
rect 6184 25372 6236 25424
rect 7748 25483 7800 25492
rect 7748 25449 7757 25483
rect 7757 25449 7791 25483
rect 7791 25449 7800 25483
rect 7748 25440 7800 25449
rect 8208 25440 8260 25492
rect 9312 25440 9364 25492
rect 10968 25440 11020 25492
rect 11612 25440 11664 25492
rect 11888 25440 11940 25492
rect 12808 25440 12860 25492
rect 13176 25440 13228 25492
rect 14740 25440 14792 25492
rect 3424 25279 3476 25288
rect 3424 25245 3433 25279
rect 3433 25245 3467 25279
rect 3467 25245 3476 25279
rect 3424 25236 3476 25245
rect 4528 25100 4580 25152
rect 5540 25143 5592 25152
rect 5540 25109 5549 25143
rect 5549 25109 5583 25143
rect 5583 25109 5592 25143
rect 5540 25100 5592 25109
rect 5632 25100 5684 25152
rect 5908 25236 5960 25288
rect 6276 25304 6328 25356
rect 7288 25304 7340 25356
rect 7472 25304 7524 25356
rect 7840 25347 7892 25356
rect 7840 25313 7849 25347
rect 7849 25313 7883 25347
rect 7883 25313 7892 25347
rect 7840 25304 7892 25313
rect 9680 25304 9732 25356
rect 10048 25304 10100 25356
rect 10324 25347 10376 25356
rect 10324 25313 10333 25347
rect 10333 25313 10367 25347
rect 10367 25313 10376 25347
rect 10324 25304 10376 25313
rect 10784 25304 10836 25356
rect 11428 25372 11480 25424
rect 13544 25372 13596 25424
rect 15476 25440 15528 25492
rect 17040 25440 17092 25492
rect 15936 25372 15988 25424
rect 16764 25372 16816 25424
rect 13452 25304 13504 25356
rect 8116 25168 8168 25220
rect 9312 25279 9364 25288
rect 9312 25245 9321 25279
rect 9321 25245 9355 25279
rect 9355 25245 9364 25279
rect 9312 25236 9364 25245
rect 11060 25236 11112 25288
rect 11520 25236 11572 25288
rect 9588 25100 9640 25152
rect 10140 25143 10192 25152
rect 10140 25109 10149 25143
rect 10149 25109 10183 25143
rect 10183 25109 10192 25143
rect 10140 25100 10192 25109
rect 10876 25143 10928 25152
rect 10876 25109 10885 25143
rect 10885 25109 10919 25143
rect 10919 25109 10928 25143
rect 10876 25100 10928 25109
rect 11152 25168 11204 25220
rect 14096 25236 14148 25288
rect 14740 25304 14792 25356
rect 17592 25304 17644 25356
rect 20536 25440 20588 25492
rect 22376 25440 22428 25492
rect 23848 25440 23900 25492
rect 22468 25415 22520 25424
rect 22468 25381 22477 25415
rect 22477 25381 22511 25415
rect 22511 25381 22520 25415
rect 22468 25372 22520 25381
rect 14464 25236 14516 25288
rect 14648 25236 14700 25288
rect 18420 25236 18472 25288
rect 14004 25100 14056 25152
rect 14556 25143 14608 25152
rect 14556 25109 14565 25143
rect 14565 25109 14599 25143
rect 14599 25109 14608 25143
rect 14556 25100 14608 25109
rect 15384 25100 15436 25152
rect 18328 25100 18380 25152
rect 22008 25304 22060 25356
rect 19524 25236 19576 25288
rect 22744 25236 22796 25288
rect 19064 25100 19116 25152
rect 20628 25143 20680 25152
rect 20628 25109 20637 25143
rect 20637 25109 20671 25143
rect 20671 25109 20680 25143
rect 20628 25100 20680 25109
rect 23940 25347 23992 25356
rect 23940 25313 23949 25347
rect 23949 25313 23983 25347
rect 23983 25313 23992 25347
rect 23940 25304 23992 25313
rect 25320 25440 25372 25492
rect 25596 25440 25648 25492
rect 25688 25483 25740 25492
rect 25688 25449 25697 25483
rect 25697 25449 25731 25483
rect 25731 25449 25740 25483
rect 25688 25440 25740 25449
rect 25964 25440 26016 25492
rect 26700 25440 26752 25492
rect 27896 25440 27948 25492
rect 30748 25440 30800 25492
rect 31392 25440 31444 25492
rect 24860 25304 24912 25356
rect 25228 25347 25280 25356
rect 25228 25313 25237 25347
rect 25237 25313 25271 25347
rect 25271 25313 25280 25347
rect 25228 25304 25280 25313
rect 25504 25304 25556 25356
rect 24952 25236 25004 25288
rect 26056 25347 26108 25356
rect 26056 25313 26065 25347
rect 26065 25313 26099 25347
rect 26099 25313 26108 25347
rect 26056 25304 26108 25313
rect 29368 25304 29420 25356
rect 29736 25304 29788 25356
rect 26332 25236 26384 25288
rect 31300 25236 31352 25288
rect 33140 25236 33192 25288
rect 25412 25168 25464 25220
rect 28172 25211 28224 25220
rect 28172 25177 28181 25211
rect 28181 25177 28215 25211
rect 28215 25177 28224 25211
rect 28172 25168 28224 25177
rect 27988 25143 28040 25152
rect 27988 25109 27997 25143
rect 27997 25109 28031 25143
rect 28031 25109 28040 25143
rect 27988 25100 28040 25109
rect 29184 25100 29236 25152
rect 30380 25100 30432 25152
rect 6286 24998 6338 25050
rect 6350 24998 6402 25050
rect 6414 24998 6466 25050
rect 6478 24998 6530 25050
rect 6542 24998 6594 25050
rect 13646 24998 13698 25050
rect 13710 24998 13762 25050
rect 13774 24998 13826 25050
rect 13838 24998 13890 25050
rect 13902 24998 13954 25050
rect 21006 24998 21058 25050
rect 21070 24998 21122 25050
rect 21134 24998 21186 25050
rect 21198 24998 21250 25050
rect 21262 24998 21314 25050
rect 28366 24998 28418 25050
rect 28430 24998 28482 25050
rect 28494 24998 28546 25050
rect 28558 24998 28610 25050
rect 28622 24998 28674 25050
rect 5816 24896 5868 24948
rect 8576 24896 8628 24948
rect 9312 24939 9364 24948
rect 9312 24905 9321 24939
rect 9321 24905 9355 24939
rect 9355 24905 9364 24939
rect 9312 24896 9364 24905
rect 9404 24939 9456 24948
rect 9404 24905 9413 24939
rect 9413 24905 9447 24939
rect 9447 24905 9456 24939
rect 9404 24896 9456 24905
rect 10048 24896 10100 24948
rect 10876 24896 10928 24948
rect 11704 24939 11756 24948
rect 11704 24905 11713 24939
rect 11713 24905 11747 24939
rect 11747 24905 11756 24939
rect 11704 24896 11756 24905
rect 1308 24760 1360 24812
rect 4252 24760 4304 24812
rect 7380 24760 7432 24812
rect 3240 24735 3292 24744
rect 3240 24701 3249 24735
rect 3249 24701 3283 24735
rect 3283 24701 3292 24735
rect 3240 24692 3292 24701
rect 5540 24692 5592 24744
rect 6184 24692 6236 24744
rect 6460 24735 6512 24744
rect 6460 24701 6469 24735
rect 6469 24701 6503 24735
rect 6503 24701 6512 24735
rect 6460 24692 6512 24701
rect 7288 24735 7340 24744
rect 7288 24701 7297 24735
rect 7297 24701 7331 24735
rect 7331 24701 7340 24735
rect 7288 24692 7340 24701
rect 9588 24735 9640 24744
rect 9588 24701 9597 24735
rect 9597 24701 9631 24735
rect 9631 24701 9640 24735
rect 9588 24692 9640 24701
rect 9680 24735 9732 24744
rect 9680 24701 9689 24735
rect 9689 24701 9723 24735
rect 9723 24701 9732 24735
rect 9680 24692 9732 24701
rect 9956 24735 10008 24744
rect 9956 24701 9965 24735
rect 9965 24701 9999 24735
rect 9999 24701 10008 24735
rect 9956 24692 10008 24701
rect 10140 24692 10192 24744
rect 10692 24828 10744 24880
rect 10784 24828 10836 24880
rect 11888 24828 11940 24880
rect 3884 24624 3936 24676
rect 4620 24599 4672 24608
rect 4620 24565 4629 24599
rect 4629 24565 4663 24599
rect 4663 24565 4672 24599
rect 4620 24556 4672 24565
rect 5264 24556 5316 24608
rect 5448 24556 5500 24608
rect 5632 24556 5684 24608
rect 9128 24624 9180 24676
rect 14280 24896 14332 24948
rect 14556 24896 14608 24948
rect 14924 24896 14976 24948
rect 15568 24939 15620 24948
rect 15568 24905 15577 24939
rect 15577 24905 15611 24939
rect 15611 24905 15620 24939
rect 15568 24896 15620 24905
rect 16304 24896 16356 24948
rect 10784 24735 10836 24744
rect 10784 24701 10793 24735
rect 10793 24701 10827 24735
rect 10827 24701 10836 24735
rect 10784 24692 10836 24701
rect 10968 24735 11020 24744
rect 10968 24701 10977 24735
rect 10977 24701 11011 24735
rect 11011 24701 11020 24735
rect 10968 24692 11020 24701
rect 11428 24692 11480 24744
rect 11520 24735 11572 24744
rect 11520 24701 11529 24735
rect 11529 24701 11563 24735
rect 11563 24701 11572 24735
rect 11520 24692 11572 24701
rect 11060 24624 11112 24676
rect 11888 24735 11940 24744
rect 11888 24701 11897 24735
rect 11897 24701 11931 24735
rect 11931 24701 11940 24735
rect 11888 24692 11940 24701
rect 13268 24760 13320 24812
rect 14464 24828 14516 24880
rect 15108 24828 15160 24880
rect 14096 24760 14148 24812
rect 18512 24896 18564 24948
rect 19524 24939 19576 24948
rect 19524 24905 19533 24939
rect 19533 24905 19567 24939
rect 19567 24905 19576 24939
rect 19524 24896 19576 24905
rect 18972 24828 19024 24880
rect 19064 24828 19116 24880
rect 27896 24896 27948 24948
rect 27988 24896 28040 24948
rect 28172 24939 28224 24948
rect 28172 24905 28181 24939
rect 28181 24905 28215 24939
rect 28215 24905 28224 24939
rect 28172 24896 28224 24905
rect 29736 24896 29788 24948
rect 23480 24828 23532 24880
rect 25504 24828 25556 24880
rect 17132 24760 17184 24812
rect 19616 24760 19668 24812
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 12256 24624 12308 24676
rect 10600 24599 10652 24608
rect 10600 24565 10609 24599
rect 10609 24565 10643 24599
rect 10643 24565 10652 24599
rect 10600 24556 10652 24565
rect 11244 24599 11296 24608
rect 11244 24565 11253 24599
rect 11253 24565 11287 24599
rect 11287 24565 11296 24599
rect 11244 24556 11296 24565
rect 11796 24556 11848 24608
rect 13912 24692 13964 24744
rect 14004 24692 14056 24744
rect 16488 24692 16540 24744
rect 19064 24692 19116 24744
rect 20628 24692 20680 24744
rect 21456 24692 21508 24744
rect 22652 24692 22704 24744
rect 22744 24692 22796 24744
rect 27712 24803 27764 24812
rect 27712 24769 27721 24803
rect 27721 24769 27755 24803
rect 27755 24769 27764 24803
rect 27712 24760 27764 24769
rect 28264 24803 28316 24812
rect 28264 24769 28273 24803
rect 28273 24769 28307 24803
rect 28307 24769 28316 24803
rect 28264 24760 28316 24769
rect 12992 24624 13044 24676
rect 14832 24556 14884 24608
rect 16120 24556 16172 24608
rect 16212 24599 16264 24608
rect 16212 24565 16221 24599
rect 16221 24565 16255 24599
rect 16255 24565 16264 24599
rect 16212 24556 16264 24565
rect 17132 24599 17184 24608
rect 17132 24565 17141 24599
rect 17141 24565 17175 24599
rect 17175 24565 17184 24599
rect 17132 24556 17184 24565
rect 17500 24599 17552 24608
rect 17500 24565 17509 24599
rect 17509 24565 17543 24599
rect 17543 24565 17552 24599
rect 17500 24556 17552 24565
rect 17960 24667 18012 24676
rect 17960 24633 17969 24667
rect 17969 24633 18003 24667
rect 18003 24633 18012 24667
rect 17960 24624 18012 24633
rect 19340 24556 19392 24608
rect 22836 24556 22888 24608
rect 24676 24556 24728 24608
rect 25780 24556 25832 24608
rect 27896 24735 27948 24744
rect 27896 24701 27905 24735
rect 27905 24701 27939 24735
rect 27939 24701 27948 24735
rect 27896 24692 27948 24701
rect 27988 24735 28040 24744
rect 27988 24701 27997 24735
rect 27997 24701 28031 24735
rect 28031 24701 28040 24735
rect 27988 24692 28040 24701
rect 30288 24735 30340 24744
rect 30288 24701 30297 24735
rect 30297 24701 30331 24735
rect 30331 24701 30340 24735
rect 30288 24692 30340 24701
rect 29184 24556 29236 24608
rect 6946 24454 6998 24506
rect 7010 24454 7062 24506
rect 7074 24454 7126 24506
rect 7138 24454 7190 24506
rect 7202 24454 7254 24506
rect 14306 24454 14358 24506
rect 14370 24454 14422 24506
rect 14434 24454 14486 24506
rect 14498 24454 14550 24506
rect 14562 24454 14614 24506
rect 21666 24454 21718 24506
rect 21730 24454 21782 24506
rect 21794 24454 21846 24506
rect 21858 24454 21910 24506
rect 21922 24454 21974 24506
rect 29026 24454 29078 24506
rect 29090 24454 29142 24506
rect 29154 24454 29206 24506
rect 29218 24454 29270 24506
rect 29282 24454 29334 24506
rect 3424 24395 3476 24404
rect 3424 24361 3433 24395
rect 3433 24361 3467 24395
rect 3467 24361 3476 24395
rect 3424 24352 3476 24361
rect 3884 24395 3936 24404
rect 3884 24361 3893 24395
rect 3893 24361 3927 24395
rect 3927 24361 3936 24395
rect 3884 24352 3936 24361
rect 4620 24352 4672 24404
rect 6460 24352 6512 24404
rect 7288 24352 7340 24404
rect 7748 24352 7800 24404
rect 8944 24352 8996 24404
rect 3240 24216 3292 24268
rect 4252 24259 4304 24268
rect 4252 24225 4261 24259
rect 4261 24225 4295 24259
rect 4295 24225 4304 24259
rect 4252 24216 4304 24225
rect 5632 24216 5684 24268
rect 4252 24080 4304 24132
rect 9128 24327 9180 24336
rect 9128 24293 9137 24327
rect 9137 24293 9171 24327
rect 9171 24293 9180 24327
rect 9128 24284 9180 24293
rect 7656 24216 7708 24268
rect 9036 24259 9088 24268
rect 9036 24225 9045 24259
rect 9045 24225 9079 24259
rect 9079 24225 9088 24259
rect 9036 24216 9088 24225
rect 10692 24352 10744 24404
rect 10784 24352 10836 24404
rect 12440 24352 12492 24404
rect 13360 24352 13412 24404
rect 21732 24352 21784 24404
rect 22652 24395 22704 24404
rect 22652 24361 22661 24395
rect 22661 24361 22695 24395
rect 22695 24361 22704 24395
rect 22652 24352 22704 24361
rect 26700 24352 26752 24404
rect 10600 24284 10652 24336
rect 13268 24284 13320 24336
rect 14372 24327 14424 24336
rect 14372 24293 14381 24327
rect 14381 24293 14415 24327
rect 14415 24293 14424 24327
rect 14372 24284 14424 24293
rect 14740 24327 14792 24336
rect 14740 24293 14749 24327
rect 14749 24293 14783 24327
rect 14783 24293 14792 24327
rect 14740 24284 14792 24293
rect 18144 24327 18196 24336
rect 18144 24293 18153 24327
rect 18153 24293 18187 24327
rect 18187 24293 18196 24327
rect 18144 24284 18196 24293
rect 19064 24327 19116 24336
rect 19064 24293 19073 24327
rect 19073 24293 19107 24327
rect 19107 24293 19116 24327
rect 19064 24284 19116 24293
rect 20076 24284 20128 24336
rect 11152 24259 11204 24268
rect 11152 24225 11161 24259
rect 11161 24225 11195 24259
rect 11195 24225 11204 24259
rect 11152 24216 11204 24225
rect 11244 24216 11296 24268
rect 11520 24216 11572 24268
rect 12624 24216 12676 24268
rect 15844 24216 15896 24268
rect 10784 24148 10836 24200
rect 13912 24148 13964 24200
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 5908 24012 5960 24064
rect 8760 24055 8812 24064
rect 8760 24021 8769 24055
rect 8769 24021 8803 24055
rect 8803 24021 8812 24055
rect 8760 24012 8812 24021
rect 11520 24012 11572 24064
rect 12256 24055 12308 24064
rect 12256 24021 12265 24055
rect 12265 24021 12299 24055
rect 12299 24021 12308 24055
rect 12256 24012 12308 24021
rect 16028 24080 16080 24132
rect 17132 24216 17184 24268
rect 14924 24012 14976 24064
rect 15292 24012 15344 24064
rect 16212 24012 16264 24064
rect 16948 24012 17000 24064
rect 17500 24148 17552 24200
rect 18880 24259 18932 24268
rect 18880 24225 18889 24259
rect 18889 24225 18923 24259
rect 18923 24225 18932 24259
rect 18880 24216 18932 24225
rect 19156 24259 19208 24268
rect 19156 24225 19165 24259
rect 19165 24225 19199 24259
rect 19199 24225 19208 24259
rect 19156 24216 19208 24225
rect 19432 24148 19484 24200
rect 17960 24080 18012 24132
rect 18880 24012 18932 24064
rect 21456 24012 21508 24064
rect 24124 24216 24176 24268
rect 25136 24259 25188 24268
rect 25136 24225 25153 24259
rect 25153 24225 25187 24259
rect 25187 24225 25188 24259
rect 25136 24216 25188 24225
rect 25412 24259 25464 24268
rect 25412 24225 25421 24259
rect 25421 24225 25455 24259
rect 25455 24225 25464 24259
rect 25412 24216 25464 24225
rect 25596 24259 25648 24268
rect 25596 24225 25605 24259
rect 25605 24225 25639 24259
rect 25639 24225 25648 24259
rect 25596 24216 25648 24225
rect 25872 24216 25924 24268
rect 26240 24259 26292 24268
rect 26240 24225 26249 24259
rect 26249 24225 26283 24259
rect 26283 24225 26292 24259
rect 26240 24216 26292 24225
rect 22192 24191 22244 24200
rect 22192 24157 22201 24191
rect 22201 24157 22235 24191
rect 22235 24157 22244 24191
rect 22192 24148 22244 24157
rect 24308 24191 24360 24200
rect 24308 24157 24317 24191
rect 24317 24157 24351 24191
rect 24351 24157 24360 24191
rect 24308 24148 24360 24157
rect 26608 24259 26660 24268
rect 26608 24225 26617 24259
rect 26617 24225 26651 24259
rect 26651 24225 26660 24259
rect 26608 24216 26660 24225
rect 27896 24284 27948 24336
rect 24216 24080 24268 24132
rect 30380 24148 30432 24200
rect 31576 24191 31628 24200
rect 31576 24157 31585 24191
rect 31585 24157 31619 24191
rect 31619 24157 31628 24191
rect 31576 24148 31628 24157
rect 33140 24148 33192 24200
rect 29460 24080 29512 24132
rect 22100 24012 22152 24064
rect 23940 24012 23992 24064
rect 24860 24055 24912 24064
rect 24860 24021 24869 24055
rect 24869 24021 24903 24055
rect 24903 24021 24912 24055
rect 24860 24012 24912 24021
rect 24952 24012 25004 24064
rect 25136 24012 25188 24064
rect 28080 24012 28132 24064
rect 6286 23910 6338 23962
rect 6350 23910 6402 23962
rect 6414 23910 6466 23962
rect 6478 23910 6530 23962
rect 6542 23910 6594 23962
rect 13646 23910 13698 23962
rect 13710 23910 13762 23962
rect 13774 23910 13826 23962
rect 13838 23910 13890 23962
rect 13902 23910 13954 23962
rect 21006 23910 21058 23962
rect 21070 23910 21122 23962
rect 21134 23910 21186 23962
rect 21198 23910 21250 23962
rect 21262 23910 21314 23962
rect 28366 23910 28418 23962
rect 28430 23910 28482 23962
rect 28494 23910 28546 23962
rect 28558 23910 28610 23962
rect 28622 23910 28674 23962
rect 3240 23808 3292 23860
rect 4160 23808 4212 23860
rect 4528 23672 4580 23724
rect 5724 23672 5776 23724
rect 7748 23808 7800 23860
rect 7840 23808 7892 23860
rect 11060 23808 11112 23860
rect 11152 23808 11204 23860
rect 11336 23808 11388 23860
rect 11428 23808 11480 23860
rect 12992 23851 13044 23860
rect 12992 23817 13001 23851
rect 13001 23817 13035 23851
rect 13035 23817 13044 23851
rect 12992 23808 13044 23817
rect 14004 23851 14056 23860
rect 14004 23817 14013 23851
rect 14013 23817 14047 23851
rect 14047 23817 14056 23851
rect 14004 23808 14056 23817
rect 14372 23808 14424 23860
rect 15844 23808 15896 23860
rect 17868 23808 17920 23860
rect 18328 23851 18380 23860
rect 18328 23817 18337 23851
rect 18337 23817 18371 23851
rect 18371 23817 18380 23851
rect 18328 23808 18380 23817
rect 18420 23851 18472 23860
rect 18420 23817 18429 23851
rect 18429 23817 18463 23851
rect 18463 23817 18472 23851
rect 18420 23808 18472 23817
rect 25320 23808 25372 23860
rect 13912 23740 13964 23792
rect 6552 23604 6604 23656
rect 7748 23604 7800 23656
rect 8392 23715 8444 23724
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 8760 23672 8812 23724
rect 11336 23672 11388 23724
rect 12256 23672 12308 23724
rect 15200 23740 15252 23792
rect 15660 23740 15712 23792
rect 11980 23604 12032 23656
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 14832 23672 14884 23724
rect 7656 23536 7708 23588
rect 8116 23579 8168 23588
rect 8116 23545 8125 23579
rect 8125 23545 8159 23579
rect 8159 23545 8168 23579
rect 8116 23536 8168 23545
rect 11888 23536 11940 23588
rect 14648 23604 14700 23656
rect 15384 23604 15436 23656
rect 16120 23604 16172 23656
rect 22284 23672 22336 23724
rect 23112 23672 23164 23724
rect 25504 23672 25556 23724
rect 25688 23672 25740 23724
rect 17592 23647 17644 23656
rect 17592 23613 17601 23647
rect 17601 23613 17635 23647
rect 17635 23613 17644 23647
rect 17592 23604 17644 23613
rect 5172 23468 5224 23520
rect 5540 23468 5592 23520
rect 6460 23511 6512 23520
rect 6460 23477 6469 23511
rect 6469 23477 6503 23511
rect 6503 23477 6512 23511
rect 6460 23468 6512 23477
rect 7748 23511 7800 23520
rect 7748 23477 7757 23511
rect 7757 23477 7791 23511
rect 7791 23477 7800 23511
rect 7748 23468 7800 23477
rect 10692 23468 10744 23520
rect 13452 23468 13504 23520
rect 14464 23536 14516 23588
rect 15752 23536 15804 23588
rect 18696 23647 18748 23656
rect 18696 23613 18705 23647
rect 18705 23613 18739 23647
rect 18739 23613 18748 23647
rect 18696 23604 18748 23613
rect 19708 23647 19760 23656
rect 19708 23613 19717 23647
rect 19717 23613 19751 23647
rect 19751 23613 19760 23647
rect 19708 23604 19760 23613
rect 20904 23604 20956 23656
rect 21732 23604 21784 23656
rect 22100 23604 22152 23656
rect 26700 23808 26752 23860
rect 26424 23783 26476 23792
rect 26424 23749 26433 23783
rect 26433 23749 26467 23783
rect 26467 23749 26476 23783
rect 26424 23740 26476 23749
rect 27988 23808 28040 23860
rect 20536 23536 20588 23588
rect 23388 23536 23440 23588
rect 24952 23536 25004 23588
rect 25136 23536 25188 23588
rect 14648 23468 14700 23520
rect 15476 23468 15528 23520
rect 15568 23468 15620 23520
rect 16028 23468 16080 23520
rect 17040 23468 17092 23520
rect 18328 23468 18380 23520
rect 18880 23511 18932 23520
rect 18880 23477 18889 23511
rect 18889 23477 18923 23511
rect 18923 23477 18932 23511
rect 18880 23468 18932 23477
rect 19064 23511 19116 23520
rect 19064 23477 19073 23511
rect 19073 23477 19107 23511
rect 19107 23477 19116 23511
rect 19064 23468 19116 23477
rect 20352 23511 20404 23520
rect 20352 23477 20361 23511
rect 20361 23477 20395 23511
rect 20395 23477 20404 23511
rect 20352 23468 20404 23477
rect 20996 23511 21048 23520
rect 20996 23477 21005 23511
rect 21005 23477 21039 23511
rect 21039 23477 21048 23511
rect 20996 23468 21048 23477
rect 23480 23468 23532 23520
rect 24400 23468 24452 23520
rect 24860 23468 24912 23520
rect 25780 23468 25832 23520
rect 26332 23647 26384 23656
rect 26332 23613 26341 23647
rect 26341 23613 26375 23647
rect 26375 23613 26384 23647
rect 26332 23604 26384 23613
rect 26424 23647 26476 23656
rect 26424 23613 26433 23647
rect 26433 23613 26467 23647
rect 26467 23613 26476 23647
rect 26424 23604 26476 23613
rect 26700 23647 26752 23656
rect 26700 23613 26709 23647
rect 26709 23613 26743 23647
rect 26743 23613 26752 23647
rect 26700 23604 26752 23613
rect 26884 23647 26936 23656
rect 26884 23613 26893 23647
rect 26893 23613 26927 23647
rect 26927 23613 26936 23647
rect 26884 23604 26936 23613
rect 29644 23740 29696 23792
rect 27804 23647 27856 23656
rect 27804 23613 27813 23647
rect 27813 23613 27847 23647
rect 27847 23613 27856 23647
rect 27804 23604 27856 23613
rect 28816 23604 28868 23656
rect 27988 23536 28040 23588
rect 26056 23468 26108 23520
rect 27344 23468 27396 23520
rect 29368 23511 29420 23520
rect 29368 23477 29377 23511
rect 29377 23477 29411 23511
rect 29411 23477 29420 23511
rect 29368 23468 29420 23477
rect 6946 23366 6998 23418
rect 7010 23366 7062 23418
rect 7074 23366 7126 23418
rect 7138 23366 7190 23418
rect 7202 23366 7254 23418
rect 14306 23366 14358 23418
rect 14370 23366 14422 23418
rect 14434 23366 14486 23418
rect 14498 23366 14550 23418
rect 14562 23366 14614 23418
rect 21666 23366 21718 23418
rect 21730 23366 21782 23418
rect 21794 23366 21846 23418
rect 21858 23366 21910 23418
rect 21922 23366 21974 23418
rect 29026 23366 29078 23418
rect 29090 23366 29142 23418
rect 29154 23366 29206 23418
rect 29218 23366 29270 23418
rect 29282 23366 29334 23418
rect 4160 23264 4212 23316
rect 4436 23264 4488 23316
rect 5264 23264 5316 23316
rect 4988 23196 5040 23248
rect 5540 23196 5592 23248
rect 6460 23264 6512 23316
rect 6552 23307 6604 23316
rect 6552 23273 6561 23307
rect 6561 23273 6595 23307
rect 6595 23273 6604 23307
rect 6552 23264 6604 23273
rect 9680 23264 9732 23316
rect 11060 23264 11112 23316
rect 7104 23196 7156 23248
rect 8208 23196 8260 23248
rect 11336 23239 11388 23248
rect 11336 23205 11345 23239
rect 11345 23205 11379 23239
rect 11379 23205 11388 23239
rect 11336 23196 11388 23205
rect 5724 23171 5776 23180
rect 5724 23137 5733 23171
rect 5733 23137 5767 23171
rect 5767 23137 5776 23171
rect 5724 23128 5776 23137
rect 7748 23171 7800 23180
rect 7748 23137 7757 23171
rect 7757 23137 7791 23171
rect 7791 23137 7800 23171
rect 7748 23128 7800 23137
rect 13544 23264 13596 23316
rect 14740 23264 14792 23316
rect 17592 23307 17644 23316
rect 17592 23273 17601 23307
rect 17601 23273 17635 23307
rect 17635 23273 17644 23307
rect 17592 23264 17644 23273
rect 18696 23264 18748 23316
rect 25228 23307 25280 23316
rect 25228 23273 25237 23307
rect 25237 23273 25271 23307
rect 25271 23273 25280 23307
rect 25228 23264 25280 23273
rect 25596 23264 25648 23316
rect 26240 23264 26292 23316
rect 14096 23196 14148 23248
rect 15292 23196 15344 23248
rect 15844 23196 15896 23248
rect 19340 23196 19392 23248
rect 20352 23196 20404 23248
rect 20996 23239 21048 23248
rect 20996 23205 21005 23239
rect 21005 23205 21039 23239
rect 21039 23205 21048 23239
rect 20996 23196 21048 23205
rect 21456 23196 21508 23248
rect 13544 23171 13596 23180
rect 13544 23137 13553 23171
rect 13553 23137 13587 23171
rect 13587 23137 13596 23171
rect 13544 23128 13596 23137
rect 5908 23103 5960 23112
rect 5908 23069 5917 23103
rect 5917 23069 5951 23103
rect 5951 23069 5960 23103
rect 5908 23060 5960 23069
rect 6736 23060 6788 23112
rect 8392 23060 8444 23112
rect 8668 23103 8720 23112
rect 8668 23069 8677 23103
rect 8677 23069 8711 23103
rect 8711 23069 8720 23103
rect 8668 23060 8720 23069
rect 10968 23060 11020 23112
rect 12532 23060 12584 23112
rect 12624 23103 12676 23112
rect 12624 23069 12633 23103
rect 12633 23069 12667 23103
rect 12667 23069 12676 23103
rect 14280 23128 14332 23180
rect 14372 23171 14424 23180
rect 14372 23137 14401 23171
rect 14401 23137 14424 23171
rect 14372 23128 14424 23137
rect 12624 23060 12676 23069
rect 8116 22992 8168 23044
rect 13268 22992 13320 23044
rect 13452 22992 13504 23044
rect 14924 23128 14976 23180
rect 17868 23128 17920 23180
rect 25504 23196 25556 23248
rect 14740 22992 14792 23044
rect 15752 23060 15804 23112
rect 16120 23103 16172 23112
rect 16120 23069 16129 23103
rect 16129 23069 16163 23103
rect 16163 23069 16172 23103
rect 16120 23060 16172 23069
rect 18052 23060 18104 23112
rect 18972 23060 19024 23112
rect 22100 23060 22152 23112
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 23112 23103 23164 23112
rect 23112 23069 23121 23103
rect 23121 23069 23155 23103
rect 23155 23069 23164 23103
rect 23112 23060 23164 23069
rect 24032 23103 24084 23112
rect 24032 23069 24041 23103
rect 24041 23069 24075 23103
rect 24075 23069 24084 23103
rect 24032 23060 24084 23069
rect 24676 23171 24728 23180
rect 24676 23137 24685 23171
rect 24685 23137 24719 23171
rect 24719 23137 24728 23171
rect 24676 23128 24728 23137
rect 26056 23196 26108 23248
rect 25872 23128 25924 23180
rect 24768 22992 24820 23044
rect 24952 23060 25004 23112
rect 26608 23128 26660 23180
rect 26700 23171 26752 23180
rect 26700 23137 26709 23171
rect 26709 23137 26743 23171
rect 26743 23137 26752 23171
rect 26700 23128 26752 23137
rect 26884 23128 26936 23180
rect 27528 23060 27580 23112
rect 30380 23307 30432 23316
rect 30380 23273 30389 23307
rect 30389 23273 30423 23307
rect 30423 23273 30432 23307
rect 30380 23264 30432 23273
rect 29920 23196 29972 23248
rect 28264 23128 28316 23180
rect 31300 23171 31352 23180
rect 31300 23137 31309 23171
rect 31309 23137 31343 23171
rect 31343 23137 31352 23171
rect 31300 23128 31352 23137
rect 25964 22992 26016 23044
rect 26240 23035 26292 23044
rect 26240 23001 26249 23035
rect 26249 23001 26283 23035
rect 26283 23001 26292 23035
rect 26240 22992 26292 23001
rect 26332 22992 26384 23044
rect 26792 22992 26844 23044
rect 28908 23103 28960 23112
rect 28908 23069 28917 23103
rect 28917 23069 28951 23103
rect 28951 23069 28960 23103
rect 28908 23060 28960 23069
rect 30288 23060 30340 23112
rect 5632 22924 5684 22976
rect 7196 22967 7248 22976
rect 7196 22933 7205 22967
rect 7205 22933 7239 22967
rect 7239 22933 7248 22967
rect 7196 22924 7248 22933
rect 7656 22924 7708 22976
rect 13544 22924 13596 22976
rect 14280 22924 14332 22976
rect 14832 22924 14884 22976
rect 15384 22924 15436 22976
rect 18880 22924 18932 22976
rect 21364 22967 21416 22976
rect 21364 22933 21373 22967
rect 21373 22933 21407 22967
rect 21407 22933 21416 22967
rect 21364 22924 21416 22933
rect 23204 22924 23256 22976
rect 24860 22924 24912 22976
rect 25780 22924 25832 22976
rect 28724 22924 28776 22976
rect 31300 22924 31352 22976
rect 6286 22822 6338 22874
rect 6350 22822 6402 22874
rect 6414 22822 6466 22874
rect 6478 22822 6530 22874
rect 6542 22822 6594 22874
rect 13646 22822 13698 22874
rect 13710 22822 13762 22874
rect 13774 22822 13826 22874
rect 13838 22822 13890 22874
rect 13902 22822 13954 22874
rect 21006 22822 21058 22874
rect 21070 22822 21122 22874
rect 21134 22822 21186 22874
rect 21198 22822 21250 22874
rect 21262 22822 21314 22874
rect 28366 22822 28418 22874
rect 28430 22822 28482 22874
rect 28494 22822 28546 22874
rect 28558 22822 28610 22874
rect 28622 22822 28674 22874
rect 4988 22720 5040 22772
rect 5724 22720 5776 22772
rect 1308 22448 1360 22500
rect 5172 22559 5224 22568
rect 5172 22525 5181 22559
rect 5181 22525 5215 22559
rect 5215 22525 5224 22559
rect 5172 22516 5224 22525
rect 6092 22559 6144 22568
rect 6092 22525 6101 22559
rect 6101 22525 6135 22559
rect 6135 22525 6144 22559
rect 6092 22516 6144 22525
rect 7196 22720 7248 22772
rect 8668 22720 8720 22772
rect 14188 22720 14240 22772
rect 14464 22763 14516 22772
rect 14464 22729 14473 22763
rect 14473 22729 14507 22763
rect 14507 22729 14516 22763
rect 14464 22720 14516 22729
rect 14740 22763 14792 22772
rect 14740 22729 14749 22763
rect 14749 22729 14783 22763
rect 14783 22729 14792 22763
rect 14740 22720 14792 22729
rect 14372 22652 14424 22704
rect 15016 22652 15068 22704
rect 7104 22627 7156 22636
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 7104 22584 7156 22593
rect 8392 22584 8444 22636
rect 12440 22584 12492 22636
rect 6644 22448 6696 22500
rect 9772 22559 9824 22568
rect 9772 22525 9781 22559
rect 9781 22525 9815 22559
rect 9815 22525 9824 22559
rect 9772 22516 9824 22525
rect 5448 22423 5500 22432
rect 5448 22389 5457 22423
rect 5457 22389 5491 22423
rect 5491 22389 5500 22423
rect 5448 22380 5500 22389
rect 6276 22423 6328 22432
rect 6276 22389 6285 22423
rect 6285 22389 6319 22423
rect 6319 22389 6328 22423
rect 6276 22380 6328 22389
rect 6552 22423 6604 22432
rect 6552 22389 6561 22423
rect 6561 22389 6595 22423
rect 6595 22389 6604 22423
rect 6552 22380 6604 22389
rect 6828 22380 6880 22432
rect 7656 22380 7708 22432
rect 11612 22559 11664 22568
rect 11612 22525 11621 22559
rect 11621 22525 11655 22559
rect 11655 22525 11664 22559
rect 11612 22516 11664 22525
rect 11704 22516 11756 22568
rect 12808 22559 12860 22568
rect 12808 22525 12817 22559
rect 12817 22525 12851 22559
rect 12851 22525 12860 22559
rect 12808 22516 12860 22525
rect 13360 22516 13412 22568
rect 12624 22448 12676 22500
rect 14556 22516 14608 22568
rect 14740 22559 14792 22568
rect 14740 22525 14749 22559
rect 14749 22525 14783 22559
rect 14783 22525 14792 22559
rect 14740 22516 14792 22525
rect 15108 22516 15160 22568
rect 15844 22695 15896 22704
rect 15844 22661 15853 22695
rect 15853 22661 15887 22695
rect 15887 22661 15896 22695
rect 15844 22652 15896 22661
rect 16120 22720 16172 22772
rect 17040 22720 17092 22772
rect 15568 22516 15620 22568
rect 15476 22448 15528 22500
rect 10140 22380 10192 22432
rect 10784 22423 10836 22432
rect 10784 22389 10793 22423
rect 10793 22389 10827 22423
rect 10827 22389 10836 22423
rect 10784 22380 10836 22389
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 11980 22423 12032 22432
rect 11980 22389 11989 22423
rect 11989 22389 12023 22423
rect 12023 22389 12032 22423
rect 11980 22380 12032 22389
rect 12532 22380 12584 22432
rect 13268 22380 13320 22432
rect 13452 22423 13504 22432
rect 13452 22389 13461 22423
rect 13461 22389 13495 22423
rect 13495 22389 13504 22423
rect 13452 22380 13504 22389
rect 14188 22380 14240 22432
rect 14648 22380 14700 22432
rect 15844 22380 15896 22432
rect 20904 22763 20956 22772
rect 20904 22729 20913 22763
rect 20913 22729 20947 22763
rect 20947 22729 20956 22763
rect 20904 22720 20956 22729
rect 21364 22720 21416 22772
rect 22192 22720 22244 22772
rect 23204 22720 23256 22772
rect 24308 22763 24360 22772
rect 24308 22729 24317 22763
rect 24317 22729 24351 22763
rect 24351 22729 24360 22763
rect 24308 22720 24360 22729
rect 24676 22720 24728 22772
rect 26056 22720 26108 22772
rect 28908 22720 28960 22772
rect 29368 22720 29420 22772
rect 29920 22720 29972 22772
rect 19156 22652 19208 22704
rect 19064 22516 19116 22568
rect 20536 22516 20588 22568
rect 20720 22559 20772 22568
rect 20720 22525 20729 22559
rect 20729 22525 20763 22559
rect 20763 22525 20772 22559
rect 20720 22516 20772 22525
rect 21640 22652 21692 22704
rect 21456 22627 21508 22636
rect 21456 22593 21465 22627
rect 21465 22593 21499 22627
rect 21499 22593 21508 22627
rect 21456 22584 21508 22593
rect 22100 22516 22152 22568
rect 24400 22559 24452 22568
rect 24400 22525 24409 22559
rect 24409 22525 24443 22559
rect 24443 22525 24452 22559
rect 24400 22516 24452 22525
rect 25412 22559 25464 22568
rect 25412 22525 25416 22559
rect 25416 22525 25450 22559
rect 25450 22525 25464 22559
rect 25412 22516 25464 22525
rect 27896 22652 27948 22704
rect 28816 22652 28868 22704
rect 25688 22516 25740 22568
rect 17960 22448 18012 22500
rect 19340 22448 19392 22500
rect 19708 22380 19760 22432
rect 19800 22423 19852 22432
rect 19800 22389 19809 22423
rect 19809 22389 19843 22423
rect 19843 22389 19852 22423
rect 19800 22380 19852 22389
rect 20076 22423 20128 22432
rect 20076 22389 20085 22423
rect 20085 22389 20119 22423
rect 20119 22389 20128 22423
rect 20076 22380 20128 22389
rect 22192 22448 22244 22500
rect 23480 22448 23532 22500
rect 21364 22423 21416 22432
rect 21364 22389 21373 22423
rect 21373 22389 21407 22423
rect 21407 22389 21416 22423
rect 21364 22380 21416 22389
rect 25228 22423 25280 22432
rect 25228 22389 25237 22423
rect 25237 22389 25271 22423
rect 25271 22389 25280 22423
rect 25228 22380 25280 22389
rect 26056 22559 26108 22568
rect 26056 22525 26065 22559
rect 26065 22525 26099 22559
rect 26099 22525 26108 22559
rect 26056 22516 26108 22525
rect 26424 22516 26476 22568
rect 26792 22559 26844 22568
rect 26792 22525 26801 22559
rect 26801 22525 26835 22559
rect 26835 22525 26844 22559
rect 26792 22516 26844 22525
rect 26332 22448 26384 22500
rect 27528 22516 27580 22568
rect 27620 22559 27672 22568
rect 27620 22525 27629 22559
rect 27629 22525 27663 22559
rect 27663 22525 27672 22559
rect 27620 22516 27672 22525
rect 27712 22559 27764 22568
rect 27712 22525 27721 22559
rect 27721 22525 27755 22559
rect 27755 22525 27764 22559
rect 27712 22516 27764 22525
rect 27896 22559 27948 22568
rect 27896 22525 27905 22559
rect 27905 22525 27939 22559
rect 27939 22525 27948 22559
rect 27896 22516 27948 22525
rect 29460 22516 29512 22568
rect 30288 22584 30340 22636
rect 29736 22448 29788 22500
rect 27160 22380 27212 22432
rect 27252 22423 27304 22432
rect 27252 22389 27261 22423
rect 27261 22389 27295 22423
rect 27295 22389 27304 22423
rect 27252 22380 27304 22389
rect 27528 22380 27580 22432
rect 27804 22423 27856 22432
rect 27804 22389 27813 22423
rect 27813 22389 27847 22423
rect 27847 22389 27856 22423
rect 27804 22380 27856 22389
rect 6946 22278 6998 22330
rect 7010 22278 7062 22330
rect 7074 22278 7126 22330
rect 7138 22278 7190 22330
rect 7202 22278 7254 22330
rect 14306 22278 14358 22330
rect 14370 22278 14422 22330
rect 14434 22278 14486 22330
rect 14498 22278 14550 22330
rect 14562 22278 14614 22330
rect 21666 22278 21718 22330
rect 21730 22278 21782 22330
rect 21794 22278 21846 22330
rect 21858 22278 21910 22330
rect 21922 22278 21974 22330
rect 29026 22278 29078 22330
rect 29090 22278 29142 22330
rect 29154 22278 29206 22330
rect 29218 22278 29270 22330
rect 29282 22278 29334 22330
rect 5448 22176 5500 22228
rect 6276 22176 6328 22228
rect 6552 22176 6604 22228
rect 6644 22176 6696 22228
rect 9772 22176 9824 22228
rect 10416 22176 10468 22228
rect 11060 22176 11112 22228
rect 11980 22176 12032 22228
rect 13360 22176 13412 22228
rect 13452 22219 13504 22228
rect 13452 22185 13461 22219
rect 13461 22185 13495 22219
rect 13495 22185 13504 22219
rect 13452 22176 13504 22185
rect 13544 22219 13596 22228
rect 13544 22185 13553 22219
rect 13553 22185 13587 22219
rect 13587 22185 13596 22219
rect 13544 22176 13596 22185
rect 7472 22040 7524 22092
rect 3240 21972 3292 22024
rect 6092 22015 6144 22024
rect 6092 21981 6101 22015
rect 6101 21981 6135 22015
rect 6135 21981 6144 22015
rect 6092 21972 6144 21981
rect 6460 21972 6512 22024
rect 11796 22108 11848 22160
rect 14648 22108 14700 22160
rect 4160 21879 4212 21888
rect 4160 21845 4169 21879
rect 4169 21845 4203 21879
rect 4203 21845 4212 21879
rect 4160 21836 4212 21845
rect 6000 21879 6052 21888
rect 6000 21845 6009 21879
rect 6009 21845 6043 21879
rect 6043 21845 6052 21879
rect 6000 21836 6052 21845
rect 7104 21836 7156 21888
rect 8116 21972 8168 22024
rect 8208 21972 8260 22024
rect 8484 21972 8536 22024
rect 10232 21972 10284 22024
rect 10876 21972 10928 22024
rect 9588 21904 9640 21956
rect 11980 21972 12032 22024
rect 14924 22040 14976 22092
rect 15200 22040 15252 22092
rect 15568 22176 15620 22228
rect 16488 22176 16540 22228
rect 17960 22219 18012 22228
rect 17960 22185 17969 22219
rect 17969 22185 18003 22219
rect 18003 22185 18012 22219
rect 17960 22176 18012 22185
rect 20076 22176 20128 22228
rect 21364 22176 21416 22228
rect 24032 22176 24084 22228
rect 24216 22176 24268 22228
rect 25412 22176 25464 22228
rect 18236 22108 18288 22160
rect 19800 22108 19852 22160
rect 21548 22108 21600 22160
rect 23572 22108 23624 22160
rect 24584 22108 24636 22160
rect 24676 22108 24728 22160
rect 15384 22040 15436 22092
rect 15568 21972 15620 22024
rect 15752 21972 15804 22024
rect 16120 22015 16172 22024
rect 16120 21981 16129 22015
rect 16129 21981 16163 22015
rect 16163 21981 16172 22015
rect 16120 21972 16172 21981
rect 18788 21972 18840 22024
rect 18972 21972 19024 22024
rect 14648 21904 14700 21956
rect 7932 21836 7984 21888
rect 9680 21836 9732 21888
rect 9956 21879 10008 21888
rect 9956 21845 9965 21879
rect 9965 21845 9999 21879
rect 9999 21845 10008 21879
rect 9956 21836 10008 21845
rect 10048 21836 10100 21888
rect 12900 21879 12952 21888
rect 12900 21845 12909 21879
rect 12909 21845 12943 21879
rect 12943 21845 12952 21879
rect 12900 21836 12952 21845
rect 14004 21879 14056 21888
rect 14004 21845 14013 21879
rect 14013 21845 14047 21879
rect 14047 21845 14056 21879
rect 14004 21836 14056 21845
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 14924 21879 14976 21888
rect 14924 21845 14933 21879
rect 14933 21845 14967 21879
rect 14967 21845 14976 21879
rect 14924 21836 14976 21845
rect 15292 21836 15344 21888
rect 18052 21904 18104 21956
rect 17960 21836 18012 21888
rect 18788 21879 18840 21888
rect 18788 21845 18797 21879
rect 18797 21845 18831 21879
rect 18831 21845 18840 21879
rect 18788 21836 18840 21845
rect 18972 21836 19024 21888
rect 19708 21972 19760 22024
rect 20904 21972 20956 22024
rect 23940 22083 23992 22092
rect 23940 22049 23949 22083
rect 23949 22049 23983 22083
rect 23983 22049 23992 22083
rect 23940 22040 23992 22049
rect 25412 22083 25464 22092
rect 22100 21972 22152 22024
rect 25412 22049 25420 22083
rect 25420 22049 25454 22083
rect 25454 22049 25464 22083
rect 25412 22040 25464 22049
rect 25872 22040 25924 22092
rect 26700 22108 26752 22160
rect 27804 22176 27856 22228
rect 27344 22151 27396 22160
rect 27344 22117 27353 22151
rect 27353 22117 27387 22151
rect 27387 22117 27396 22151
rect 27344 22108 27396 22117
rect 24492 22015 24544 22024
rect 24492 21981 24501 22015
rect 24501 21981 24535 22015
rect 24535 21981 24544 22015
rect 24492 21972 24544 21981
rect 24768 21972 24820 22024
rect 25228 21972 25280 22024
rect 27528 22040 27580 22092
rect 27988 22083 28040 22092
rect 27988 22049 27997 22083
rect 27997 22049 28031 22083
rect 28031 22049 28040 22083
rect 27988 22040 28040 22049
rect 28080 22040 28132 22092
rect 20076 21836 20128 21888
rect 20628 21879 20680 21888
rect 20628 21845 20637 21879
rect 20637 21845 20671 21879
rect 20671 21845 20680 21879
rect 20628 21836 20680 21845
rect 24676 21836 24728 21888
rect 25504 21904 25556 21956
rect 26332 21972 26384 22024
rect 27436 22015 27488 22024
rect 27436 21981 27445 22015
rect 27445 21981 27479 22015
rect 27479 21981 27488 22015
rect 27436 21972 27488 21981
rect 31668 22083 31720 22092
rect 31668 22049 31677 22083
rect 31677 22049 31711 22083
rect 31711 22049 31720 22083
rect 31668 22040 31720 22049
rect 25780 21879 25832 21888
rect 25780 21845 25789 21879
rect 25789 21845 25823 21879
rect 25823 21845 25832 21879
rect 25780 21836 25832 21845
rect 26056 21836 26108 21888
rect 26700 21836 26752 21888
rect 26792 21836 26844 21888
rect 26976 21836 27028 21888
rect 6286 21734 6338 21786
rect 6350 21734 6402 21786
rect 6414 21734 6466 21786
rect 6478 21734 6530 21786
rect 6542 21734 6594 21786
rect 13646 21734 13698 21786
rect 13710 21734 13762 21786
rect 13774 21734 13826 21786
rect 13838 21734 13890 21786
rect 13902 21734 13954 21786
rect 21006 21734 21058 21786
rect 21070 21734 21122 21786
rect 21134 21734 21186 21786
rect 21198 21734 21250 21786
rect 21262 21734 21314 21786
rect 28366 21734 28418 21786
rect 28430 21734 28482 21786
rect 28494 21734 28546 21786
rect 28558 21734 28610 21786
rect 28622 21734 28674 21786
rect 3240 21632 3292 21684
rect 6184 21632 6236 21684
rect 7472 21675 7524 21684
rect 7472 21641 7481 21675
rect 7481 21641 7515 21675
rect 7515 21641 7524 21675
rect 7472 21632 7524 21641
rect 7932 21675 7984 21684
rect 7932 21641 7941 21675
rect 7941 21641 7975 21675
rect 7975 21641 7984 21675
rect 7932 21632 7984 21641
rect 8116 21632 8168 21684
rect 11336 21632 11388 21684
rect 11796 21675 11848 21684
rect 11796 21641 11805 21675
rect 11805 21641 11839 21675
rect 11839 21641 11848 21675
rect 11796 21632 11848 21641
rect 12808 21632 12860 21684
rect 14004 21632 14056 21684
rect 6828 21564 6880 21616
rect 6000 21539 6052 21548
rect 6000 21505 6009 21539
rect 6009 21505 6043 21539
rect 6043 21505 6052 21539
rect 6000 21496 6052 21505
rect 6736 21496 6788 21548
rect 4620 21403 4672 21412
rect 4620 21369 4629 21403
rect 4629 21369 4663 21403
rect 4663 21369 4672 21403
rect 4620 21360 4672 21369
rect 4712 21292 4764 21344
rect 5724 21292 5776 21344
rect 7104 21471 7156 21480
rect 7104 21437 7113 21471
rect 7113 21437 7147 21471
rect 7147 21437 7156 21471
rect 7104 21428 7156 21437
rect 7288 21471 7340 21480
rect 7288 21437 7297 21471
rect 7297 21437 7331 21471
rect 7331 21437 7340 21471
rect 8484 21564 8536 21616
rect 8392 21496 8444 21548
rect 9588 21496 9640 21548
rect 9680 21496 9732 21548
rect 7288 21428 7340 21437
rect 7932 21428 7984 21480
rect 9956 21428 10008 21480
rect 8024 21292 8076 21344
rect 10232 21360 10284 21412
rect 9680 21292 9732 21344
rect 10416 21335 10468 21344
rect 10416 21301 10425 21335
rect 10425 21301 10459 21335
rect 10459 21301 10468 21335
rect 10416 21292 10468 21301
rect 12072 21292 12124 21344
rect 12900 21360 12952 21412
rect 13452 21360 13504 21412
rect 14188 21496 14240 21548
rect 14004 21360 14056 21412
rect 14832 21632 14884 21684
rect 15200 21675 15252 21684
rect 15200 21641 15209 21675
rect 15209 21641 15243 21675
rect 15243 21641 15252 21675
rect 15200 21632 15252 21641
rect 16120 21632 16172 21684
rect 18236 21675 18288 21684
rect 18236 21641 18245 21675
rect 18245 21641 18279 21675
rect 18279 21641 18288 21675
rect 18236 21632 18288 21641
rect 18420 21632 18472 21684
rect 20720 21632 20772 21684
rect 20904 21675 20956 21684
rect 20904 21641 20913 21675
rect 20913 21641 20947 21675
rect 20947 21641 20956 21675
rect 20904 21632 20956 21641
rect 15568 21564 15620 21616
rect 16212 21564 16264 21616
rect 17132 21564 17184 21616
rect 23756 21564 23808 21616
rect 24124 21564 24176 21616
rect 15108 21428 15160 21480
rect 15292 21471 15344 21480
rect 15292 21437 15301 21471
rect 15301 21437 15335 21471
rect 15335 21437 15344 21471
rect 15292 21428 15344 21437
rect 18788 21496 18840 21548
rect 15476 21428 15528 21480
rect 15844 21428 15896 21480
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 15016 21292 15068 21344
rect 16028 21403 16080 21412
rect 16028 21369 16037 21403
rect 16037 21369 16071 21403
rect 16071 21369 16080 21403
rect 16028 21360 16080 21369
rect 16396 21360 16448 21412
rect 16672 21360 16724 21412
rect 17500 21428 17552 21480
rect 18052 21428 18104 21480
rect 17132 21403 17184 21412
rect 17132 21369 17141 21403
rect 17141 21369 17175 21403
rect 17175 21369 17184 21403
rect 17132 21360 17184 21369
rect 15660 21292 15712 21344
rect 15844 21292 15896 21344
rect 16580 21335 16632 21344
rect 16580 21301 16589 21335
rect 16589 21301 16623 21335
rect 16623 21301 16632 21335
rect 16580 21292 16632 21301
rect 17224 21292 17276 21344
rect 20628 21496 20680 21548
rect 20076 21428 20128 21480
rect 20536 21471 20588 21480
rect 20536 21437 20545 21471
rect 20545 21437 20579 21471
rect 20579 21437 20588 21471
rect 20536 21428 20588 21437
rect 19800 21360 19852 21412
rect 21456 21292 21508 21344
rect 22100 21292 22152 21344
rect 23296 21471 23348 21480
rect 23296 21437 23305 21471
rect 23305 21437 23339 21471
rect 23339 21437 23348 21471
rect 23296 21428 23348 21437
rect 24492 21632 24544 21684
rect 26056 21632 26108 21684
rect 24676 21564 24728 21616
rect 25228 21564 25280 21616
rect 27988 21632 28040 21684
rect 26148 21496 26200 21548
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 26792 21496 26844 21548
rect 27068 21496 27120 21548
rect 24952 21428 25004 21480
rect 25044 21428 25096 21480
rect 30196 21496 30248 21548
rect 22836 21360 22888 21412
rect 23388 21360 23440 21412
rect 25688 21403 25740 21412
rect 25688 21369 25697 21403
rect 25697 21369 25731 21403
rect 25731 21369 25740 21403
rect 25688 21360 25740 21369
rect 25872 21403 25924 21412
rect 25872 21369 25881 21403
rect 25881 21369 25915 21403
rect 25915 21369 25924 21403
rect 25872 21360 25924 21369
rect 26976 21360 27028 21412
rect 24032 21292 24084 21344
rect 24216 21292 24268 21344
rect 24952 21292 25004 21344
rect 25412 21292 25464 21344
rect 26516 21292 26568 21344
rect 26792 21292 26844 21344
rect 27712 21292 27764 21344
rect 28172 21335 28224 21344
rect 28172 21301 28181 21335
rect 28181 21301 28215 21335
rect 28215 21301 28224 21335
rect 28172 21292 28224 21301
rect 28724 21292 28776 21344
rect 6946 21190 6998 21242
rect 7010 21190 7062 21242
rect 7074 21190 7126 21242
rect 7138 21190 7190 21242
rect 7202 21190 7254 21242
rect 14306 21190 14358 21242
rect 14370 21190 14422 21242
rect 14434 21190 14486 21242
rect 14498 21190 14550 21242
rect 14562 21190 14614 21242
rect 21666 21190 21718 21242
rect 21730 21190 21782 21242
rect 21794 21190 21846 21242
rect 21858 21190 21910 21242
rect 21922 21190 21974 21242
rect 29026 21190 29078 21242
rect 29090 21190 29142 21242
rect 29154 21190 29206 21242
rect 29218 21190 29270 21242
rect 29282 21190 29334 21242
rect 4160 21088 4212 21140
rect 4620 21088 4672 21140
rect 11060 21088 11112 21140
rect 10048 21063 10100 21072
rect 10048 21029 10057 21063
rect 10057 21029 10091 21063
rect 10091 21029 10100 21063
rect 10048 21020 10100 21029
rect 10784 21020 10836 21072
rect 11612 21088 11664 21140
rect 14096 21088 14148 21140
rect 15108 21088 15160 21140
rect 11980 21020 12032 21072
rect 12440 21020 12492 21072
rect 13360 21020 13412 21072
rect 13544 21020 13596 21072
rect 3332 20995 3384 21004
rect 3332 20961 3341 20995
rect 3341 20961 3375 20995
rect 3375 20961 3384 20995
rect 3332 20952 3384 20961
rect 5908 20952 5960 21004
rect 9588 20952 9640 21004
rect 3056 20927 3108 20936
rect 3056 20893 3065 20927
rect 3065 20893 3099 20927
rect 3099 20893 3108 20927
rect 3056 20884 3108 20893
rect 4252 20927 4304 20936
rect 4252 20893 4261 20927
rect 4261 20893 4295 20927
rect 4295 20893 4304 20927
rect 4252 20884 4304 20893
rect 5816 20927 5868 20936
rect 5816 20893 5825 20927
rect 5825 20893 5859 20927
rect 5859 20893 5868 20927
rect 5816 20884 5868 20893
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 8208 20884 8260 20936
rect 13268 20952 13320 21004
rect 14004 20995 14056 21004
rect 14004 20961 14038 20995
rect 14038 20961 14056 20995
rect 14004 20952 14056 20961
rect 14188 20952 14240 21004
rect 14464 20952 14516 21004
rect 15016 20952 15068 21004
rect 12256 20927 12308 20936
rect 12256 20893 12265 20927
rect 12265 20893 12299 20927
rect 12299 20893 12308 20927
rect 12256 20884 12308 20893
rect 12992 20884 13044 20936
rect 12624 20816 12676 20868
rect 5264 20791 5316 20800
rect 5264 20757 5273 20791
rect 5273 20757 5307 20791
rect 5307 20757 5316 20791
rect 5264 20748 5316 20757
rect 12808 20748 12860 20800
rect 13820 20927 13872 20936
rect 13820 20893 13829 20927
rect 13829 20893 13863 20927
rect 13863 20893 13872 20927
rect 13820 20884 13872 20893
rect 15936 21020 15988 21072
rect 16856 21020 16908 21072
rect 19064 21020 19116 21072
rect 20628 21088 20680 21140
rect 23296 21088 23348 21140
rect 20904 21020 20956 21072
rect 21548 21063 21600 21072
rect 21548 21029 21557 21063
rect 21557 21029 21591 21063
rect 21591 21029 21600 21063
rect 21548 21020 21600 21029
rect 24676 21088 24728 21140
rect 27804 21088 27856 21140
rect 28172 21088 28224 21140
rect 15660 20952 15712 21004
rect 20812 20952 20864 21004
rect 23572 20952 23624 21004
rect 24032 20952 24084 21004
rect 24216 20952 24268 21004
rect 24400 20995 24452 21004
rect 24400 20961 24409 20995
rect 24409 20961 24443 20995
rect 24443 20961 24452 20995
rect 24400 20952 24452 20961
rect 18328 20927 18380 20936
rect 18328 20893 18337 20927
rect 18337 20893 18371 20927
rect 18371 20893 18380 20927
rect 18328 20884 18380 20893
rect 14556 20748 14608 20800
rect 14924 20748 14976 20800
rect 16672 20748 16724 20800
rect 17040 20748 17092 20800
rect 20720 20884 20772 20936
rect 22100 20816 22152 20868
rect 23020 20816 23072 20868
rect 18696 20748 18748 20800
rect 23940 20791 23992 20800
rect 23940 20757 23949 20791
rect 23949 20757 23983 20791
rect 23983 20757 23992 20791
rect 23940 20748 23992 20757
rect 24124 20816 24176 20868
rect 25504 21020 25556 21072
rect 27712 21020 27764 21072
rect 24584 20995 24636 21004
rect 24584 20961 24593 20995
rect 24593 20961 24627 20995
rect 24627 20961 24636 20995
rect 24584 20952 24636 20961
rect 24768 20995 24820 21004
rect 24768 20961 24777 20995
rect 24777 20961 24811 20995
rect 24811 20961 24820 20995
rect 24768 20952 24820 20961
rect 24860 20952 24912 21004
rect 25320 20884 25372 20936
rect 25688 20952 25740 21004
rect 25504 20927 25556 20936
rect 25504 20893 25513 20927
rect 25513 20893 25547 20927
rect 25547 20893 25556 20927
rect 25504 20884 25556 20893
rect 24952 20748 25004 20800
rect 25688 20791 25740 20800
rect 25688 20757 25697 20791
rect 25697 20757 25731 20791
rect 25731 20757 25740 20791
rect 25688 20748 25740 20757
rect 26056 20927 26108 20936
rect 26056 20893 26065 20927
rect 26065 20893 26099 20927
rect 26099 20893 26108 20927
rect 26056 20884 26108 20893
rect 26148 20884 26200 20936
rect 29552 20884 29604 20936
rect 29644 20884 29696 20936
rect 33048 20884 33100 20936
rect 26424 20748 26476 20800
rect 27620 20791 27672 20800
rect 27620 20757 27629 20791
rect 27629 20757 27663 20791
rect 27663 20757 27672 20791
rect 27620 20748 27672 20757
rect 27712 20748 27764 20800
rect 30012 20791 30064 20800
rect 30012 20757 30021 20791
rect 30021 20757 30055 20791
rect 30055 20757 30064 20791
rect 30012 20748 30064 20757
rect 30104 20791 30156 20800
rect 30104 20757 30113 20791
rect 30113 20757 30147 20791
rect 30147 20757 30156 20791
rect 30104 20748 30156 20757
rect 6286 20646 6338 20698
rect 6350 20646 6402 20698
rect 6414 20646 6466 20698
rect 6478 20646 6530 20698
rect 6542 20646 6594 20698
rect 13646 20646 13698 20698
rect 13710 20646 13762 20698
rect 13774 20646 13826 20698
rect 13838 20646 13890 20698
rect 13902 20646 13954 20698
rect 21006 20646 21058 20698
rect 21070 20646 21122 20698
rect 21134 20646 21186 20698
rect 21198 20646 21250 20698
rect 21262 20646 21314 20698
rect 28366 20646 28418 20698
rect 28430 20646 28482 20698
rect 28494 20646 28546 20698
rect 28558 20646 28610 20698
rect 28622 20646 28674 20698
rect 4252 20544 4304 20596
rect 5816 20544 5868 20596
rect 9680 20544 9732 20596
rect 8024 20476 8076 20528
rect 10508 20544 10560 20596
rect 11152 20544 11204 20596
rect 11612 20587 11664 20596
rect 5816 20408 5868 20460
rect 6092 20451 6144 20460
rect 6092 20417 6101 20451
rect 6101 20417 6135 20451
rect 6135 20417 6144 20451
rect 6092 20408 6144 20417
rect 8392 20408 8444 20460
rect 9588 20408 9640 20460
rect 10876 20408 10928 20460
rect 5908 20340 5960 20392
rect 6000 20204 6052 20256
rect 10048 20340 10100 20392
rect 11612 20553 11621 20587
rect 11621 20553 11655 20587
rect 11655 20553 11664 20587
rect 11612 20544 11664 20553
rect 14188 20587 14240 20596
rect 14188 20553 14197 20587
rect 14197 20553 14231 20587
rect 14231 20553 14240 20587
rect 14188 20544 14240 20553
rect 14556 20544 14608 20596
rect 15292 20544 15344 20596
rect 15384 20544 15436 20596
rect 18696 20544 18748 20596
rect 19064 20544 19116 20596
rect 20720 20544 20772 20596
rect 23940 20544 23992 20596
rect 24124 20544 24176 20596
rect 11980 20451 12032 20460
rect 11980 20417 11989 20451
rect 11989 20417 12023 20451
rect 12023 20417 12032 20451
rect 11980 20408 12032 20417
rect 6368 20315 6420 20324
rect 6368 20281 6377 20315
rect 6377 20281 6411 20315
rect 6411 20281 6420 20315
rect 6368 20272 6420 20281
rect 7380 20272 7432 20324
rect 8944 20315 8996 20324
rect 8944 20281 8953 20315
rect 8953 20281 8987 20315
rect 8987 20281 8996 20315
rect 8944 20272 8996 20281
rect 11060 20315 11112 20324
rect 11060 20281 11069 20315
rect 11069 20281 11103 20315
rect 11103 20281 11112 20315
rect 11060 20272 11112 20281
rect 7288 20204 7340 20256
rect 8116 20204 8168 20256
rect 9312 20204 9364 20256
rect 16580 20476 16632 20528
rect 12256 20408 12308 20460
rect 12440 20451 12492 20460
rect 12440 20417 12474 20451
rect 12474 20417 12492 20451
rect 12440 20408 12492 20417
rect 12624 20340 12676 20392
rect 14648 20408 14700 20460
rect 15200 20408 15252 20460
rect 18696 20408 18748 20460
rect 14740 20340 14792 20392
rect 15384 20340 15436 20392
rect 15936 20340 15988 20392
rect 19064 20383 19116 20392
rect 19064 20349 19073 20383
rect 19073 20349 19107 20383
rect 19107 20349 19116 20383
rect 19800 20408 19852 20460
rect 21364 20408 21416 20460
rect 22100 20408 22152 20460
rect 24032 20451 24084 20460
rect 24032 20417 24041 20451
rect 24041 20417 24075 20451
rect 24075 20417 24084 20451
rect 24032 20408 24084 20417
rect 24676 20451 24728 20460
rect 24676 20417 24685 20451
rect 24685 20417 24719 20451
rect 24719 20417 24728 20451
rect 24676 20408 24728 20417
rect 19064 20340 19116 20349
rect 22928 20340 22980 20392
rect 19984 20272 20036 20324
rect 22008 20272 22060 20324
rect 12716 20204 12768 20256
rect 13084 20204 13136 20256
rect 13544 20204 13596 20256
rect 14096 20204 14148 20256
rect 14648 20247 14700 20256
rect 14648 20213 14657 20247
rect 14657 20213 14691 20247
rect 14691 20213 14700 20247
rect 14648 20204 14700 20213
rect 14740 20204 14792 20256
rect 15660 20204 15712 20256
rect 20444 20204 20496 20256
rect 21088 20247 21140 20256
rect 21088 20213 21097 20247
rect 21097 20213 21131 20247
rect 21131 20213 21140 20247
rect 21088 20204 21140 20213
rect 23388 20383 23440 20392
rect 23388 20349 23397 20383
rect 23397 20349 23431 20383
rect 23431 20349 23440 20383
rect 23388 20340 23440 20349
rect 23756 20340 23808 20392
rect 23848 20383 23900 20392
rect 23848 20349 23857 20383
rect 23857 20349 23891 20383
rect 23891 20349 23900 20383
rect 23848 20340 23900 20349
rect 24124 20383 24176 20392
rect 24124 20349 24133 20383
rect 24133 20349 24167 20383
rect 24167 20349 24176 20383
rect 24124 20340 24176 20349
rect 23940 20204 23992 20256
rect 24308 20247 24360 20256
rect 24308 20213 24317 20247
rect 24317 20213 24351 20247
rect 24351 20213 24360 20247
rect 24308 20204 24360 20213
rect 24676 20204 24728 20256
rect 25044 20544 25096 20596
rect 25504 20544 25556 20596
rect 25596 20587 25648 20596
rect 25596 20553 25605 20587
rect 25605 20553 25639 20587
rect 25639 20553 25648 20587
rect 25596 20544 25648 20553
rect 25688 20544 25740 20596
rect 26792 20544 26844 20596
rect 27988 20544 28040 20596
rect 29644 20544 29696 20596
rect 29828 20544 29880 20596
rect 26148 20519 26200 20528
rect 26148 20485 26157 20519
rect 26157 20485 26191 20519
rect 26191 20485 26200 20519
rect 26148 20476 26200 20485
rect 25136 20408 25188 20460
rect 25504 20451 25556 20460
rect 25504 20417 25513 20451
rect 25513 20417 25547 20451
rect 25547 20417 25556 20451
rect 25504 20408 25556 20417
rect 26424 20451 26476 20460
rect 26424 20417 26433 20451
rect 26433 20417 26467 20451
rect 26467 20417 26476 20451
rect 26424 20408 26476 20417
rect 29368 20408 29420 20460
rect 24860 20340 24912 20392
rect 25688 20383 25740 20392
rect 25688 20349 25697 20383
rect 25697 20349 25731 20383
rect 25731 20349 25740 20383
rect 25688 20340 25740 20349
rect 25780 20340 25832 20392
rect 26332 20340 26384 20392
rect 28172 20340 28224 20392
rect 26700 20204 26752 20256
rect 28080 20272 28132 20324
rect 29460 20272 29512 20324
rect 30012 20315 30064 20324
rect 30012 20281 30021 20315
rect 30021 20281 30055 20315
rect 30055 20281 30064 20315
rect 30012 20272 30064 20281
rect 28172 20204 28224 20256
rect 30104 20204 30156 20256
rect 30656 20204 30708 20256
rect 31208 20204 31260 20256
rect 6946 20102 6998 20154
rect 7010 20102 7062 20154
rect 7074 20102 7126 20154
rect 7138 20102 7190 20154
rect 7202 20102 7254 20154
rect 14306 20102 14358 20154
rect 14370 20102 14422 20154
rect 14434 20102 14486 20154
rect 14498 20102 14550 20154
rect 14562 20102 14614 20154
rect 21666 20102 21718 20154
rect 21730 20102 21782 20154
rect 21794 20102 21846 20154
rect 21858 20102 21910 20154
rect 21922 20102 21974 20154
rect 29026 20102 29078 20154
rect 29090 20102 29142 20154
rect 29154 20102 29206 20154
rect 29218 20102 29270 20154
rect 29282 20102 29334 20154
rect 6368 20000 6420 20052
rect 6736 20000 6788 20052
rect 7380 20000 7432 20052
rect 5264 19932 5316 19984
rect 5724 19932 5776 19984
rect 8944 20000 8996 20052
rect 10048 20000 10100 20052
rect 11612 20000 11664 20052
rect 14740 20000 14792 20052
rect 15108 20000 15160 20052
rect 16488 20000 16540 20052
rect 19064 20000 19116 20052
rect 19248 20043 19300 20052
rect 19248 20009 19257 20043
rect 19257 20009 19291 20043
rect 19291 20009 19300 20043
rect 19248 20000 19300 20009
rect 20444 20043 20496 20052
rect 20444 20009 20453 20043
rect 20453 20009 20487 20043
rect 20487 20009 20496 20043
rect 20444 20000 20496 20009
rect 21088 20000 21140 20052
rect 22008 20000 22060 20052
rect 23664 20043 23716 20052
rect 8116 19932 8168 19984
rect 9864 19932 9916 19984
rect 14280 19932 14332 19984
rect 15476 19932 15528 19984
rect 15660 19932 15712 19984
rect 16764 19932 16816 19984
rect 6920 19864 6972 19916
rect 7288 19864 7340 19916
rect 7380 19864 7432 19916
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 5724 19796 5776 19848
rect 8024 19796 8076 19848
rect 9312 19864 9364 19916
rect 9588 19907 9640 19916
rect 9588 19873 9597 19907
rect 9597 19873 9631 19907
rect 9631 19873 9640 19907
rect 9588 19864 9640 19873
rect 9680 19907 9732 19916
rect 9680 19873 9689 19907
rect 9689 19873 9723 19907
rect 9723 19873 9732 19907
rect 9680 19864 9732 19873
rect 9772 19907 9824 19916
rect 9772 19873 9781 19907
rect 9781 19873 9815 19907
rect 9815 19873 9824 19907
rect 9772 19864 9824 19873
rect 10232 19907 10284 19916
rect 10232 19873 10241 19907
rect 10241 19873 10275 19907
rect 10275 19873 10284 19907
rect 10232 19864 10284 19873
rect 10416 19864 10468 19916
rect 11060 19864 11112 19916
rect 12256 19864 12308 19916
rect 12808 19864 12860 19916
rect 12900 19864 12952 19916
rect 6000 19728 6052 19780
rect 9772 19728 9824 19780
rect 11336 19728 11388 19780
rect 11612 19728 11664 19780
rect 12624 19728 12676 19780
rect 13268 19839 13320 19848
rect 13268 19805 13277 19839
rect 13277 19805 13311 19839
rect 13311 19805 13320 19839
rect 13268 19796 13320 19805
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 14740 19907 14792 19916
rect 14740 19873 14749 19907
rect 14749 19873 14783 19907
rect 14783 19873 14792 19907
rect 14740 19864 14792 19873
rect 14924 19796 14976 19848
rect 15568 19907 15620 19916
rect 15568 19873 15579 19907
rect 15579 19873 15613 19907
rect 15613 19873 15620 19907
rect 15568 19864 15620 19873
rect 18420 19864 18472 19916
rect 15200 19796 15252 19848
rect 18144 19796 18196 19848
rect 9220 19703 9272 19712
rect 9220 19669 9229 19703
rect 9229 19669 9263 19703
rect 9263 19669 9272 19703
rect 9220 19660 9272 19669
rect 10232 19660 10284 19712
rect 14004 19703 14056 19712
rect 14004 19669 14013 19703
rect 14013 19669 14047 19703
rect 14047 19669 14056 19703
rect 14004 19660 14056 19669
rect 14740 19728 14792 19780
rect 16672 19728 16724 19780
rect 16764 19728 16816 19780
rect 20168 19728 20220 19780
rect 21732 19839 21784 19848
rect 21732 19805 21741 19839
rect 21741 19805 21775 19839
rect 21775 19805 21784 19839
rect 21732 19796 21784 19805
rect 15292 19660 15344 19712
rect 15476 19660 15528 19712
rect 16212 19660 16264 19712
rect 17684 19660 17736 19712
rect 18420 19703 18472 19712
rect 18420 19669 18429 19703
rect 18429 19669 18463 19703
rect 18463 19669 18472 19703
rect 18420 19660 18472 19669
rect 20260 19660 20312 19712
rect 21548 19660 21600 19712
rect 23664 20009 23673 20043
rect 23673 20009 23707 20043
rect 23707 20009 23716 20043
rect 23664 20000 23716 20009
rect 23848 20000 23900 20052
rect 24584 20000 24636 20052
rect 26332 20043 26384 20052
rect 26332 20009 26341 20043
rect 26341 20009 26375 20043
rect 26375 20009 26384 20043
rect 26332 20000 26384 20009
rect 27436 20000 27488 20052
rect 27528 20000 27580 20052
rect 23940 19932 23992 19984
rect 22836 19864 22888 19916
rect 23020 19907 23072 19916
rect 23020 19873 23029 19907
rect 23029 19873 23063 19907
rect 23063 19873 23072 19907
rect 23020 19864 23072 19873
rect 23204 19907 23256 19916
rect 23204 19873 23213 19907
rect 23213 19873 23247 19907
rect 23247 19873 23256 19907
rect 23204 19864 23256 19873
rect 23572 19864 23624 19916
rect 25688 19864 25740 19916
rect 23848 19796 23900 19848
rect 24768 19796 24820 19848
rect 22928 19728 22980 19780
rect 24216 19728 24268 19780
rect 22744 19660 22796 19712
rect 23204 19660 23256 19712
rect 25688 19728 25740 19780
rect 26332 19864 26384 19916
rect 27712 19932 27764 19984
rect 26700 19796 26752 19848
rect 27620 19864 27672 19916
rect 28172 20000 28224 20052
rect 29552 20000 29604 20052
rect 29828 20000 29880 20052
rect 28264 19932 28316 19984
rect 28908 19975 28960 19984
rect 28908 19941 28917 19975
rect 28917 19941 28951 19975
rect 28951 19941 28960 19975
rect 28908 19932 28960 19941
rect 27988 19864 28040 19916
rect 24768 19660 24820 19712
rect 25136 19703 25188 19712
rect 25136 19669 25145 19703
rect 25145 19669 25179 19703
rect 25179 19669 25188 19703
rect 25136 19660 25188 19669
rect 25964 19703 26016 19712
rect 25964 19669 25973 19703
rect 25973 19669 26007 19703
rect 26007 19669 26016 19703
rect 25964 19660 26016 19669
rect 26608 19660 26660 19712
rect 27252 19703 27304 19712
rect 27252 19669 27261 19703
rect 27261 19669 27295 19703
rect 27295 19669 27304 19703
rect 27252 19660 27304 19669
rect 27804 19660 27856 19712
rect 29000 19796 29052 19848
rect 29920 19932 29972 19984
rect 28724 19728 28776 19780
rect 30656 19907 30708 19916
rect 30656 19873 30665 19907
rect 30665 19873 30699 19907
rect 30699 19873 30708 19907
rect 30656 19864 30708 19873
rect 30840 19907 30892 19916
rect 30840 19873 30858 19907
rect 30858 19873 30892 19907
rect 30840 19864 30892 19873
rect 31484 19796 31536 19848
rect 31208 19771 31260 19780
rect 31208 19737 31217 19771
rect 31217 19737 31251 19771
rect 31251 19737 31260 19771
rect 31208 19728 31260 19737
rect 31392 19728 31444 19780
rect 28264 19703 28316 19712
rect 28264 19669 28273 19703
rect 28273 19669 28307 19703
rect 28307 19669 28316 19703
rect 28264 19660 28316 19669
rect 29460 19660 29512 19712
rect 30012 19703 30064 19712
rect 30012 19669 30021 19703
rect 30021 19669 30055 19703
rect 30055 19669 30064 19703
rect 30012 19660 30064 19669
rect 30656 19660 30708 19712
rect 6286 19558 6338 19610
rect 6350 19558 6402 19610
rect 6414 19558 6466 19610
rect 6478 19558 6530 19610
rect 6542 19558 6594 19610
rect 13646 19558 13698 19610
rect 13710 19558 13762 19610
rect 13774 19558 13826 19610
rect 13838 19558 13890 19610
rect 13902 19558 13954 19610
rect 21006 19558 21058 19610
rect 21070 19558 21122 19610
rect 21134 19558 21186 19610
rect 21198 19558 21250 19610
rect 21262 19558 21314 19610
rect 28366 19558 28418 19610
rect 28430 19558 28482 19610
rect 28494 19558 28546 19610
rect 28558 19558 28610 19610
rect 28622 19558 28674 19610
rect 14188 19456 14240 19508
rect 1308 19252 1360 19304
rect 7840 19295 7892 19304
rect 7840 19261 7849 19295
rect 7849 19261 7883 19295
rect 7883 19261 7892 19295
rect 7840 19252 7892 19261
rect 9588 19320 9640 19372
rect 10048 19320 10100 19372
rect 9220 19252 9272 19304
rect 3240 19159 3292 19168
rect 3240 19125 3249 19159
rect 3249 19125 3283 19159
rect 3283 19125 3292 19159
rect 3240 19116 3292 19125
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 8852 19116 8904 19168
rect 8944 19116 8996 19168
rect 10508 19252 10560 19304
rect 10692 19295 10744 19304
rect 10692 19261 10701 19295
rect 10701 19261 10735 19295
rect 10735 19261 10744 19295
rect 10692 19252 10744 19261
rect 11796 19295 11848 19304
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 12164 19252 12216 19304
rect 11888 19184 11940 19236
rect 9404 19116 9456 19168
rect 9772 19116 9824 19168
rect 9956 19116 10008 19168
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 11428 19116 11480 19168
rect 11980 19159 12032 19168
rect 11980 19125 11989 19159
rect 11989 19125 12023 19159
rect 12023 19125 12032 19159
rect 11980 19116 12032 19125
rect 14464 19320 14516 19372
rect 12532 19295 12584 19304
rect 12532 19261 12541 19295
rect 12541 19261 12575 19295
rect 12575 19261 12584 19295
rect 12532 19252 12584 19261
rect 14740 19252 14792 19304
rect 12808 19227 12860 19236
rect 12808 19193 12817 19227
rect 12817 19193 12851 19227
rect 12851 19193 12860 19227
rect 12808 19184 12860 19193
rect 14096 19184 14148 19236
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 16856 19252 16908 19304
rect 15200 19184 15252 19236
rect 15752 19184 15804 19236
rect 14728 19116 14780 19168
rect 15016 19116 15068 19168
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15292 19116 15344 19125
rect 16028 19116 16080 19168
rect 16120 19159 16172 19168
rect 16120 19125 16129 19159
rect 16129 19125 16163 19159
rect 16163 19125 16172 19159
rect 16120 19116 16172 19125
rect 16948 19159 17000 19168
rect 16948 19125 16957 19159
rect 16957 19125 16991 19159
rect 16991 19125 17000 19159
rect 16948 19116 17000 19125
rect 18420 19252 18472 19304
rect 19800 19456 19852 19508
rect 17408 19227 17460 19236
rect 17408 19193 17417 19227
rect 17417 19193 17451 19227
rect 17451 19193 17460 19227
rect 17408 19184 17460 19193
rect 19156 19227 19208 19236
rect 19156 19193 19165 19227
rect 19165 19193 19199 19227
rect 19199 19193 19208 19227
rect 19156 19184 19208 19193
rect 21732 19456 21784 19508
rect 22744 19456 22796 19508
rect 23664 19456 23716 19508
rect 24032 19456 24084 19508
rect 24584 19456 24636 19508
rect 24676 19456 24728 19508
rect 24768 19456 24820 19508
rect 26332 19456 26384 19508
rect 20628 19320 20680 19372
rect 23480 19320 23532 19372
rect 25504 19388 25556 19440
rect 26608 19456 26660 19508
rect 28080 19456 28132 19508
rect 28908 19499 28960 19508
rect 28908 19465 28917 19499
rect 28917 19465 28951 19499
rect 28951 19465 28960 19499
rect 28908 19456 28960 19465
rect 18052 19116 18104 19168
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 20352 19116 20404 19168
rect 20904 19184 20956 19236
rect 23756 19252 23808 19304
rect 25964 19320 26016 19372
rect 22652 19184 22704 19236
rect 21272 19116 21324 19168
rect 21548 19116 21600 19168
rect 24400 19159 24452 19168
rect 24400 19125 24409 19159
rect 24409 19125 24443 19159
rect 24443 19125 24452 19159
rect 24400 19116 24452 19125
rect 24584 19116 24636 19168
rect 25412 19252 25464 19304
rect 27252 19320 27304 19372
rect 27436 19295 27488 19304
rect 27436 19261 27445 19295
rect 27445 19261 27479 19295
rect 27479 19261 27488 19295
rect 27436 19252 27488 19261
rect 27804 19363 27856 19372
rect 27804 19329 27813 19363
rect 27813 19329 27847 19363
rect 27847 19329 27856 19363
rect 27804 19320 27856 19329
rect 27896 19363 27948 19372
rect 27896 19329 27905 19363
rect 27905 19329 27939 19363
rect 27939 19329 27948 19363
rect 27896 19320 27948 19329
rect 28264 19320 28316 19372
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 25872 19116 25924 19168
rect 27712 19184 27764 19236
rect 27344 19116 27396 19168
rect 27988 19116 28040 19168
rect 28356 19116 28408 19168
rect 28724 19252 28776 19304
rect 29552 19227 29604 19236
rect 29552 19193 29561 19227
rect 29561 19193 29595 19227
rect 29595 19193 29604 19227
rect 29552 19184 29604 19193
rect 30288 19184 30340 19236
rect 29368 19116 29420 19168
rect 31024 19159 31076 19168
rect 31024 19125 31033 19159
rect 31033 19125 31067 19159
rect 31067 19125 31076 19159
rect 31024 19116 31076 19125
rect 31208 19159 31260 19168
rect 31208 19125 31217 19159
rect 31217 19125 31251 19159
rect 31251 19125 31260 19159
rect 31208 19116 31260 19125
rect 6946 19014 6998 19066
rect 7010 19014 7062 19066
rect 7074 19014 7126 19066
rect 7138 19014 7190 19066
rect 7202 19014 7254 19066
rect 14306 19014 14358 19066
rect 14370 19014 14422 19066
rect 14434 19014 14486 19066
rect 14498 19014 14550 19066
rect 14562 19014 14614 19066
rect 21666 19014 21718 19066
rect 21730 19014 21782 19066
rect 21794 19014 21846 19066
rect 21858 19014 21910 19066
rect 21922 19014 21974 19066
rect 29026 19014 29078 19066
rect 29090 19014 29142 19066
rect 29154 19014 29206 19066
rect 29218 19014 29270 19066
rect 29282 19014 29334 19066
rect 8944 18844 8996 18896
rect 9864 18844 9916 18896
rect 12808 18912 12860 18964
rect 13820 18912 13872 18964
rect 14096 18912 14148 18964
rect 14556 18912 14608 18964
rect 14740 18912 14792 18964
rect 15292 18912 15344 18964
rect 17408 18912 17460 18964
rect 17592 18912 17644 18964
rect 6092 18776 6144 18828
rect 9680 18776 9732 18828
rect 10968 18776 11020 18828
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 4988 18751 5040 18760
rect 4988 18717 4997 18751
rect 4997 18717 5031 18751
rect 5031 18717 5040 18751
rect 4988 18708 5040 18717
rect 6184 18640 6236 18692
rect 5172 18572 5224 18624
rect 6000 18572 6052 18624
rect 7932 18708 7984 18760
rect 8852 18640 8904 18692
rect 9772 18708 9824 18760
rect 9864 18751 9916 18760
rect 9864 18717 9873 18751
rect 9873 18717 9907 18751
rect 9907 18717 9916 18751
rect 9864 18708 9916 18717
rect 10048 18708 10100 18760
rect 12532 18844 12584 18896
rect 13452 18844 13504 18896
rect 15752 18844 15804 18896
rect 16948 18844 17000 18896
rect 19248 18844 19300 18896
rect 21088 18844 21140 18896
rect 12072 18819 12124 18828
rect 12072 18785 12081 18819
rect 12081 18785 12115 18819
rect 12115 18785 12124 18819
rect 12072 18776 12124 18785
rect 12900 18776 12952 18828
rect 13360 18776 13412 18828
rect 14188 18776 14240 18828
rect 15016 18819 15068 18828
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 12624 18708 12676 18717
rect 12992 18751 13044 18760
rect 12992 18717 13001 18751
rect 13001 18717 13035 18751
rect 13035 18717 13044 18751
rect 12992 18708 13044 18717
rect 13452 18708 13504 18760
rect 15016 18785 15025 18819
rect 15025 18785 15059 18819
rect 15059 18785 15068 18819
rect 15016 18776 15068 18785
rect 15200 18819 15252 18828
rect 15200 18785 15209 18819
rect 15209 18785 15243 18819
rect 15243 18785 15252 18819
rect 15200 18776 15252 18785
rect 8116 18615 8168 18624
rect 8116 18581 8125 18615
rect 8125 18581 8159 18615
rect 8159 18581 8168 18615
rect 8116 18572 8168 18581
rect 10140 18640 10192 18692
rect 14280 18640 14332 18692
rect 10508 18615 10560 18624
rect 10508 18581 10517 18615
rect 10517 18581 10551 18615
rect 10551 18581 10560 18615
rect 10508 18572 10560 18581
rect 12440 18572 12492 18624
rect 13084 18572 13136 18624
rect 14096 18615 14148 18624
rect 14096 18581 14105 18615
rect 14105 18581 14139 18615
rect 14139 18581 14148 18615
rect 14096 18572 14148 18581
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 16948 18708 17000 18760
rect 17776 18751 17828 18760
rect 17776 18717 17785 18751
rect 17785 18717 17819 18751
rect 17819 18717 17828 18751
rect 17776 18708 17828 18717
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 19156 18708 19208 18760
rect 19340 18751 19392 18760
rect 19340 18717 19349 18751
rect 19349 18717 19383 18751
rect 19383 18717 19392 18751
rect 19340 18708 19392 18717
rect 16488 18640 16540 18692
rect 16120 18572 16172 18624
rect 16764 18572 16816 18624
rect 18512 18640 18564 18692
rect 20352 18708 20404 18760
rect 22652 18955 22704 18964
rect 22652 18921 22661 18955
rect 22661 18921 22695 18955
rect 22695 18921 22704 18955
rect 22652 18912 22704 18921
rect 23388 18912 23440 18964
rect 23848 18912 23900 18964
rect 24124 18912 24176 18964
rect 22744 18819 22796 18828
rect 21456 18708 21508 18760
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 23756 18844 23808 18896
rect 26424 18912 26476 18964
rect 26516 18912 26568 18964
rect 27804 18912 27856 18964
rect 29552 18912 29604 18964
rect 30288 18955 30340 18964
rect 30288 18921 30297 18955
rect 30297 18921 30331 18955
rect 30331 18921 30340 18955
rect 30288 18912 30340 18921
rect 31208 18912 31260 18964
rect 24032 18776 24084 18828
rect 24676 18776 24728 18828
rect 24768 18819 24820 18828
rect 24768 18785 24777 18819
rect 24777 18785 24811 18819
rect 24811 18785 24820 18819
rect 24768 18776 24820 18785
rect 25136 18887 25188 18896
rect 25136 18853 25145 18887
rect 25145 18853 25179 18887
rect 25179 18853 25188 18887
rect 25136 18844 25188 18853
rect 25596 18844 25648 18896
rect 26792 18844 26844 18896
rect 33140 18844 33192 18896
rect 28356 18819 28408 18828
rect 25872 18708 25924 18760
rect 28356 18785 28365 18819
rect 28365 18785 28399 18819
rect 28399 18785 28408 18819
rect 28356 18776 28408 18785
rect 28908 18776 28960 18828
rect 30196 18819 30248 18828
rect 30196 18785 30205 18819
rect 30205 18785 30239 18819
rect 30239 18785 30248 18819
rect 30196 18776 30248 18785
rect 31024 18776 31076 18828
rect 29828 18751 29880 18760
rect 29828 18717 29837 18751
rect 29837 18717 29871 18751
rect 29871 18717 29880 18751
rect 29828 18708 29880 18717
rect 20076 18572 20128 18624
rect 21088 18572 21140 18624
rect 23572 18572 23624 18624
rect 26240 18640 26292 18692
rect 26976 18640 27028 18692
rect 27528 18683 27580 18692
rect 27528 18649 27537 18683
rect 27537 18649 27571 18683
rect 27571 18649 27580 18683
rect 27528 18640 27580 18649
rect 28908 18640 28960 18692
rect 27896 18572 27948 18624
rect 28724 18572 28776 18624
rect 29828 18572 29880 18624
rect 6286 18470 6338 18522
rect 6350 18470 6402 18522
rect 6414 18470 6466 18522
rect 6478 18470 6530 18522
rect 6542 18470 6594 18522
rect 13646 18470 13698 18522
rect 13710 18470 13762 18522
rect 13774 18470 13826 18522
rect 13838 18470 13890 18522
rect 13902 18470 13954 18522
rect 21006 18470 21058 18522
rect 21070 18470 21122 18522
rect 21134 18470 21186 18522
rect 21198 18470 21250 18522
rect 21262 18470 21314 18522
rect 28366 18470 28418 18522
rect 28430 18470 28482 18522
rect 28494 18470 28546 18522
rect 28558 18470 28610 18522
rect 28622 18470 28674 18522
rect 4988 18368 5040 18420
rect 6092 18368 6144 18420
rect 6460 18368 6512 18420
rect 6920 18368 6972 18420
rect 8208 18368 8260 18420
rect 8760 18368 8812 18420
rect 9864 18411 9916 18420
rect 9864 18377 9873 18411
rect 9873 18377 9907 18411
rect 9907 18377 9916 18411
rect 9864 18368 9916 18377
rect 11888 18411 11940 18420
rect 11888 18377 11897 18411
rect 11897 18377 11931 18411
rect 11931 18377 11940 18411
rect 11888 18368 11940 18377
rect 12992 18368 13044 18420
rect 5172 18300 5224 18352
rect 5632 18232 5684 18284
rect 6092 18232 6144 18284
rect 6368 18232 6420 18284
rect 6184 18164 6236 18216
rect 6920 18232 6972 18284
rect 9680 18300 9732 18352
rect 14372 18368 14424 18420
rect 14740 18368 14792 18420
rect 15476 18368 15528 18420
rect 15844 18368 15896 18420
rect 16488 18300 16540 18352
rect 7932 18275 7984 18284
rect 7932 18241 7941 18275
rect 7941 18241 7975 18275
rect 7975 18241 7984 18275
rect 7932 18232 7984 18241
rect 8392 18232 8444 18284
rect 10048 18164 10100 18216
rect 4068 18096 4120 18148
rect 8392 18096 8444 18148
rect 9128 18096 9180 18148
rect 10600 18164 10652 18216
rect 10968 18096 11020 18148
rect 7196 18028 7248 18080
rect 7380 18028 7432 18080
rect 7472 18028 7524 18080
rect 7656 18071 7708 18080
rect 7656 18037 7665 18071
rect 7665 18037 7699 18071
rect 7699 18037 7708 18071
rect 7656 18028 7708 18037
rect 10140 18028 10192 18080
rect 11520 18071 11572 18080
rect 11520 18037 11529 18071
rect 11529 18037 11563 18071
rect 11563 18037 11572 18071
rect 11520 18028 11572 18037
rect 12072 18028 12124 18080
rect 14648 18164 14700 18216
rect 12532 18096 12584 18148
rect 12624 18139 12676 18148
rect 12624 18105 12633 18139
rect 12633 18105 12667 18139
rect 12667 18105 12676 18139
rect 12624 18096 12676 18105
rect 13084 18096 13136 18148
rect 16028 18207 16080 18216
rect 16028 18173 16037 18207
rect 16037 18173 16071 18207
rect 16071 18173 16080 18207
rect 16028 18164 16080 18173
rect 16212 18164 16264 18216
rect 16488 18207 16540 18216
rect 16488 18173 16497 18207
rect 16497 18173 16531 18207
rect 16531 18173 16540 18207
rect 16488 18164 16540 18173
rect 12716 18028 12768 18080
rect 12992 18028 13044 18080
rect 15844 18096 15896 18148
rect 14924 18028 14976 18080
rect 15752 18028 15804 18080
rect 16396 18071 16448 18080
rect 16396 18037 16405 18071
rect 16405 18037 16439 18071
rect 16439 18037 16448 18071
rect 16396 18028 16448 18037
rect 16856 18207 16908 18216
rect 16856 18173 16865 18207
rect 16865 18173 16899 18207
rect 16899 18173 16908 18207
rect 16856 18164 16908 18173
rect 17776 18368 17828 18420
rect 18328 18368 18380 18420
rect 23480 18411 23532 18420
rect 23480 18377 23489 18411
rect 23489 18377 23523 18411
rect 23523 18377 23532 18411
rect 23480 18368 23532 18377
rect 23664 18368 23716 18420
rect 23848 18368 23900 18420
rect 23940 18368 23992 18420
rect 24400 18368 24452 18420
rect 24584 18411 24636 18420
rect 24584 18377 24593 18411
rect 24593 18377 24627 18411
rect 24627 18377 24636 18411
rect 24584 18368 24636 18377
rect 25596 18368 25648 18420
rect 25688 18368 25740 18420
rect 26516 18368 26568 18420
rect 27436 18368 27488 18420
rect 19064 18343 19116 18352
rect 19064 18309 19073 18343
rect 19073 18309 19107 18343
rect 19107 18309 19116 18343
rect 19064 18300 19116 18309
rect 19156 18300 19208 18352
rect 19432 18300 19484 18352
rect 19616 18232 19668 18284
rect 20628 18232 20680 18284
rect 26056 18232 26108 18284
rect 26792 18275 26844 18284
rect 26792 18241 26801 18275
rect 26801 18241 26835 18275
rect 26835 18241 26844 18275
rect 26792 18232 26844 18241
rect 26884 18275 26936 18284
rect 26884 18241 26893 18275
rect 26893 18241 26927 18275
rect 26927 18241 26936 18275
rect 26884 18232 26936 18241
rect 30288 18232 30340 18284
rect 19524 18164 19576 18216
rect 19800 18164 19852 18216
rect 19984 18207 20036 18216
rect 19984 18173 19993 18207
rect 19993 18173 20027 18207
rect 20027 18173 20036 18207
rect 19984 18164 20036 18173
rect 20076 18207 20128 18216
rect 20076 18173 20085 18207
rect 20085 18173 20119 18207
rect 20119 18173 20128 18207
rect 20076 18164 20128 18173
rect 20260 18207 20312 18216
rect 20260 18173 20269 18207
rect 20269 18173 20303 18207
rect 20303 18173 20312 18207
rect 20260 18164 20312 18173
rect 22560 18207 22612 18216
rect 22560 18173 22569 18207
rect 22569 18173 22603 18207
rect 22603 18173 22612 18207
rect 22560 18164 22612 18173
rect 19432 18139 19484 18148
rect 19432 18105 19441 18139
rect 19441 18105 19475 18139
rect 19475 18105 19484 18139
rect 19432 18096 19484 18105
rect 20352 18096 20404 18148
rect 22836 18096 22888 18148
rect 16856 18028 16908 18080
rect 17040 18071 17092 18080
rect 17040 18037 17049 18071
rect 17049 18037 17083 18071
rect 17083 18037 17092 18071
rect 17040 18028 17092 18037
rect 17316 18028 17368 18080
rect 19248 18028 19300 18080
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 22008 18028 22060 18080
rect 23112 18028 23164 18080
rect 23848 18207 23900 18216
rect 23848 18173 23857 18207
rect 23857 18173 23891 18207
rect 23891 18173 23900 18207
rect 23848 18164 23900 18173
rect 24492 18164 24544 18216
rect 24952 18207 25004 18216
rect 24952 18173 24961 18207
rect 24961 18173 24995 18207
rect 24995 18173 25004 18207
rect 24952 18164 25004 18173
rect 25320 18207 25372 18216
rect 25320 18173 25329 18207
rect 25329 18173 25363 18207
rect 25363 18173 25372 18207
rect 25320 18164 25372 18173
rect 25964 18164 26016 18216
rect 26424 18207 26476 18216
rect 26424 18173 26433 18207
rect 26433 18173 26467 18207
rect 26467 18173 26476 18207
rect 26424 18164 26476 18173
rect 27528 18164 27580 18216
rect 29460 18164 29512 18216
rect 30380 18096 30432 18148
rect 30748 18096 30800 18148
rect 25780 18028 25832 18080
rect 28080 18071 28132 18080
rect 28080 18037 28089 18071
rect 28089 18037 28123 18071
rect 28123 18037 28132 18071
rect 28080 18028 28132 18037
rect 6946 17926 6998 17978
rect 7010 17926 7062 17978
rect 7074 17926 7126 17978
rect 7138 17926 7190 17978
rect 7202 17926 7254 17978
rect 14306 17926 14358 17978
rect 14370 17926 14422 17978
rect 14434 17926 14486 17978
rect 14498 17926 14550 17978
rect 14562 17926 14614 17978
rect 21666 17926 21718 17978
rect 21730 17926 21782 17978
rect 21794 17926 21846 17978
rect 21858 17926 21910 17978
rect 21922 17926 21974 17978
rect 29026 17926 29078 17978
rect 29090 17926 29142 17978
rect 29154 17926 29206 17978
rect 29218 17926 29270 17978
rect 29282 17926 29334 17978
rect 7288 17824 7340 17876
rect 7932 17756 7984 17808
rect 7380 17688 7432 17740
rect 9772 17824 9824 17876
rect 8852 17756 8904 17808
rect 10140 17799 10192 17808
rect 10140 17765 10149 17799
rect 10149 17765 10183 17799
rect 10183 17765 10192 17799
rect 10140 17756 10192 17765
rect 10508 17756 10560 17808
rect 11888 17824 11940 17876
rect 12624 17824 12676 17876
rect 12716 17824 12768 17876
rect 9680 17688 9732 17740
rect 13176 17799 13228 17808
rect 12440 17688 12492 17740
rect 13176 17765 13185 17799
rect 13185 17765 13219 17799
rect 13219 17765 13228 17799
rect 13176 17756 13228 17765
rect 13268 17756 13320 17808
rect 14832 17824 14884 17876
rect 16304 17824 16356 17876
rect 22560 17824 22612 17876
rect 22836 17867 22888 17876
rect 22836 17833 22845 17867
rect 22845 17833 22879 17867
rect 22879 17833 22888 17867
rect 22836 17824 22888 17833
rect 23848 17824 23900 17876
rect 25320 17824 25372 17876
rect 25688 17824 25740 17876
rect 14648 17756 14700 17808
rect 15016 17756 15068 17808
rect 16396 17756 16448 17808
rect 13544 17688 13596 17740
rect 8300 17663 8352 17672
rect 8300 17629 8309 17663
rect 8309 17629 8343 17663
rect 8343 17629 8352 17663
rect 8300 17620 8352 17629
rect 10140 17620 10192 17672
rect 7840 17595 7892 17604
rect 7840 17561 7849 17595
rect 7849 17561 7883 17595
rect 7883 17561 7892 17595
rect 7840 17552 7892 17561
rect 11980 17620 12032 17672
rect 14004 17620 14056 17672
rect 14188 17620 14240 17672
rect 14740 17688 14792 17740
rect 15752 17731 15804 17740
rect 15752 17697 15761 17731
rect 15761 17697 15795 17731
rect 15795 17697 15804 17731
rect 15752 17688 15804 17697
rect 12072 17552 12124 17604
rect 11520 17484 11572 17536
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 13452 17552 13504 17604
rect 15660 17620 15712 17672
rect 15476 17552 15528 17604
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 14004 17527 14056 17536
rect 14004 17493 14013 17527
rect 14013 17493 14047 17527
rect 14047 17493 14056 17527
rect 14004 17484 14056 17493
rect 14096 17484 14148 17536
rect 14372 17484 14424 17536
rect 14464 17484 14516 17536
rect 16120 17688 16172 17740
rect 16672 17756 16724 17808
rect 18052 17756 18104 17808
rect 19064 17756 19116 17808
rect 22008 17756 22060 17808
rect 24308 17756 24360 17808
rect 25044 17756 25096 17808
rect 16948 17731 17000 17740
rect 16948 17697 16957 17731
rect 16957 17697 16991 17731
rect 16991 17697 17000 17731
rect 16948 17688 17000 17697
rect 17592 17731 17644 17740
rect 17592 17697 17601 17731
rect 17601 17697 17635 17731
rect 17635 17697 17644 17731
rect 17592 17688 17644 17697
rect 17132 17663 17184 17672
rect 17132 17629 17141 17663
rect 17141 17629 17175 17663
rect 17175 17629 17184 17663
rect 17132 17620 17184 17629
rect 16488 17552 16540 17604
rect 16856 17552 16908 17604
rect 17224 17552 17276 17604
rect 17684 17552 17736 17604
rect 17960 17620 18012 17672
rect 19432 17688 19484 17740
rect 20628 17688 20680 17740
rect 28724 17824 28776 17876
rect 28816 17867 28868 17876
rect 28816 17833 28825 17867
rect 28825 17833 28859 17867
rect 28859 17833 28868 17867
rect 28816 17824 28868 17833
rect 27896 17756 27948 17808
rect 28080 17756 28132 17808
rect 28908 17756 28960 17808
rect 25688 17688 25740 17740
rect 26884 17688 26936 17740
rect 19616 17620 19668 17672
rect 21272 17620 21324 17672
rect 22100 17620 22152 17672
rect 23572 17620 23624 17672
rect 23756 17663 23808 17672
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 25412 17620 25464 17672
rect 26792 17620 26844 17672
rect 29000 17620 29052 17672
rect 29368 17620 29420 17672
rect 29920 17731 29972 17740
rect 29920 17697 29929 17731
rect 29929 17697 29963 17731
rect 29963 17697 29972 17731
rect 29920 17688 29972 17697
rect 30840 17688 30892 17740
rect 33140 17620 33192 17672
rect 18144 17552 18196 17604
rect 17316 17484 17368 17536
rect 17868 17484 17920 17536
rect 17960 17527 18012 17536
rect 17960 17493 17969 17527
rect 17969 17493 18003 17527
rect 18003 17493 18012 17527
rect 17960 17484 18012 17493
rect 18236 17484 18288 17536
rect 20076 17527 20128 17536
rect 20076 17493 20085 17527
rect 20085 17493 20119 17527
rect 20119 17493 20128 17527
rect 20076 17484 20128 17493
rect 26332 17527 26384 17536
rect 26332 17493 26341 17527
rect 26341 17493 26375 17527
rect 26375 17493 26384 17527
rect 26332 17484 26384 17493
rect 29552 17527 29604 17536
rect 29552 17493 29561 17527
rect 29561 17493 29595 17527
rect 29595 17493 29604 17527
rect 29552 17484 29604 17493
rect 6286 17382 6338 17434
rect 6350 17382 6402 17434
rect 6414 17382 6466 17434
rect 6478 17382 6530 17434
rect 6542 17382 6594 17434
rect 13646 17382 13698 17434
rect 13710 17382 13762 17434
rect 13774 17382 13826 17434
rect 13838 17382 13890 17434
rect 13902 17382 13954 17434
rect 21006 17382 21058 17434
rect 21070 17382 21122 17434
rect 21134 17382 21186 17434
rect 21198 17382 21250 17434
rect 21262 17382 21314 17434
rect 28366 17382 28418 17434
rect 28430 17382 28482 17434
rect 28494 17382 28546 17434
rect 28558 17382 28610 17434
rect 28622 17382 28674 17434
rect 8300 17280 8352 17332
rect 10600 17280 10652 17332
rect 11704 17280 11756 17332
rect 12992 17280 13044 17332
rect 13268 17323 13320 17332
rect 13268 17289 13277 17323
rect 13277 17289 13311 17323
rect 13311 17289 13320 17323
rect 13268 17280 13320 17289
rect 13544 17280 13596 17332
rect 8116 17144 8168 17196
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 10048 17144 10100 17196
rect 12164 17144 12216 17196
rect 7288 17076 7340 17128
rect 9680 17076 9732 17128
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 12256 17119 12308 17128
rect 12256 17085 12265 17119
rect 12265 17085 12299 17119
rect 12299 17085 12308 17119
rect 12256 17076 12308 17085
rect 12348 17119 12400 17128
rect 12348 17085 12358 17119
rect 12358 17085 12392 17119
rect 12392 17085 12400 17119
rect 12348 17076 12400 17085
rect 8484 17008 8536 17060
rect 9956 17008 10008 17060
rect 11520 17008 11572 17060
rect 14004 17280 14056 17332
rect 14372 17280 14424 17332
rect 16028 17280 16080 17332
rect 16212 17280 16264 17332
rect 16396 17280 16448 17332
rect 17592 17280 17644 17332
rect 20628 17280 20680 17332
rect 25044 17280 25096 17332
rect 28908 17280 28960 17332
rect 29460 17280 29512 17332
rect 29920 17280 29972 17332
rect 14556 17212 14608 17264
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 14280 17144 14332 17196
rect 16120 17212 16172 17264
rect 17960 17212 18012 17264
rect 18144 17212 18196 17264
rect 13544 17119 13596 17128
rect 13544 17085 13553 17119
rect 13553 17085 13587 17119
rect 13587 17085 13596 17119
rect 13544 17076 13596 17085
rect 14004 17076 14056 17128
rect 14464 17119 14516 17128
rect 14464 17085 14487 17119
rect 14487 17085 14516 17119
rect 14464 17076 14516 17085
rect 15016 17144 15068 17196
rect 10232 16940 10284 16992
rect 11980 16940 12032 16992
rect 12624 16983 12676 16992
rect 12624 16949 12633 16983
rect 12633 16949 12667 16983
rect 12667 16949 12676 16983
rect 12624 16940 12676 16949
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 13544 16940 13596 16992
rect 14924 17119 14976 17128
rect 14924 17085 14933 17119
rect 14933 17085 14967 17119
rect 14967 17085 14976 17119
rect 14924 17076 14976 17085
rect 15108 17076 15160 17128
rect 15752 17144 15804 17196
rect 16304 17144 16356 17196
rect 17040 17144 17092 17196
rect 17132 17144 17184 17196
rect 18052 17144 18104 17196
rect 16580 17076 16632 17128
rect 16764 17119 16816 17128
rect 16764 17085 16773 17119
rect 16773 17085 16807 17119
rect 16807 17085 16816 17119
rect 16764 17076 16816 17085
rect 17316 17076 17368 17128
rect 17592 17119 17644 17128
rect 17592 17085 17601 17119
rect 17601 17085 17635 17119
rect 17635 17085 17644 17119
rect 17592 17076 17644 17085
rect 19340 17144 19392 17196
rect 22100 17144 22152 17196
rect 29000 17144 29052 17196
rect 17040 17051 17092 17060
rect 17040 17017 17049 17051
rect 17049 17017 17083 17051
rect 17083 17017 17092 17051
rect 17040 17008 17092 17017
rect 18512 17076 18564 17128
rect 19248 17076 19300 17128
rect 21456 17076 21508 17128
rect 23112 17076 23164 17128
rect 18052 17051 18104 17060
rect 18052 17017 18061 17051
rect 18061 17017 18095 17051
rect 18095 17017 18104 17051
rect 18052 17008 18104 17017
rect 20352 17051 20404 17060
rect 20352 17017 20361 17051
rect 20361 17017 20395 17051
rect 20395 17017 20404 17051
rect 20352 17008 20404 17017
rect 14832 16940 14884 16992
rect 15016 16940 15068 16992
rect 15292 16940 15344 16992
rect 15384 16940 15436 16992
rect 15936 16940 15988 16992
rect 16672 16940 16724 16992
rect 17316 16940 17368 16992
rect 17868 16940 17920 16992
rect 17960 16940 18012 16992
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 24952 17119 25004 17128
rect 24952 17085 24961 17119
rect 24961 17085 24995 17119
rect 24995 17085 25004 17119
rect 24952 17076 25004 17085
rect 23664 17008 23716 17060
rect 27344 17008 27396 17060
rect 25412 16983 25464 16992
rect 25412 16949 25421 16983
rect 25421 16949 25455 16983
rect 25455 16949 25464 16983
rect 25412 16940 25464 16949
rect 25504 16940 25556 16992
rect 26516 16940 26568 16992
rect 27068 16940 27120 16992
rect 30656 17119 30708 17128
rect 30656 17085 30665 17119
rect 30665 17085 30699 17119
rect 30699 17085 30708 17119
rect 30656 17076 30708 17085
rect 30932 17076 30984 17128
rect 28908 16940 28960 16992
rect 30380 16940 30432 16992
rect 6946 16838 6998 16890
rect 7010 16838 7062 16890
rect 7074 16838 7126 16890
rect 7138 16838 7190 16890
rect 7202 16838 7254 16890
rect 14306 16838 14358 16890
rect 14370 16838 14422 16890
rect 14434 16838 14486 16890
rect 14498 16838 14550 16890
rect 14562 16838 14614 16890
rect 21666 16838 21718 16890
rect 21730 16838 21782 16890
rect 21794 16838 21846 16890
rect 21858 16838 21910 16890
rect 21922 16838 21974 16890
rect 29026 16838 29078 16890
rect 29090 16838 29142 16890
rect 29154 16838 29206 16890
rect 29218 16838 29270 16890
rect 29282 16838 29334 16890
rect 7932 16736 7984 16788
rect 8300 16736 8352 16788
rect 8484 16736 8536 16788
rect 8852 16779 8904 16788
rect 8852 16745 8861 16779
rect 8861 16745 8895 16779
rect 8895 16745 8904 16779
rect 8852 16736 8904 16745
rect 9128 16779 9180 16788
rect 9128 16745 9137 16779
rect 9137 16745 9171 16779
rect 9171 16745 9180 16779
rect 9128 16736 9180 16745
rect 10968 16736 11020 16788
rect 5908 16643 5960 16652
rect 5908 16609 5917 16643
rect 5917 16609 5951 16643
rect 5951 16609 5960 16643
rect 5908 16600 5960 16609
rect 10140 16600 10192 16652
rect 10968 16643 11020 16652
rect 10968 16609 10977 16643
rect 10977 16609 11011 16643
rect 11011 16609 11020 16643
rect 10968 16600 11020 16609
rect 11612 16600 11664 16652
rect 11704 16600 11756 16652
rect 13084 16736 13136 16788
rect 14096 16779 14148 16788
rect 14096 16745 14105 16779
rect 14105 16745 14139 16779
rect 14139 16745 14148 16779
rect 14096 16736 14148 16745
rect 14832 16736 14884 16788
rect 15568 16736 15620 16788
rect 12808 16600 12860 16652
rect 13360 16600 13412 16652
rect 14004 16668 14056 16720
rect 11520 16532 11572 16584
rect 15200 16600 15252 16652
rect 6736 16507 6788 16516
rect 6736 16473 6745 16507
rect 6745 16473 6779 16507
rect 6779 16473 6788 16507
rect 6736 16464 6788 16473
rect 5264 16439 5316 16448
rect 5264 16405 5273 16439
rect 5273 16405 5307 16439
rect 5307 16405 5316 16439
rect 5264 16396 5316 16405
rect 10416 16464 10468 16516
rect 12072 16464 12124 16516
rect 12164 16464 12216 16516
rect 12532 16396 12584 16448
rect 12624 16396 12676 16448
rect 15752 16575 15804 16584
rect 15752 16541 15761 16575
rect 15761 16541 15795 16575
rect 15795 16541 15804 16575
rect 16488 16736 16540 16788
rect 20076 16736 20128 16788
rect 21272 16736 21324 16788
rect 17592 16668 17644 16720
rect 16212 16600 16264 16652
rect 16580 16600 16632 16652
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 15752 16532 15804 16541
rect 17776 16668 17828 16720
rect 17316 16532 17368 16584
rect 19432 16600 19484 16652
rect 19524 16600 19576 16652
rect 22836 16779 22888 16788
rect 22836 16745 22845 16779
rect 22845 16745 22879 16779
rect 22879 16745 22888 16779
rect 22836 16736 22888 16745
rect 26332 16736 26384 16788
rect 27068 16779 27120 16788
rect 27068 16745 27077 16779
rect 27077 16745 27111 16779
rect 27111 16745 27120 16779
rect 27068 16736 27120 16745
rect 27344 16779 27396 16788
rect 27344 16745 27353 16779
rect 27353 16745 27387 16779
rect 27387 16745 27396 16779
rect 27344 16736 27396 16745
rect 30656 16736 30708 16788
rect 26516 16668 26568 16720
rect 28908 16668 28960 16720
rect 29552 16668 29604 16720
rect 31300 16668 31352 16720
rect 17868 16532 17920 16584
rect 16948 16464 17000 16516
rect 15568 16396 15620 16448
rect 15660 16396 15712 16448
rect 15936 16396 15988 16448
rect 16120 16396 16172 16448
rect 19984 16575 20036 16584
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 19984 16532 20036 16541
rect 17408 16439 17460 16448
rect 17408 16405 17417 16439
rect 17417 16405 17451 16439
rect 17451 16405 17460 16439
rect 17408 16396 17460 16405
rect 18420 16396 18472 16448
rect 29368 16575 29420 16584
rect 29368 16541 29377 16575
rect 29377 16541 29411 16575
rect 29411 16541 29420 16575
rect 29368 16532 29420 16541
rect 31852 16575 31904 16584
rect 31852 16541 31861 16575
rect 31861 16541 31895 16575
rect 31895 16541 31904 16575
rect 31852 16532 31904 16541
rect 30840 16464 30892 16516
rect 30380 16396 30432 16448
rect 6286 16294 6338 16346
rect 6350 16294 6402 16346
rect 6414 16294 6466 16346
rect 6478 16294 6530 16346
rect 6542 16294 6594 16346
rect 13646 16294 13698 16346
rect 13710 16294 13762 16346
rect 13774 16294 13826 16346
rect 13838 16294 13890 16346
rect 13902 16294 13954 16346
rect 21006 16294 21058 16346
rect 21070 16294 21122 16346
rect 21134 16294 21186 16346
rect 21198 16294 21250 16346
rect 21262 16294 21314 16346
rect 28366 16294 28418 16346
rect 28430 16294 28482 16346
rect 28494 16294 28546 16346
rect 28558 16294 28610 16346
rect 28622 16294 28674 16346
rect 12164 16192 12216 16244
rect 13084 16235 13136 16244
rect 13084 16201 13093 16235
rect 13093 16201 13127 16235
rect 13127 16201 13136 16235
rect 13084 16192 13136 16201
rect 13176 16192 13228 16244
rect 14188 16235 14240 16244
rect 14188 16201 14197 16235
rect 14197 16201 14231 16235
rect 14231 16201 14240 16235
rect 14188 16192 14240 16201
rect 5632 16056 5684 16108
rect 6644 16056 6696 16108
rect 1308 15920 1360 15972
rect 6736 15988 6788 16040
rect 5816 15920 5868 15972
rect 6184 15920 6236 15972
rect 8484 16031 8536 16040
rect 8484 15997 8493 16031
rect 8493 15997 8527 16031
rect 8527 15997 8536 16031
rect 8484 15988 8536 15997
rect 10968 15988 11020 16040
rect 12348 16124 12400 16176
rect 12532 16167 12584 16176
rect 12532 16133 12541 16167
rect 12541 16133 12575 16167
rect 12575 16133 12584 16167
rect 12532 16124 12584 16133
rect 15016 16192 15068 16244
rect 15476 16235 15528 16244
rect 15476 16201 15485 16235
rect 15485 16201 15519 16235
rect 15519 16201 15528 16235
rect 15476 16192 15528 16201
rect 16672 16192 16724 16244
rect 17408 16192 17460 16244
rect 17684 16192 17736 16244
rect 19984 16192 20036 16244
rect 12072 16056 12124 16108
rect 8576 15963 8628 15972
rect 8576 15929 8585 15963
rect 8585 15929 8619 15963
rect 8619 15929 8628 15963
rect 8576 15920 8628 15929
rect 10416 15920 10468 15972
rect 3424 15852 3476 15904
rect 5448 15852 5500 15904
rect 6828 15852 6880 15904
rect 7564 15895 7616 15904
rect 7564 15861 7573 15895
rect 7573 15861 7607 15895
rect 7607 15861 7616 15895
rect 7564 15852 7616 15861
rect 7932 15852 7984 15904
rect 10692 15852 10744 15904
rect 11888 15988 11940 16040
rect 12440 15988 12492 16040
rect 13452 16056 13504 16108
rect 17132 16167 17184 16176
rect 17132 16133 17141 16167
rect 17141 16133 17175 16167
rect 17175 16133 17184 16167
rect 17132 16124 17184 16133
rect 19800 16124 19852 16176
rect 23112 16124 23164 16176
rect 14648 16099 14700 16108
rect 14648 16065 14657 16099
rect 14657 16065 14691 16099
rect 14691 16065 14700 16099
rect 14648 16056 14700 16065
rect 15292 16056 15344 16108
rect 12624 15988 12676 16040
rect 13360 15988 13412 16040
rect 14004 15988 14056 16040
rect 13544 15920 13596 15972
rect 14648 15920 14700 15972
rect 15476 15988 15528 16040
rect 15660 15988 15712 16040
rect 16856 16056 16908 16108
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 20904 16056 20956 16108
rect 11520 15895 11572 15904
rect 11520 15861 11529 15895
rect 11529 15861 11563 15895
rect 11563 15861 11572 15895
rect 11520 15852 11572 15861
rect 12348 15852 12400 15904
rect 15016 15852 15068 15904
rect 16580 15988 16632 16040
rect 16672 15988 16724 16040
rect 18144 16031 18196 16040
rect 18144 15997 18153 16031
rect 18153 15997 18187 16031
rect 18187 15997 18196 16031
rect 18144 15988 18196 15997
rect 30012 16192 30064 16244
rect 31852 16235 31904 16244
rect 31852 16201 31861 16235
rect 31861 16201 31895 16235
rect 31895 16201 31904 16235
rect 31852 16192 31904 16201
rect 25504 16056 25556 16108
rect 29368 16056 29420 16108
rect 16304 15920 16356 15972
rect 17776 15920 17828 15972
rect 19156 15920 19208 15972
rect 17040 15852 17092 15904
rect 24124 16031 24176 16040
rect 24124 15997 24133 16031
rect 24133 15997 24167 16031
rect 24167 15997 24176 16031
rect 24124 15988 24176 15997
rect 26608 15988 26660 16040
rect 29828 16056 29880 16108
rect 30196 15920 30248 15972
rect 24400 15852 24452 15904
rect 24584 15852 24636 15904
rect 26332 15895 26384 15904
rect 26332 15861 26341 15895
rect 26341 15861 26375 15895
rect 26375 15861 26384 15895
rect 26332 15852 26384 15861
rect 6946 15750 6998 15802
rect 7010 15750 7062 15802
rect 7074 15750 7126 15802
rect 7138 15750 7190 15802
rect 7202 15750 7254 15802
rect 14306 15750 14358 15802
rect 14370 15750 14422 15802
rect 14434 15750 14486 15802
rect 14498 15750 14550 15802
rect 14562 15750 14614 15802
rect 21666 15750 21718 15802
rect 21730 15750 21782 15802
rect 21794 15750 21846 15802
rect 21858 15750 21910 15802
rect 21922 15750 21974 15802
rect 29026 15750 29078 15802
rect 29090 15750 29142 15802
rect 29154 15750 29206 15802
rect 29218 15750 29270 15802
rect 29282 15750 29334 15802
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 5448 15648 5500 15700
rect 5264 15580 5316 15632
rect 6828 15648 6880 15700
rect 12256 15648 12308 15700
rect 12348 15648 12400 15700
rect 12164 15580 12216 15632
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 11152 15555 11204 15564
rect 11152 15521 11161 15555
rect 11161 15521 11195 15555
rect 11195 15521 11204 15555
rect 11152 15512 11204 15521
rect 12348 15512 12400 15564
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 12808 15555 12860 15564
rect 12808 15521 12817 15555
rect 12817 15521 12851 15555
rect 12851 15521 12860 15555
rect 12808 15512 12860 15521
rect 12900 15555 12952 15564
rect 12900 15521 12909 15555
rect 12909 15521 12943 15555
rect 12943 15521 12952 15555
rect 12900 15512 12952 15521
rect 5448 15444 5500 15496
rect 7288 15444 7340 15496
rect 7656 15487 7708 15496
rect 7656 15453 7665 15487
rect 7665 15453 7699 15487
rect 7699 15453 7708 15487
rect 7656 15444 7708 15453
rect 9036 15487 9088 15496
rect 9036 15453 9045 15487
rect 9045 15453 9079 15487
rect 9079 15453 9088 15487
rect 9036 15444 9088 15453
rect 11796 15444 11848 15496
rect 12532 15444 12584 15496
rect 13176 15648 13228 15700
rect 14188 15648 14240 15700
rect 14648 15648 14700 15700
rect 15292 15648 15344 15700
rect 17500 15648 17552 15700
rect 19156 15648 19208 15700
rect 13268 15623 13320 15632
rect 13268 15589 13277 15623
rect 13277 15589 13311 15623
rect 13311 15589 13320 15623
rect 13268 15580 13320 15589
rect 14004 15555 14056 15564
rect 14004 15521 14013 15555
rect 14013 15521 14047 15555
rect 14047 15521 14056 15555
rect 14004 15512 14056 15521
rect 14096 15512 14148 15564
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 15660 15580 15712 15632
rect 14832 15512 14884 15564
rect 15200 15444 15252 15496
rect 15384 15555 15436 15564
rect 15384 15521 15393 15555
rect 15393 15521 15427 15555
rect 15427 15521 15436 15555
rect 15384 15512 15436 15521
rect 15568 15555 15620 15564
rect 15568 15521 15577 15555
rect 15577 15521 15611 15555
rect 15611 15521 15620 15555
rect 15568 15512 15620 15521
rect 16120 15512 16172 15564
rect 16672 15555 16724 15564
rect 16672 15521 16681 15555
rect 16681 15521 16715 15555
rect 16715 15521 16724 15555
rect 16672 15512 16724 15521
rect 17040 15580 17092 15632
rect 17224 15512 17276 15564
rect 15844 15444 15896 15496
rect 16580 15444 16632 15496
rect 15568 15376 15620 15428
rect 5724 15308 5776 15360
rect 8576 15308 8628 15360
rect 8944 15308 8996 15360
rect 10692 15308 10744 15360
rect 10968 15308 11020 15360
rect 11796 15308 11848 15360
rect 11980 15308 12032 15360
rect 12164 15308 12216 15360
rect 14004 15351 14056 15360
rect 14004 15317 14013 15351
rect 14013 15317 14047 15351
rect 14047 15317 14056 15351
rect 14004 15308 14056 15317
rect 14188 15308 14240 15360
rect 15476 15308 15528 15360
rect 23112 15648 23164 15700
rect 24124 15648 24176 15700
rect 24400 15648 24452 15700
rect 30196 15691 30248 15700
rect 30196 15657 30205 15691
rect 30205 15657 30239 15691
rect 30239 15657 30248 15691
rect 30196 15648 30248 15657
rect 30472 15648 30524 15700
rect 21548 15580 21600 15632
rect 23572 15580 23624 15632
rect 20536 15444 20588 15496
rect 17592 15376 17644 15428
rect 19156 15376 19208 15428
rect 17500 15308 17552 15360
rect 23112 15512 23164 15564
rect 24584 15555 24636 15564
rect 24584 15521 24593 15555
rect 24593 15521 24627 15555
rect 24627 15521 24636 15555
rect 24584 15512 24636 15521
rect 26056 15580 26108 15632
rect 27804 15580 27856 15632
rect 30748 15580 30800 15632
rect 33140 15580 33192 15632
rect 26884 15444 26936 15496
rect 30380 15512 30432 15564
rect 19524 15308 19576 15360
rect 19800 15351 19852 15360
rect 19800 15317 19809 15351
rect 19809 15317 19843 15351
rect 19843 15317 19852 15351
rect 19800 15308 19852 15317
rect 19892 15308 19944 15360
rect 21364 15308 21416 15360
rect 22468 15308 22520 15360
rect 24584 15308 24636 15360
rect 27988 15308 28040 15360
rect 28172 15308 28224 15360
rect 6286 15206 6338 15258
rect 6350 15206 6402 15258
rect 6414 15206 6466 15258
rect 6478 15206 6530 15258
rect 6542 15206 6594 15258
rect 13646 15206 13698 15258
rect 13710 15206 13762 15258
rect 13774 15206 13826 15258
rect 13838 15206 13890 15258
rect 13902 15206 13954 15258
rect 21006 15206 21058 15258
rect 21070 15206 21122 15258
rect 21134 15206 21186 15258
rect 21198 15206 21250 15258
rect 21262 15206 21314 15258
rect 28366 15206 28418 15258
rect 28430 15206 28482 15258
rect 28494 15206 28546 15258
rect 28558 15206 28610 15258
rect 28622 15206 28674 15258
rect 5908 15104 5960 15156
rect 7380 15104 7432 15156
rect 9036 15104 9088 15156
rect 9220 15104 9272 15156
rect 9956 15104 10008 15156
rect 11980 15104 12032 15156
rect 12808 15104 12860 15156
rect 12900 15104 12952 15156
rect 13452 15104 13504 15156
rect 15384 15147 15436 15156
rect 15384 15113 15393 15147
rect 15393 15113 15427 15147
rect 15427 15113 15436 15147
rect 15384 15104 15436 15113
rect 16856 15147 16908 15156
rect 16856 15113 16865 15147
rect 16865 15113 16899 15147
rect 16899 15113 16908 15147
rect 16856 15104 16908 15113
rect 17040 15147 17092 15156
rect 17040 15113 17049 15147
rect 17049 15113 17083 15147
rect 17083 15113 17092 15147
rect 17040 15104 17092 15113
rect 17960 15104 18012 15156
rect 19248 15104 19300 15156
rect 10876 15036 10928 15088
rect 12992 15036 13044 15088
rect 22560 15104 22612 15156
rect 26884 15104 26936 15156
rect 31300 15147 31352 15156
rect 31300 15113 31309 15147
rect 31309 15113 31343 15147
rect 31343 15113 31352 15147
rect 31300 15104 31352 15113
rect 5632 15011 5684 15020
rect 5632 14977 5641 15011
rect 5641 14977 5675 15011
rect 5675 14977 5684 15011
rect 5632 14968 5684 14977
rect 5724 14968 5776 15020
rect 7288 14968 7340 15020
rect 10692 14968 10744 15020
rect 12532 14968 12584 15020
rect 5816 14943 5868 14952
rect 5816 14909 5825 14943
rect 5825 14909 5859 14943
rect 5859 14909 5868 14943
rect 5816 14900 5868 14909
rect 6092 14900 6144 14952
rect 11336 14900 11388 14952
rect 11520 14943 11572 14952
rect 11520 14909 11529 14943
rect 11529 14909 11563 14943
rect 11563 14909 11572 14943
rect 11520 14900 11572 14909
rect 11796 14900 11848 14952
rect 13084 14900 13136 14952
rect 13360 14943 13412 14952
rect 13360 14909 13369 14943
rect 13369 14909 13403 14943
rect 13403 14909 13412 14943
rect 13360 14900 13412 14909
rect 4252 14764 4304 14816
rect 4436 14807 4488 14816
rect 4436 14773 4445 14807
rect 4445 14773 4479 14807
rect 4479 14773 4488 14807
rect 4436 14764 4488 14773
rect 6552 14764 6604 14816
rect 7564 14832 7616 14884
rect 8024 14832 8076 14884
rect 11888 14832 11940 14884
rect 14648 14943 14700 14952
rect 14648 14909 14657 14943
rect 14657 14909 14691 14943
rect 14691 14909 14700 14943
rect 14648 14900 14700 14909
rect 14832 14943 14884 14952
rect 14832 14909 14841 14943
rect 14841 14909 14875 14943
rect 14875 14909 14884 14943
rect 14832 14900 14884 14909
rect 14924 14900 14976 14952
rect 15476 14900 15528 14952
rect 15844 14968 15896 15020
rect 16120 14943 16172 14952
rect 16120 14909 16129 14943
rect 16129 14909 16163 14943
rect 16163 14909 16172 14943
rect 16120 14900 16172 14909
rect 17592 14968 17644 15020
rect 9036 14764 9088 14816
rect 10784 14764 10836 14816
rect 11244 14764 11296 14816
rect 11336 14807 11388 14816
rect 11336 14773 11345 14807
rect 11345 14773 11379 14807
rect 11379 14773 11388 14807
rect 11336 14764 11388 14773
rect 12348 14764 12400 14816
rect 12808 14764 12860 14816
rect 13084 14764 13136 14816
rect 13544 14764 13596 14816
rect 15752 14764 15804 14816
rect 16120 14764 16172 14816
rect 16212 14764 16264 14816
rect 17500 14900 17552 14952
rect 16580 14832 16632 14884
rect 18144 14968 18196 15020
rect 19892 14968 19944 15020
rect 22192 14968 22244 15020
rect 22928 14968 22980 15020
rect 17684 14875 17736 14884
rect 17684 14841 17693 14875
rect 17693 14841 17727 14875
rect 17727 14841 17736 14875
rect 17684 14832 17736 14841
rect 17224 14764 17276 14816
rect 17408 14764 17460 14816
rect 17960 14807 18012 14816
rect 17960 14773 17969 14807
rect 17969 14773 18003 14807
rect 18003 14773 18012 14807
rect 17960 14764 18012 14773
rect 18052 14764 18104 14816
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 20352 14900 20404 14952
rect 20628 14900 20680 14952
rect 18328 14832 18380 14884
rect 19524 14832 19576 14884
rect 20996 14764 21048 14816
rect 21456 14764 21508 14816
rect 21548 14764 21600 14816
rect 22008 14764 22060 14816
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 22560 14943 22612 14952
rect 22560 14909 22569 14943
rect 22569 14909 22603 14943
rect 22603 14909 22612 14943
rect 22560 14900 22612 14909
rect 24308 14943 24360 14952
rect 24308 14909 24317 14943
rect 24317 14909 24351 14943
rect 24351 14909 24360 14943
rect 24308 14900 24360 14909
rect 22836 14764 22888 14816
rect 23020 14807 23072 14816
rect 23020 14773 23029 14807
rect 23029 14773 23063 14807
rect 23063 14773 23072 14807
rect 23020 14764 23072 14773
rect 23204 14764 23256 14816
rect 24768 14807 24820 14816
rect 24768 14773 24777 14807
rect 24777 14773 24811 14807
rect 24811 14773 24820 14807
rect 24768 14764 24820 14773
rect 30932 15036 30984 15088
rect 26332 15011 26384 15020
rect 26332 14977 26341 15011
rect 26341 14977 26375 15011
rect 26375 14977 26384 15011
rect 26332 14968 26384 14977
rect 28080 14968 28132 15020
rect 25872 14900 25924 14952
rect 26056 14943 26108 14952
rect 26056 14909 26065 14943
rect 26065 14909 26099 14943
rect 26099 14909 26108 14943
rect 26056 14900 26108 14909
rect 28448 14943 28500 14952
rect 28448 14909 28457 14943
rect 28457 14909 28491 14943
rect 28491 14909 28500 14943
rect 28448 14900 28500 14909
rect 28632 14900 28684 14952
rect 29736 14900 29788 14952
rect 28540 14832 28592 14884
rect 30748 14900 30800 14952
rect 27896 14764 27948 14816
rect 29460 14764 29512 14816
rect 29920 14807 29972 14816
rect 29920 14773 29929 14807
rect 29929 14773 29963 14807
rect 29963 14773 29972 14807
rect 29920 14764 29972 14773
rect 30840 14832 30892 14884
rect 31668 14832 31720 14884
rect 30656 14764 30708 14816
rect 6946 14662 6998 14714
rect 7010 14662 7062 14714
rect 7074 14662 7126 14714
rect 7138 14662 7190 14714
rect 7202 14662 7254 14714
rect 14306 14662 14358 14714
rect 14370 14662 14422 14714
rect 14434 14662 14486 14714
rect 14498 14662 14550 14714
rect 14562 14662 14614 14714
rect 21666 14662 21718 14714
rect 21730 14662 21782 14714
rect 21794 14662 21846 14714
rect 21858 14662 21910 14714
rect 21922 14662 21974 14714
rect 29026 14662 29078 14714
rect 29090 14662 29142 14714
rect 29154 14662 29206 14714
rect 29218 14662 29270 14714
rect 29282 14662 29334 14714
rect 6184 14492 6236 14544
rect 6552 14560 6604 14612
rect 7656 14560 7708 14612
rect 8024 14560 8076 14612
rect 8484 14560 8536 14612
rect 8944 14603 8996 14612
rect 8944 14569 8953 14603
rect 8953 14569 8987 14603
rect 8987 14569 8996 14603
rect 8944 14560 8996 14569
rect 9864 14560 9916 14612
rect 10324 14560 10376 14612
rect 11152 14560 11204 14612
rect 7380 14535 7432 14544
rect 7380 14501 7389 14535
rect 7389 14501 7423 14535
rect 7423 14501 7432 14535
rect 7380 14492 7432 14501
rect 4436 14356 4488 14408
rect 5448 14356 5500 14408
rect 8024 14467 8076 14476
rect 8024 14433 8033 14467
rect 8033 14433 8067 14467
rect 8067 14433 8076 14467
rect 8024 14424 8076 14433
rect 7748 14331 7800 14340
rect 7748 14297 7757 14331
rect 7757 14297 7791 14331
rect 7791 14297 7800 14331
rect 7748 14288 7800 14297
rect 9036 14399 9088 14408
rect 9036 14365 9045 14399
rect 9045 14365 9079 14399
rect 9079 14365 9088 14399
rect 9036 14356 9088 14365
rect 9128 14356 9180 14408
rect 9680 14288 9732 14340
rect 4252 14220 4304 14272
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 10232 14220 10284 14272
rect 11152 14424 11204 14476
rect 11336 14535 11388 14544
rect 11336 14501 11345 14535
rect 11345 14501 11379 14535
rect 11379 14501 11388 14535
rect 12900 14560 12952 14612
rect 13268 14560 13320 14612
rect 13360 14560 13412 14612
rect 14004 14560 14056 14612
rect 14648 14560 14700 14612
rect 17040 14560 17092 14612
rect 11336 14492 11388 14501
rect 11428 14424 11480 14476
rect 11980 14467 12032 14476
rect 11980 14433 11989 14467
rect 11989 14433 12023 14467
rect 12023 14433 12032 14467
rect 11980 14424 12032 14433
rect 10876 14356 10928 14408
rect 11796 14356 11848 14408
rect 12624 14424 12676 14476
rect 13084 14424 13136 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 14648 14467 14700 14476
rect 14648 14433 14657 14467
rect 14657 14433 14691 14467
rect 14691 14433 14700 14467
rect 14648 14424 14700 14433
rect 14096 14356 14148 14408
rect 14556 14356 14608 14408
rect 15476 14492 15528 14544
rect 15844 14492 15896 14544
rect 17684 14560 17736 14612
rect 18696 14560 18748 14612
rect 20352 14560 20404 14612
rect 15568 14424 15620 14476
rect 16672 14424 16724 14476
rect 16948 14424 17000 14476
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 10692 14220 10744 14272
rect 11612 14263 11664 14272
rect 11612 14229 11621 14263
rect 11621 14229 11655 14263
rect 11655 14229 11664 14263
rect 11612 14220 11664 14229
rect 11888 14220 11940 14272
rect 17316 14424 17368 14476
rect 20904 14492 20956 14544
rect 20996 14535 21048 14544
rect 20996 14501 21005 14535
rect 21005 14501 21039 14535
rect 21039 14501 21048 14535
rect 20996 14492 21048 14501
rect 23020 14560 23072 14612
rect 23572 14603 23624 14612
rect 23572 14569 23581 14603
rect 23581 14569 23615 14603
rect 23615 14569 23624 14603
rect 23572 14560 23624 14569
rect 25872 14560 25924 14612
rect 18328 14424 18380 14476
rect 19156 14424 19208 14476
rect 20628 14424 20680 14476
rect 17500 14399 17552 14408
rect 17500 14365 17509 14399
rect 17509 14365 17543 14399
rect 17543 14365 17552 14399
rect 17500 14356 17552 14365
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 18880 14331 18932 14340
rect 14096 14220 14148 14272
rect 14832 14263 14884 14272
rect 14832 14229 14841 14263
rect 14841 14229 14875 14263
rect 14875 14229 14884 14263
rect 14832 14220 14884 14229
rect 14924 14220 14976 14272
rect 18880 14297 18889 14331
rect 18889 14297 18923 14331
rect 18923 14297 18932 14331
rect 18880 14288 18932 14297
rect 22928 14424 22980 14476
rect 23664 14467 23716 14476
rect 23664 14433 23673 14467
rect 23673 14433 23707 14467
rect 23707 14433 23716 14467
rect 23664 14424 23716 14433
rect 24032 14467 24084 14476
rect 24032 14433 24041 14467
rect 24041 14433 24075 14467
rect 24075 14433 24084 14467
rect 24032 14424 24084 14433
rect 26056 14492 26108 14544
rect 27160 14560 27212 14612
rect 27804 14560 27856 14612
rect 28448 14560 28500 14612
rect 28540 14560 28592 14612
rect 27528 14424 27580 14476
rect 27712 14467 27764 14476
rect 27712 14433 27721 14467
rect 27721 14433 27755 14467
rect 27755 14433 27764 14467
rect 27712 14424 27764 14433
rect 28816 14535 28868 14544
rect 28816 14501 28843 14535
rect 28843 14501 28868 14535
rect 28816 14492 28868 14501
rect 28632 14424 28684 14476
rect 20812 14356 20864 14408
rect 21364 14399 21416 14408
rect 21364 14365 21373 14399
rect 21373 14365 21407 14399
rect 21407 14365 21416 14399
rect 21364 14356 21416 14365
rect 20904 14288 20956 14340
rect 25412 14356 25464 14408
rect 25780 14399 25832 14408
rect 25780 14365 25789 14399
rect 25789 14365 25823 14399
rect 25823 14365 25832 14399
rect 25780 14356 25832 14365
rect 27620 14356 27672 14408
rect 27988 14356 28040 14408
rect 30288 14535 30340 14544
rect 30288 14501 30297 14535
rect 30297 14501 30331 14535
rect 30331 14501 30340 14535
rect 30288 14492 30340 14501
rect 30656 14467 30708 14476
rect 30656 14433 30665 14467
rect 30665 14433 30699 14467
rect 30699 14433 30708 14467
rect 30656 14424 30708 14433
rect 30840 14424 30892 14476
rect 29276 14399 29328 14408
rect 29276 14365 29285 14399
rect 29285 14365 29319 14399
rect 29319 14365 29328 14399
rect 29276 14356 29328 14365
rect 29920 14356 29972 14408
rect 31024 14356 31076 14408
rect 31300 14399 31352 14408
rect 31300 14365 31309 14399
rect 31309 14365 31343 14399
rect 31343 14365 31352 14399
rect 31300 14356 31352 14365
rect 33140 14356 33192 14408
rect 16580 14263 16632 14272
rect 16580 14229 16589 14263
rect 16589 14229 16623 14263
rect 16623 14229 16632 14263
rect 16580 14220 16632 14229
rect 17408 14220 17460 14272
rect 18604 14220 18656 14272
rect 18696 14263 18748 14272
rect 18696 14229 18705 14263
rect 18705 14229 18739 14263
rect 18739 14229 18748 14263
rect 18696 14220 18748 14229
rect 20076 14263 20128 14272
rect 20076 14229 20085 14263
rect 20085 14229 20119 14263
rect 20119 14229 20128 14263
rect 24308 14288 24360 14340
rect 27804 14288 27856 14340
rect 20076 14220 20128 14229
rect 22652 14220 22704 14272
rect 24768 14220 24820 14272
rect 26148 14220 26200 14272
rect 27344 14220 27396 14272
rect 28908 14288 28960 14340
rect 29644 14220 29696 14272
rect 30748 14263 30800 14272
rect 30748 14229 30757 14263
rect 30757 14229 30791 14263
rect 30791 14229 30800 14263
rect 30748 14220 30800 14229
rect 6286 14118 6338 14170
rect 6350 14118 6402 14170
rect 6414 14118 6466 14170
rect 6478 14118 6530 14170
rect 6542 14118 6594 14170
rect 13646 14118 13698 14170
rect 13710 14118 13762 14170
rect 13774 14118 13826 14170
rect 13838 14118 13890 14170
rect 13902 14118 13954 14170
rect 21006 14118 21058 14170
rect 21070 14118 21122 14170
rect 21134 14118 21186 14170
rect 21198 14118 21250 14170
rect 21262 14118 21314 14170
rect 28366 14118 28418 14170
rect 28430 14118 28482 14170
rect 28494 14118 28546 14170
rect 28558 14118 28610 14170
rect 28622 14118 28674 14170
rect 5632 14059 5684 14068
rect 5632 14025 5641 14059
rect 5641 14025 5675 14059
rect 5675 14025 5684 14059
rect 5632 14016 5684 14025
rect 6644 14016 6696 14068
rect 8484 14016 8536 14068
rect 9128 14016 9180 14068
rect 11060 14016 11112 14068
rect 12440 14016 12492 14068
rect 11336 13948 11388 14000
rect 13084 14016 13136 14068
rect 14648 14016 14700 14068
rect 14832 14016 14884 14068
rect 15108 14016 15160 14068
rect 17500 14059 17552 14068
rect 17500 14025 17509 14059
rect 17509 14025 17543 14059
rect 17543 14025 17552 14059
rect 17500 14016 17552 14025
rect 14280 13948 14332 14000
rect 1308 13880 1360 13932
rect 5448 13880 5500 13932
rect 7288 13880 7340 13932
rect 8208 13880 8260 13932
rect 10048 13880 10100 13932
rect 4252 13855 4304 13864
rect 4252 13821 4261 13855
rect 4261 13821 4295 13855
rect 4295 13821 4304 13855
rect 4252 13812 4304 13821
rect 7656 13744 7708 13796
rect 10600 13855 10652 13864
rect 10600 13821 10609 13855
rect 10609 13821 10643 13855
rect 10643 13821 10652 13855
rect 10600 13812 10652 13821
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 10876 13880 10928 13889
rect 14188 13880 14240 13932
rect 16580 13880 16632 13932
rect 18144 14016 18196 14068
rect 18604 14016 18656 14068
rect 19432 14059 19484 14068
rect 19432 14025 19441 14059
rect 19441 14025 19475 14059
rect 19475 14025 19484 14059
rect 19432 14016 19484 14025
rect 20812 14016 20864 14068
rect 18052 13880 18104 13932
rect 11060 13812 11112 13864
rect 11152 13812 11204 13864
rect 11244 13855 11296 13864
rect 11244 13821 11253 13855
rect 11253 13821 11287 13855
rect 11287 13821 11296 13855
rect 11244 13812 11296 13821
rect 13544 13812 13596 13864
rect 14280 13855 14332 13864
rect 14280 13821 14322 13855
rect 14322 13821 14332 13855
rect 14280 13812 14332 13821
rect 14924 13812 14976 13864
rect 15660 13812 15712 13864
rect 20076 13855 20128 13864
rect 20076 13821 20085 13855
rect 20085 13821 20119 13855
rect 20119 13821 20128 13855
rect 20076 13812 20128 13821
rect 20904 13880 20956 13932
rect 22284 13880 22336 13932
rect 22652 13923 22704 13932
rect 22652 13889 22661 13923
rect 22661 13889 22695 13923
rect 22695 13889 22704 13923
rect 22652 13880 22704 13889
rect 20812 13812 20864 13864
rect 22100 13812 22152 13864
rect 10416 13744 10468 13796
rect 9772 13719 9824 13728
rect 9772 13685 9781 13719
rect 9781 13685 9815 13719
rect 9815 13685 9824 13719
rect 9772 13676 9824 13685
rect 11796 13744 11848 13796
rect 11888 13787 11940 13796
rect 11888 13753 11897 13787
rect 11897 13753 11931 13787
rect 11931 13753 11940 13787
rect 11888 13744 11940 13753
rect 12624 13744 12676 13796
rect 14096 13744 14148 13796
rect 11428 13676 11480 13728
rect 11980 13676 12032 13728
rect 13912 13676 13964 13728
rect 14280 13676 14332 13728
rect 15016 13744 15068 13796
rect 17960 13744 18012 13796
rect 18696 13744 18748 13796
rect 25780 14016 25832 14068
rect 26608 14016 26660 14068
rect 27160 14016 27212 14068
rect 27712 14016 27764 14068
rect 29276 14016 29328 14068
rect 29368 14016 29420 14068
rect 29552 14016 29604 14068
rect 30196 14016 30248 14068
rect 30748 14016 30800 14068
rect 31024 14059 31076 14068
rect 31024 14025 31033 14059
rect 31033 14025 31067 14059
rect 31067 14025 31076 14059
rect 31024 14016 31076 14025
rect 27528 13948 27580 14000
rect 23480 13812 23532 13864
rect 25872 13855 25924 13864
rect 25872 13821 25881 13855
rect 25881 13821 25915 13855
rect 25915 13821 25924 13855
rect 25872 13812 25924 13821
rect 26148 13812 26200 13864
rect 27344 13812 27396 13864
rect 27804 13923 27856 13932
rect 27804 13889 27813 13923
rect 27813 13889 27847 13923
rect 27847 13889 27856 13923
rect 27804 13880 27856 13889
rect 28816 13948 28868 14000
rect 27896 13812 27948 13864
rect 24124 13787 24176 13796
rect 24124 13753 24133 13787
rect 24133 13753 24167 13787
rect 24167 13753 24176 13787
rect 24124 13744 24176 13753
rect 24860 13787 24912 13796
rect 24860 13753 24869 13787
rect 24869 13753 24903 13787
rect 24903 13753 24912 13787
rect 24860 13744 24912 13753
rect 26976 13744 27028 13796
rect 28632 13812 28684 13864
rect 28724 13855 28776 13864
rect 28724 13821 28733 13855
rect 28733 13821 28767 13855
rect 28767 13821 28776 13855
rect 28724 13812 28776 13821
rect 16672 13676 16724 13728
rect 17684 13676 17736 13728
rect 19524 13719 19576 13728
rect 19524 13685 19533 13719
rect 19533 13685 19567 13719
rect 19567 13685 19576 13719
rect 19524 13676 19576 13685
rect 20904 13719 20956 13728
rect 20904 13685 20913 13719
rect 20913 13685 20947 13719
rect 20947 13685 20956 13719
rect 20904 13676 20956 13685
rect 21548 13676 21600 13728
rect 23388 13676 23440 13728
rect 27988 13676 28040 13728
rect 29000 13855 29052 13864
rect 29000 13821 29009 13855
rect 29009 13821 29043 13855
rect 29043 13821 29052 13855
rect 29000 13812 29052 13821
rect 30840 13744 30892 13796
rect 31760 13855 31812 13864
rect 31760 13821 31769 13855
rect 31769 13821 31803 13855
rect 31803 13821 31812 13855
rect 31760 13812 31812 13821
rect 31576 13744 31628 13796
rect 30288 13676 30340 13728
rect 6946 13574 6998 13626
rect 7010 13574 7062 13626
rect 7074 13574 7126 13626
rect 7138 13574 7190 13626
rect 7202 13574 7254 13626
rect 14306 13574 14358 13626
rect 14370 13574 14422 13626
rect 14434 13574 14486 13626
rect 14498 13574 14550 13626
rect 14562 13574 14614 13626
rect 21666 13574 21718 13626
rect 21730 13574 21782 13626
rect 21794 13574 21846 13626
rect 21858 13574 21910 13626
rect 21922 13574 21974 13626
rect 29026 13574 29078 13626
rect 29090 13574 29142 13626
rect 29154 13574 29206 13626
rect 29218 13574 29270 13626
rect 29282 13574 29334 13626
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 10416 13515 10468 13524
rect 10416 13481 10425 13515
rect 10425 13481 10459 13515
rect 10459 13481 10468 13515
rect 10416 13472 10468 13481
rect 9772 13404 9824 13456
rect 6000 13336 6052 13388
rect 1308 13268 1360 13320
rect 10048 13379 10100 13388
rect 10048 13345 10057 13379
rect 10057 13345 10091 13379
rect 10091 13345 10100 13379
rect 10048 13336 10100 13345
rect 11152 13404 11204 13456
rect 11336 13404 11388 13456
rect 12624 13404 12676 13456
rect 12900 13379 12952 13388
rect 12900 13345 12909 13379
rect 12909 13345 12943 13379
rect 12943 13345 12952 13379
rect 12900 13336 12952 13345
rect 13912 13472 13964 13524
rect 14188 13447 14240 13456
rect 14188 13413 14197 13447
rect 14197 13413 14231 13447
rect 14231 13413 14240 13447
rect 14188 13404 14240 13413
rect 14096 13336 14148 13388
rect 15108 13472 15160 13524
rect 15936 13472 15988 13524
rect 16580 13472 16632 13524
rect 16856 13472 16908 13524
rect 17960 13472 18012 13524
rect 18512 13472 18564 13524
rect 18880 13472 18932 13524
rect 19524 13472 19576 13524
rect 14924 13404 14976 13456
rect 20904 13472 20956 13524
rect 22100 13472 22152 13524
rect 24032 13472 24084 13524
rect 24768 13515 24820 13524
rect 24768 13481 24777 13515
rect 24777 13481 24811 13515
rect 24811 13481 24820 13515
rect 24768 13472 24820 13481
rect 24860 13472 24912 13524
rect 25872 13472 25924 13524
rect 14556 13336 14608 13388
rect 14740 13379 14792 13388
rect 14740 13345 14749 13379
rect 14749 13345 14783 13379
rect 14783 13345 14792 13379
rect 14740 13336 14792 13345
rect 16028 13379 16080 13388
rect 16028 13345 16037 13379
rect 16037 13345 16071 13379
rect 16071 13345 16080 13379
rect 16028 13336 16080 13345
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 21456 13404 21508 13456
rect 22652 13404 22704 13456
rect 24124 13404 24176 13456
rect 16856 13379 16908 13388
rect 16856 13345 16865 13379
rect 16865 13345 16899 13379
rect 16899 13345 16908 13379
rect 16856 13336 16908 13345
rect 8024 13268 8076 13320
rect 9772 13311 9824 13320
rect 9772 13277 9781 13311
rect 9781 13277 9815 13311
rect 9815 13277 9824 13311
rect 9772 13268 9824 13277
rect 10968 13268 11020 13320
rect 12532 13268 12584 13320
rect 17408 13336 17460 13388
rect 17224 13311 17276 13320
rect 17224 13277 17233 13311
rect 17233 13277 17267 13311
rect 17267 13277 17276 13311
rect 17224 13268 17276 13277
rect 7288 13200 7340 13252
rect 8300 13175 8352 13184
rect 8300 13141 8309 13175
rect 8309 13141 8343 13175
rect 8343 13141 8352 13175
rect 8300 13132 8352 13141
rect 14004 13200 14056 13252
rect 14740 13200 14792 13252
rect 15752 13132 15804 13184
rect 16580 13200 16632 13252
rect 18972 13336 19024 13388
rect 18696 13268 18748 13320
rect 23480 13336 23532 13388
rect 25596 13379 25648 13388
rect 25596 13345 25605 13379
rect 25605 13345 25639 13379
rect 25639 13345 25648 13379
rect 26976 13404 27028 13456
rect 25596 13336 25648 13345
rect 21364 13268 21416 13320
rect 21824 13311 21876 13320
rect 21824 13277 21833 13311
rect 21833 13277 21867 13311
rect 21867 13277 21876 13311
rect 21824 13268 21876 13277
rect 26424 13311 26476 13320
rect 26424 13277 26433 13311
rect 26433 13277 26467 13311
rect 26467 13277 26476 13311
rect 26424 13268 26476 13277
rect 26700 13268 26752 13320
rect 27620 13268 27672 13320
rect 28632 13404 28684 13456
rect 29368 13404 29420 13456
rect 30564 13404 30616 13456
rect 29000 13379 29052 13388
rect 29000 13345 29009 13379
rect 29009 13345 29043 13379
rect 29043 13345 29052 13379
rect 29000 13336 29052 13345
rect 30932 13472 30984 13524
rect 31760 13472 31812 13524
rect 31024 13404 31076 13456
rect 31668 13379 31720 13388
rect 31668 13345 31677 13379
rect 31677 13345 31711 13379
rect 31711 13345 31720 13379
rect 31668 13336 31720 13345
rect 30840 13268 30892 13320
rect 30932 13311 30984 13320
rect 30932 13277 30941 13311
rect 30941 13277 30975 13311
rect 30975 13277 30984 13311
rect 30932 13268 30984 13277
rect 31760 13311 31812 13320
rect 31760 13277 31769 13311
rect 31769 13277 31803 13311
rect 31803 13277 31812 13311
rect 31760 13268 31812 13277
rect 18604 13175 18656 13184
rect 18604 13141 18613 13175
rect 18613 13141 18647 13175
rect 18647 13141 18656 13175
rect 18604 13132 18656 13141
rect 27988 13200 28040 13252
rect 19524 13132 19576 13184
rect 26792 13175 26844 13184
rect 26792 13141 26801 13175
rect 26801 13141 26835 13175
rect 26835 13141 26844 13175
rect 26792 13132 26844 13141
rect 29000 13200 29052 13252
rect 28448 13175 28500 13184
rect 28448 13141 28457 13175
rect 28457 13141 28491 13175
rect 28491 13141 28500 13175
rect 28448 13132 28500 13141
rect 28724 13132 28776 13184
rect 29828 13132 29880 13184
rect 31760 13132 31812 13184
rect 6286 13030 6338 13082
rect 6350 13030 6402 13082
rect 6414 13030 6466 13082
rect 6478 13030 6530 13082
rect 6542 13030 6594 13082
rect 13646 13030 13698 13082
rect 13710 13030 13762 13082
rect 13774 13030 13826 13082
rect 13838 13030 13890 13082
rect 13902 13030 13954 13082
rect 21006 13030 21058 13082
rect 21070 13030 21122 13082
rect 21134 13030 21186 13082
rect 21198 13030 21250 13082
rect 21262 13030 21314 13082
rect 28366 13030 28418 13082
rect 28430 13030 28482 13082
rect 28494 13030 28546 13082
rect 28558 13030 28610 13082
rect 28622 13030 28674 13082
rect 6644 12971 6696 12980
rect 6644 12937 6653 12971
rect 6653 12937 6687 12971
rect 6687 12937 6696 12971
rect 6644 12928 6696 12937
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 8300 12928 8352 12980
rect 5724 12724 5776 12776
rect 8760 12724 8812 12776
rect 10416 12928 10468 12980
rect 11612 12928 11664 12980
rect 11888 12928 11940 12980
rect 13176 12928 13228 12980
rect 14556 12928 14608 12980
rect 16856 12928 16908 12980
rect 17040 12928 17092 12980
rect 17316 12928 17368 12980
rect 17684 12971 17736 12980
rect 17684 12937 17693 12971
rect 17693 12937 17727 12971
rect 17727 12937 17736 12971
rect 17684 12928 17736 12937
rect 18144 12928 18196 12980
rect 20812 12928 20864 12980
rect 12348 12860 12400 12912
rect 13544 12860 13596 12912
rect 17132 12860 17184 12912
rect 17500 12860 17552 12912
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 12072 12792 12124 12844
rect 12992 12835 13044 12844
rect 12992 12801 13001 12835
rect 13001 12801 13035 12835
rect 13035 12801 13044 12835
rect 12992 12792 13044 12801
rect 14188 12792 14240 12844
rect 15016 12835 15068 12844
rect 15016 12801 15025 12835
rect 15025 12801 15059 12835
rect 15059 12801 15068 12835
rect 15016 12792 15068 12801
rect 10784 12724 10836 12776
rect 11612 12724 11664 12776
rect 8024 12656 8076 12708
rect 8484 12656 8536 12708
rect 12164 12699 12216 12708
rect 12164 12665 12173 12699
rect 12173 12665 12207 12699
rect 12207 12665 12216 12699
rect 12164 12656 12216 12665
rect 13176 12656 13228 12708
rect 14004 12656 14056 12708
rect 14648 12656 14700 12708
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 6920 12588 6972 12640
rect 7932 12588 7984 12640
rect 8576 12588 8628 12640
rect 11152 12588 11204 12640
rect 11704 12588 11756 12640
rect 16948 12792 17000 12844
rect 16672 12724 16724 12776
rect 17040 12767 17092 12776
rect 17040 12733 17049 12767
rect 17049 12733 17083 12767
rect 17083 12733 17092 12767
rect 17040 12724 17092 12733
rect 18604 12792 18656 12844
rect 17960 12724 18012 12776
rect 21548 12928 21600 12980
rect 21824 12971 21876 12980
rect 21824 12937 21833 12971
rect 21833 12937 21867 12971
rect 21867 12937 21876 12971
rect 21824 12928 21876 12937
rect 25596 12928 25648 12980
rect 26792 12928 26844 12980
rect 26884 12928 26936 12980
rect 29460 12928 29512 12980
rect 30656 12928 30708 12980
rect 21364 12860 21416 12912
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 16856 12631 16908 12640
rect 16856 12597 16865 12631
rect 16865 12597 16899 12631
rect 16899 12597 16908 12631
rect 16856 12588 16908 12597
rect 18052 12656 18104 12708
rect 18236 12656 18288 12708
rect 18420 12656 18472 12708
rect 20168 12656 20220 12708
rect 22008 12792 22060 12844
rect 26056 12835 26108 12844
rect 26056 12801 26065 12835
rect 26065 12801 26099 12835
rect 26099 12801 26108 12835
rect 26056 12792 26108 12801
rect 26332 12792 26384 12844
rect 27804 12792 27856 12844
rect 28172 12835 28224 12844
rect 28172 12801 28181 12835
rect 28181 12801 28215 12835
rect 28215 12801 28224 12835
rect 28172 12792 28224 12801
rect 29092 12835 29144 12844
rect 29092 12801 29101 12835
rect 29101 12801 29135 12835
rect 29135 12801 29144 12835
rect 29092 12792 29144 12801
rect 30104 12792 30156 12844
rect 22376 12767 22428 12776
rect 22376 12733 22385 12767
rect 22385 12733 22419 12767
rect 22419 12733 22428 12767
rect 22376 12724 22428 12733
rect 23940 12724 23992 12776
rect 25780 12724 25832 12776
rect 22836 12699 22888 12708
rect 22836 12665 22845 12699
rect 22845 12665 22879 12699
rect 22879 12665 22888 12699
rect 22836 12656 22888 12665
rect 20076 12588 20128 12640
rect 26240 12656 26292 12708
rect 27620 12656 27672 12708
rect 27804 12631 27856 12640
rect 27804 12597 27813 12631
rect 27813 12597 27847 12631
rect 27847 12597 27856 12631
rect 27804 12588 27856 12597
rect 28080 12656 28132 12708
rect 28356 12767 28408 12776
rect 28356 12733 28365 12767
rect 28365 12733 28399 12767
rect 28399 12733 28408 12767
rect 28356 12724 28408 12733
rect 28172 12588 28224 12640
rect 28632 12588 28684 12640
rect 28816 12699 28868 12708
rect 28816 12665 28825 12699
rect 28825 12665 28859 12699
rect 28859 12665 28868 12699
rect 28816 12656 28868 12665
rect 29276 12656 29328 12708
rect 29644 12656 29696 12708
rect 29828 12656 29880 12708
rect 30656 12588 30708 12640
rect 6946 12486 6998 12538
rect 7010 12486 7062 12538
rect 7074 12486 7126 12538
rect 7138 12486 7190 12538
rect 7202 12486 7254 12538
rect 14306 12486 14358 12538
rect 14370 12486 14422 12538
rect 14434 12486 14486 12538
rect 14498 12486 14550 12538
rect 14562 12486 14614 12538
rect 21666 12486 21718 12538
rect 21730 12486 21782 12538
rect 21794 12486 21846 12538
rect 21858 12486 21910 12538
rect 21922 12486 21974 12538
rect 29026 12486 29078 12538
rect 29090 12486 29142 12538
rect 29154 12486 29206 12538
rect 29218 12486 29270 12538
rect 29282 12486 29334 12538
rect 5724 12427 5776 12436
rect 5724 12393 5733 12427
rect 5733 12393 5767 12427
rect 5767 12393 5776 12427
rect 5724 12384 5776 12393
rect 7932 12384 7984 12436
rect 8116 12384 8168 12436
rect 8576 12384 8628 12436
rect 4344 12316 4396 12368
rect 5632 12316 5684 12368
rect 6920 12359 6972 12368
rect 6920 12325 6929 12359
rect 6929 12325 6963 12359
rect 6963 12325 6972 12359
rect 6920 12316 6972 12325
rect 7840 12316 7892 12368
rect 8760 12316 8812 12368
rect 9772 12384 9824 12436
rect 11612 12384 11664 12436
rect 12440 12384 12492 12436
rect 11152 12359 11204 12368
rect 11152 12325 11161 12359
rect 11161 12325 11195 12359
rect 11195 12325 11204 12359
rect 11152 12316 11204 12325
rect 11704 12316 11756 12368
rect 12256 12359 12308 12368
rect 12256 12325 12265 12359
rect 12265 12325 12299 12359
rect 12299 12325 12308 12359
rect 12256 12316 12308 12325
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 14096 12359 14148 12368
rect 14096 12325 14105 12359
rect 14105 12325 14139 12359
rect 14139 12325 14148 12359
rect 14096 12316 14148 12325
rect 14648 12316 14700 12368
rect 15384 12316 15436 12368
rect 15752 12316 15804 12368
rect 18420 12384 18472 12436
rect 18972 12384 19024 12436
rect 20168 12427 20220 12436
rect 20168 12393 20177 12427
rect 20177 12393 20211 12427
rect 20211 12393 20220 12427
rect 20168 12384 20220 12393
rect 20628 12384 20680 12436
rect 22376 12384 22428 12436
rect 22652 12427 22704 12436
rect 22652 12393 22661 12427
rect 22661 12393 22695 12427
rect 22695 12393 22704 12427
rect 22652 12384 22704 12393
rect 22744 12384 22796 12436
rect 22928 12427 22980 12436
rect 22928 12393 22937 12427
rect 22937 12393 22971 12427
rect 22971 12393 22980 12427
rect 22928 12384 22980 12393
rect 5724 12248 5776 12300
rect 5632 12223 5684 12232
rect 5632 12189 5641 12223
rect 5641 12189 5675 12223
rect 5675 12189 5684 12223
rect 5632 12180 5684 12189
rect 6644 12180 6696 12232
rect 6828 12291 6880 12300
rect 6828 12257 6837 12291
rect 6837 12257 6871 12291
rect 6871 12257 6880 12291
rect 6828 12248 6880 12257
rect 7104 12291 7156 12300
rect 7104 12257 7113 12291
rect 7113 12257 7147 12291
rect 7147 12257 7156 12291
rect 7104 12248 7156 12257
rect 7380 12248 7432 12300
rect 7932 12248 7984 12300
rect 8024 12291 8076 12300
rect 8024 12257 8033 12291
rect 8033 12257 8067 12291
rect 8067 12257 8076 12291
rect 8024 12248 8076 12257
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 4712 12044 4764 12096
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10876 12248 10928 12300
rect 16856 12291 16908 12300
rect 16856 12257 16865 12291
rect 16865 12257 16899 12291
rect 16899 12257 16908 12291
rect 16856 12248 16908 12257
rect 18604 12248 18656 12300
rect 19248 12248 19300 12300
rect 21456 12316 21508 12368
rect 22100 12316 22152 12368
rect 22284 12316 22336 12368
rect 23756 12384 23808 12436
rect 23940 12384 23992 12436
rect 24124 12384 24176 12436
rect 24860 12427 24912 12436
rect 24860 12393 24869 12427
rect 24869 12393 24903 12427
rect 24903 12393 24912 12427
rect 24860 12384 24912 12393
rect 25688 12384 25740 12436
rect 26700 12384 26752 12436
rect 23480 12316 23532 12368
rect 10048 12180 10100 12189
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 12624 12180 12676 12232
rect 13084 12180 13136 12232
rect 9680 12112 9732 12164
rect 15292 12180 15344 12232
rect 16304 12223 16356 12232
rect 16304 12189 16313 12223
rect 16313 12189 16347 12223
rect 16347 12189 16356 12223
rect 16304 12180 16356 12189
rect 16948 12180 17000 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 8852 12044 8904 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 16672 12087 16724 12096
rect 16672 12053 16681 12087
rect 16681 12053 16715 12087
rect 16715 12053 16724 12087
rect 16672 12044 16724 12053
rect 16856 12044 16908 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 18144 12087 18196 12096
rect 18144 12053 18153 12087
rect 18153 12053 18187 12087
rect 18187 12053 18196 12087
rect 18144 12044 18196 12053
rect 19064 12044 19116 12096
rect 19984 12087 20036 12096
rect 19984 12053 19993 12087
rect 19993 12053 20027 12087
rect 20027 12053 20036 12087
rect 19984 12044 20036 12053
rect 22836 12291 22888 12300
rect 22836 12257 22845 12291
rect 22845 12257 22879 12291
rect 22879 12257 22888 12291
rect 22836 12248 22888 12257
rect 23388 12248 23440 12300
rect 26332 12359 26384 12368
rect 26332 12325 26341 12359
rect 26341 12325 26375 12359
rect 26375 12325 26384 12359
rect 26332 12316 26384 12325
rect 26608 12316 26660 12368
rect 26884 12316 26936 12368
rect 23756 12180 23808 12232
rect 24952 12248 25004 12300
rect 25688 12291 25740 12300
rect 25688 12257 25697 12291
rect 25697 12257 25731 12291
rect 25731 12257 25740 12291
rect 25688 12248 25740 12257
rect 26976 12248 27028 12300
rect 28632 12384 28684 12436
rect 29736 12384 29788 12436
rect 28356 12316 28408 12368
rect 28724 12316 28776 12368
rect 27804 12291 27856 12300
rect 27804 12257 27813 12291
rect 27813 12257 27847 12291
rect 27847 12257 27856 12291
rect 27804 12248 27856 12257
rect 29184 12291 29236 12300
rect 29184 12257 29193 12291
rect 29193 12257 29227 12291
rect 29227 12257 29236 12291
rect 29184 12248 29236 12257
rect 29552 12316 29604 12368
rect 27436 12180 27488 12232
rect 30104 12316 30156 12368
rect 29736 12248 29788 12300
rect 30196 12291 30248 12300
rect 30196 12257 30205 12291
rect 30205 12257 30239 12291
rect 30239 12257 30248 12291
rect 30196 12248 30248 12257
rect 26148 12112 26200 12164
rect 26240 12112 26292 12164
rect 33140 12248 33192 12300
rect 22836 12044 22888 12096
rect 23480 12087 23532 12096
rect 23480 12053 23489 12087
rect 23489 12053 23523 12087
rect 23523 12053 23532 12087
rect 23480 12044 23532 12053
rect 25136 12044 25188 12096
rect 25872 12044 25924 12096
rect 26608 12044 26660 12096
rect 28816 12044 28868 12096
rect 29184 12044 29236 12096
rect 29828 12044 29880 12096
rect 6286 11942 6338 11994
rect 6350 11942 6402 11994
rect 6414 11942 6466 11994
rect 6478 11942 6530 11994
rect 6542 11942 6594 11994
rect 13646 11942 13698 11994
rect 13710 11942 13762 11994
rect 13774 11942 13826 11994
rect 13838 11942 13890 11994
rect 13902 11942 13954 11994
rect 21006 11942 21058 11994
rect 21070 11942 21122 11994
rect 21134 11942 21186 11994
rect 21198 11942 21250 11994
rect 21262 11942 21314 11994
rect 28366 11942 28418 11994
rect 28430 11942 28482 11994
rect 28494 11942 28546 11994
rect 28558 11942 28610 11994
rect 28622 11942 28674 11994
rect 4344 11840 4396 11892
rect 4712 11840 4764 11892
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 6828 11840 6880 11892
rect 7840 11840 7892 11892
rect 8024 11840 8076 11892
rect 8484 11747 8536 11756
rect 8484 11713 8493 11747
rect 8493 11713 8527 11747
rect 8527 11713 8536 11747
rect 8484 11704 8536 11713
rect 8668 11704 8720 11756
rect 6092 11636 6144 11688
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 9496 11636 9548 11688
rect 9772 11840 9824 11892
rect 10600 11840 10652 11892
rect 14096 11840 14148 11892
rect 19708 11840 19760 11892
rect 11060 11704 11112 11756
rect 15384 11815 15436 11824
rect 15384 11781 15393 11815
rect 15393 11781 15427 11815
rect 15427 11781 15436 11815
rect 15384 11772 15436 11781
rect 16948 11815 17000 11824
rect 16948 11781 16957 11815
rect 16957 11781 16991 11815
rect 16991 11781 17000 11815
rect 16948 11772 17000 11781
rect 17224 11772 17276 11824
rect 17408 11772 17460 11824
rect 19432 11772 19484 11824
rect 10508 11636 10560 11688
rect 4436 11500 4488 11552
rect 5264 11543 5316 11552
rect 5264 11509 5273 11543
rect 5273 11509 5307 11543
rect 5307 11509 5316 11543
rect 5264 11500 5316 11509
rect 5540 11543 5592 11552
rect 5540 11509 5549 11543
rect 5549 11509 5583 11543
rect 5583 11509 5592 11543
rect 5540 11500 5592 11509
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 7748 11568 7800 11620
rect 8576 11568 8628 11620
rect 11704 11611 11756 11620
rect 11704 11577 11713 11611
rect 11713 11577 11747 11611
rect 11747 11577 11756 11611
rect 11704 11568 11756 11577
rect 12072 11636 12124 11688
rect 12900 11704 12952 11756
rect 12256 11679 12308 11688
rect 12256 11645 12265 11679
rect 12265 11645 12299 11679
rect 12299 11645 12308 11679
rect 12256 11636 12308 11645
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 14004 11636 14056 11688
rect 14924 11704 14976 11756
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 19064 11747 19116 11756
rect 19064 11713 19073 11747
rect 19073 11713 19107 11747
rect 19107 11713 19116 11747
rect 19064 11704 19116 11713
rect 8392 11500 8444 11552
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 10600 11543 10652 11552
rect 10600 11509 10609 11543
rect 10609 11509 10643 11543
rect 10643 11509 10652 11543
rect 10600 11500 10652 11509
rect 12072 11543 12124 11552
rect 12072 11509 12081 11543
rect 12081 11509 12115 11543
rect 12115 11509 12124 11543
rect 12072 11500 12124 11509
rect 12348 11500 12400 11552
rect 12992 11543 13044 11552
rect 12992 11509 13001 11543
rect 13001 11509 13035 11543
rect 13035 11509 13044 11543
rect 12992 11500 13044 11509
rect 15476 11500 15528 11552
rect 15844 11636 15896 11688
rect 18696 11679 18748 11688
rect 18696 11645 18705 11679
rect 18705 11645 18739 11679
rect 18739 11645 18748 11679
rect 18696 11636 18748 11645
rect 20168 11636 20220 11688
rect 17960 11568 18012 11620
rect 18420 11568 18472 11620
rect 20536 11636 20588 11688
rect 23480 11840 23532 11892
rect 26608 11840 26660 11892
rect 27436 11840 27488 11892
rect 29736 11840 29788 11892
rect 30932 11840 30984 11892
rect 24216 11772 24268 11824
rect 24492 11815 24544 11824
rect 24492 11781 24501 11815
rect 24501 11781 24535 11815
rect 24535 11781 24544 11815
rect 24492 11772 24544 11781
rect 24952 11772 25004 11824
rect 27252 11772 27304 11824
rect 21364 11704 21416 11756
rect 30288 11772 30340 11824
rect 30840 11815 30892 11824
rect 30840 11781 30849 11815
rect 30849 11781 30883 11815
rect 30883 11781 30892 11815
rect 30840 11772 30892 11781
rect 20720 11636 20772 11688
rect 24584 11636 24636 11688
rect 24860 11636 24912 11688
rect 24952 11679 25004 11688
rect 24952 11645 24961 11679
rect 24961 11645 24995 11679
rect 24995 11645 25004 11679
rect 24952 11636 25004 11645
rect 25136 11679 25188 11688
rect 25136 11645 25145 11679
rect 25145 11645 25179 11679
rect 25179 11645 25188 11679
rect 25136 11636 25188 11645
rect 25413 11679 25465 11688
rect 25413 11645 25421 11679
rect 25421 11645 25455 11679
rect 25455 11645 25465 11679
rect 25413 11636 25465 11645
rect 25872 11679 25924 11688
rect 25872 11645 25881 11679
rect 25881 11645 25915 11679
rect 25915 11645 25924 11679
rect 25872 11636 25924 11645
rect 26976 11679 27028 11688
rect 26976 11645 26982 11679
rect 26982 11645 27016 11679
rect 27016 11645 27028 11679
rect 26976 11636 27028 11645
rect 25504 11611 25556 11620
rect 25504 11577 25513 11611
rect 25513 11577 25547 11611
rect 25547 11577 25556 11611
rect 25504 11568 25556 11577
rect 25596 11611 25648 11620
rect 25596 11577 25605 11611
rect 25605 11577 25639 11611
rect 25639 11577 25648 11611
rect 25596 11568 25648 11577
rect 26148 11568 26200 11620
rect 26424 11568 26476 11620
rect 26884 11568 26936 11620
rect 27436 11636 27488 11688
rect 27712 11636 27764 11688
rect 27804 11636 27856 11688
rect 27988 11636 28040 11688
rect 29368 11704 29420 11756
rect 29460 11704 29512 11756
rect 31760 11747 31812 11756
rect 31760 11713 31769 11747
rect 31769 11713 31803 11747
rect 31803 11713 31812 11747
rect 31760 11704 31812 11713
rect 28172 11679 28224 11688
rect 28172 11645 28181 11679
rect 28181 11645 28215 11679
rect 28215 11645 28224 11679
rect 28172 11636 28224 11645
rect 16212 11500 16264 11552
rect 16764 11543 16816 11552
rect 16764 11509 16773 11543
rect 16773 11509 16807 11543
rect 16807 11509 16816 11543
rect 16764 11500 16816 11509
rect 18788 11500 18840 11552
rect 25136 11543 25188 11552
rect 25136 11509 25145 11543
rect 25145 11509 25179 11543
rect 25179 11509 25188 11543
rect 25136 11500 25188 11509
rect 25228 11543 25280 11552
rect 25228 11509 25237 11543
rect 25237 11509 25271 11543
rect 25271 11509 25280 11543
rect 25228 11500 25280 11509
rect 26332 11500 26384 11552
rect 27804 11543 27856 11552
rect 27804 11509 27813 11543
rect 27813 11509 27847 11543
rect 27847 11509 27856 11543
rect 27804 11500 27856 11509
rect 28080 11500 28132 11552
rect 30472 11611 30524 11620
rect 30472 11577 30481 11611
rect 30481 11577 30515 11611
rect 30515 11577 30524 11611
rect 30472 11568 30524 11577
rect 28908 11500 28960 11552
rect 30196 11500 30248 11552
rect 30380 11543 30432 11552
rect 30380 11509 30389 11543
rect 30389 11509 30423 11543
rect 30423 11509 30432 11543
rect 30380 11500 30432 11509
rect 6946 11398 6998 11450
rect 7010 11398 7062 11450
rect 7074 11398 7126 11450
rect 7138 11398 7190 11450
rect 7202 11398 7254 11450
rect 14306 11398 14358 11450
rect 14370 11398 14422 11450
rect 14434 11398 14486 11450
rect 14498 11398 14550 11450
rect 14562 11398 14614 11450
rect 21666 11398 21718 11450
rect 21730 11398 21782 11450
rect 21794 11398 21846 11450
rect 21858 11398 21910 11450
rect 21922 11398 21974 11450
rect 29026 11398 29078 11450
rect 29090 11398 29142 11450
rect 29154 11398 29206 11450
rect 29218 11398 29270 11450
rect 29282 11398 29334 11450
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 5632 11296 5684 11348
rect 6092 11296 6144 11348
rect 6644 11296 6696 11348
rect 7748 11339 7800 11348
rect 7748 11305 7757 11339
rect 7757 11305 7791 11339
rect 7791 11305 7800 11339
rect 7748 11296 7800 11305
rect 7840 11296 7892 11348
rect 8392 11339 8444 11348
rect 8392 11305 8401 11339
rect 8401 11305 8435 11339
rect 8435 11305 8444 11339
rect 8392 11296 8444 11305
rect 9128 11296 9180 11348
rect 12256 11296 12308 11348
rect 12348 11339 12400 11348
rect 12348 11305 12357 11339
rect 12357 11305 12391 11339
rect 12391 11305 12400 11339
rect 12348 11296 12400 11305
rect 13544 11296 13596 11348
rect 17960 11339 18012 11348
rect 17960 11305 17969 11339
rect 17969 11305 18003 11339
rect 18003 11305 18012 11339
rect 17960 11296 18012 11305
rect 5264 11271 5316 11280
rect 5264 11237 5273 11271
rect 5273 11237 5307 11271
rect 5307 11237 5316 11271
rect 5264 11228 5316 11237
rect 5816 11228 5868 11280
rect 6736 11160 6788 11212
rect 8668 11228 8720 11280
rect 3240 11135 3292 11144
rect 3240 11101 3249 11135
rect 3249 11101 3283 11135
rect 3283 11101 3292 11135
rect 3240 11092 3292 11101
rect 8852 11092 8904 11144
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 9128 11160 9180 11169
rect 9312 11160 9364 11212
rect 9680 11160 9732 11212
rect 9864 11203 9916 11212
rect 9864 11169 9873 11203
rect 9873 11169 9907 11203
rect 9907 11169 9916 11203
rect 9864 11160 9916 11169
rect 10416 11228 10468 11280
rect 10600 11228 10652 11280
rect 12072 11228 12124 11280
rect 8024 10999 8076 11008
rect 8024 10965 8033 10999
rect 8033 10965 8067 10999
rect 8067 10965 8076 10999
rect 8024 10956 8076 10965
rect 9496 11135 9548 11144
rect 9496 11101 9505 11135
rect 9505 11101 9539 11135
rect 9539 11101 9548 11135
rect 9496 11092 9548 11101
rect 9588 11135 9640 11144
rect 9588 11101 9597 11135
rect 9597 11101 9631 11135
rect 9631 11101 9640 11135
rect 9588 11092 9640 11101
rect 10048 11092 10100 11144
rect 10508 11092 10560 11144
rect 18972 11296 19024 11348
rect 22560 11296 22612 11348
rect 18880 11228 18932 11280
rect 19984 11228 20036 11280
rect 26424 11296 26476 11348
rect 28908 11296 28960 11348
rect 12440 11024 12492 11076
rect 10140 10999 10192 11008
rect 10140 10965 10149 10999
rect 10149 10965 10183 10999
rect 10183 10965 10192 10999
rect 10140 10956 10192 10965
rect 11520 10956 11572 11008
rect 14004 11203 14056 11212
rect 14004 11169 14013 11203
rect 14013 11169 14047 11203
rect 14047 11169 14056 11203
rect 14004 11160 14056 11169
rect 15108 11160 15160 11212
rect 12624 11092 12676 11144
rect 13452 11024 13504 11076
rect 14924 11092 14976 11144
rect 16764 11160 16816 11212
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 20168 11203 20220 11212
rect 20168 11169 20177 11203
rect 20177 11169 20211 11203
rect 20211 11169 20220 11203
rect 20168 11160 20220 11169
rect 20260 11160 20312 11212
rect 22100 11203 22152 11212
rect 22100 11169 22109 11203
rect 22109 11169 22143 11203
rect 22143 11169 22152 11203
rect 22100 11160 22152 11169
rect 22376 11160 22428 11212
rect 25136 11228 25188 11280
rect 25412 11228 25464 11280
rect 26884 11228 26936 11280
rect 27160 11228 27212 11280
rect 28632 11228 28684 11280
rect 29368 11296 29420 11348
rect 30380 11296 30432 11348
rect 30748 11339 30800 11348
rect 30748 11305 30757 11339
rect 30757 11305 30791 11339
rect 30791 11305 30800 11339
rect 30748 11296 30800 11305
rect 30840 11296 30892 11348
rect 31300 11296 31352 11348
rect 31576 11339 31628 11348
rect 31576 11305 31585 11339
rect 31585 11305 31619 11339
rect 31619 11305 31628 11339
rect 31576 11296 31628 11305
rect 26240 11160 26292 11212
rect 29736 11160 29788 11212
rect 30104 11203 30156 11212
rect 30104 11169 30113 11203
rect 30113 11169 30147 11203
rect 30147 11169 30156 11203
rect 30104 11160 30156 11169
rect 30288 11203 30340 11212
rect 30288 11169 30297 11203
rect 30297 11169 30331 11203
rect 30331 11169 30340 11203
rect 30288 11160 30340 11169
rect 31392 11203 31444 11212
rect 31392 11169 31401 11203
rect 31401 11169 31435 11203
rect 31435 11169 31444 11203
rect 31392 11160 31444 11169
rect 31668 11203 31720 11212
rect 31668 11169 31677 11203
rect 31677 11169 31711 11203
rect 31711 11169 31720 11203
rect 31668 11160 31720 11169
rect 19248 11092 19300 11144
rect 20812 11092 20864 11144
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 25136 11135 25188 11144
rect 25136 11101 25145 11135
rect 25145 11101 25179 11135
rect 25179 11101 25188 11135
rect 25136 11092 25188 11101
rect 27068 11092 27120 11144
rect 16856 11024 16908 11076
rect 18420 11067 18472 11076
rect 18420 11033 18429 11067
rect 18429 11033 18463 11067
rect 18463 11033 18472 11067
rect 18420 11024 18472 11033
rect 21364 11024 21416 11076
rect 16672 10956 16724 11008
rect 18788 10956 18840 11008
rect 24400 10956 24452 11008
rect 25320 10956 25372 11008
rect 31484 11024 31536 11076
rect 27712 10956 27764 11008
rect 28724 10956 28776 11008
rect 28816 10999 28868 11008
rect 28816 10965 28825 10999
rect 28825 10965 28859 10999
rect 28859 10965 28868 10999
rect 28816 10956 28868 10965
rect 31024 10956 31076 11008
rect 6286 10854 6338 10906
rect 6350 10854 6402 10906
rect 6414 10854 6466 10906
rect 6478 10854 6530 10906
rect 6542 10854 6594 10906
rect 13646 10854 13698 10906
rect 13710 10854 13762 10906
rect 13774 10854 13826 10906
rect 13838 10854 13890 10906
rect 13902 10854 13954 10906
rect 21006 10854 21058 10906
rect 21070 10854 21122 10906
rect 21134 10854 21186 10906
rect 21198 10854 21250 10906
rect 21262 10854 21314 10906
rect 28366 10854 28418 10906
rect 28430 10854 28482 10906
rect 28494 10854 28546 10906
rect 28558 10854 28610 10906
rect 28622 10854 28674 10906
rect 5908 10752 5960 10804
rect 6368 10752 6420 10804
rect 8576 10795 8628 10804
rect 8576 10761 8585 10795
rect 8585 10761 8619 10795
rect 8619 10761 8628 10795
rect 8576 10752 8628 10761
rect 6000 10616 6052 10668
rect 8024 10659 8076 10668
rect 8024 10625 8033 10659
rect 8033 10625 8067 10659
rect 8067 10625 8076 10659
rect 8024 10616 8076 10625
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 10140 10616 10192 10625
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 12992 10752 13044 10804
rect 13176 10752 13228 10804
rect 14004 10752 14056 10804
rect 18880 10752 18932 10804
rect 20260 10752 20312 10804
rect 20720 10795 20772 10804
rect 20720 10761 20729 10795
rect 20729 10761 20763 10795
rect 20763 10761 20772 10795
rect 20720 10752 20772 10761
rect 20904 10752 20956 10804
rect 23756 10795 23808 10804
rect 23756 10761 23765 10795
rect 23765 10761 23799 10795
rect 23799 10761 23808 10795
rect 23756 10752 23808 10761
rect 25136 10752 25188 10804
rect 27068 10752 27120 10804
rect 29460 10752 29512 10804
rect 30104 10752 30156 10804
rect 30196 10752 30248 10804
rect 30288 10795 30340 10804
rect 30288 10761 30297 10795
rect 30297 10761 30331 10795
rect 30331 10761 30340 10795
rect 30288 10752 30340 10761
rect 15660 10684 15712 10736
rect 19340 10684 19392 10736
rect 12532 10616 12584 10668
rect 13452 10616 13504 10668
rect 15016 10616 15068 10668
rect 16304 10659 16356 10668
rect 16304 10625 16313 10659
rect 16313 10625 16347 10659
rect 16347 10625 16356 10659
rect 16304 10616 16356 10625
rect 16672 10616 16724 10668
rect 4344 10548 4396 10600
rect 9680 10480 9732 10532
rect 6276 10455 6328 10464
rect 6276 10421 6285 10455
rect 6285 10421 6319 10455
rect 6319 10421 6328 10455
rect 6276 10412 6328 10421
rect 8668 10455 8720 10464
rect 8668 10421 8677 10455
rect 8677 10421 8711 10455
rect 8711 10421 8720 10455
rect 8668 10412 8720 10421
rect 11520 10412 11572 10464
rect 13084 10591 13136 10600
rect 13084 10557 13093 10591
rect 13093 10557 13127 10591
rect 13127 10557 13136 10591
rect 13084 10548 13136 10557
rect 14648 10548 14700 10600
rect 15200 10591 15252 10600
rect 15200 10557 15209 10591
rect 15209 10557 15243 10591
rect 15243 10557 15252 10591
rect 15200 10548 15252 10557
rect 19248 10616 19300 10668
rect 22928 10684 22980 10736
rect 14096 10480 14148 10532
rect 12716 10412 12768 10464
rect 15568 10480 15620 10532
rect 18420 10480 18472 10532
rect 20720 10480 20772 10532
rect 22284 10591 22336 10600
rect 22284 10557 22293 10591
rect 22293 10557 22327 10591
rect 22327 10557 22336 10591
rect 22284 10548 22336 10557
rect 21456 10523 21508 10532
rect 21456 10489 21465 10523
rect 21465 10489 21499 10523
rect 21499 10489 21508 10523
rect 21456 10480 21508 10489
rect 22008 10480 22060 10532
rect 25228 10616 25280 10668
rect 27160 10616 27212 10668
rect 29368 10616 29420 10668
rect 23204 10548 23256 10600
rect 23664 10480 23716 10532
rect 24124 10548 24176 10600
rect 26424 10548 26476 10600
rect 28724 10548 28776 10600
rect 15292 10412 15344 10464
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 15936 10412 15988 10464
rect 19248 10412 19300 10464
rect 20996 10412 21048 10464
rect 22376 10412 22428 10464
rect 23020 10455 23072 10464
rect 23020 10421 23029 10455
rect 23029 10421 23063 10455
rect 23063 10421 23072 10455
rect 23020 10412 23072 10421
rect 24860 10480 24912 10532
rect 29552 10591 29604 10600
rect 29552 10557 29561 10591
rect 29561 10557 29595 10591
rect 29595 10557 29604 10591
rect 29552 10548 29604 10557
rect 30748 10548 30800 10600
rect 30932 10591 30984 10600
rect 30932 10557 30941 10591
rect 30941 10557 30975 10591
rect 30975 10557 30984 10591
rect 30932 10548 30984 10557
rect 24308 10412 24360 10464
rect 24400 10412 24452 10464
rect 29644 10480 29696 10532
rect 30288 10480 30340 10532
rect 31392 10480 31444 10532
rect 29736 10412 29788 10464
rect 29920 10412 29972 10464
rect 6946 10310 6998 10362
rect 7010 10310 7062 10362
rect 7074 10310 7126 10362
rect 7138 10310 7190 10362
rect 7202 10310 7254 10362
rect 14306 10310 14358 10362
rect 14370 10310 14422 10362
rect 14434 10310 14486 10362
rect 14498 10310 14550 10362
rect 14562 10310 14614 10362
rect 21666 10310 21718 10362
rect 21730 10310 21782 10362
rect 21794 10310 21846 10362
rect 21858 10310 21910 10362
rect 21922 10310 21974 10362
rect 29026 10310 29078 10362
rect 29090 10310 29142 10362
rect 29154 10310 29206 10362
rect 29218 10310 29270 10362
rect 29282 10310 29334 10362
rect 6276 10208 6328 10260
rect 6368 10251 6420 10260
rect 6368 10217 6377 10251
rect 6377 10217 6411 10251
rect 6411 10217 6420 10251
rect 6368 10208 6420 10217
rect 9312 10208 9364 10260
rect 9680 10208 9732 10260
rect 10508 10251 10560 10260
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 12440 10208 12492 10260
rect 14096 10251 14148 10260
rect 14096 10217 14105 10251
rect 14105 10217 14139 10251
rect 14139 10217 14148 10251
rect 14096 10208 14148 10217
rect 5540 10140 5592 10192
rect 9772 10140 9824 10192
rect 3056 10115 3108 10124
rect 3056 10081 3065 10115
rect 3065 10081 3099 10115
rect 3099 10081 3108 10115
rect 3056 10072 3108 10081
rect 12716 10072 12768 10124
rect 14924 10208 14976 10260
rect 15568 10208 15620 10260
rect 17316 10208 17368 10260
rect 18420 10251 18472 10260
rect 18420 10217 18429 10251
rect 18429 10217 18463 10251
rect 18463 10217 18472 10251
rect 18420 10208 18472 10217
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 19340 10208 19392 10260
rect 22284 10208 22336 10260
rect 20996 10140 21048 10192
rect 24124 10140 24176 10192
rect 26240 10208 26292 10260
rect 26424 10251 26476 10260
rect 26424 10217 26433 10251
rect 26433 10217 26467 10251
rect 26467 10217 26476 10251
rect 26424 10208 26476 10217
rect 28080 10208 28132 10260
rect 29552 10208 29604 10260
rect 29920 10208 29972 10260
rect 30932 10208 30984 10260
rect 16764 10072 16816 10124
rect 18788 10072 18840 10124
rect 6092 10047 6144 10056
rect 6092 10013 6101 10047
rect 6101 10013 6135 10047
rect 6135 10013 6144 10047
rect 6092 10004 6144 10013
rect 14648 10047 14700 10056
rect 14648 10013 14657 10047
rect 14657 10013 14691 10047
rect 14691 10013 14700 10047
rect 14648 10004 14700 10013
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 15384 10004 15436 10056
rect 16580 10004 16632 10056
rect 19248 10004 19300 10056
rect 23388 10072 23440 10124
rect 25504 10140 25556 10192
rect 24860 10072 24912 10124
rect 25412 10072 25464 10124
rect 25780 10072 25832 10124
rect 26884 10115 26936 10124
rect 26884 10081 26893 10115
rect 26893 10081 26927 10115
rect 26927 10081 26936 10115
rect 26884 10072 26936 10081
rect 27620 10140 27672 10192
rect 27804 10140 27856 10192
rect 28172 10140 28224 10192
rect 27252 10072 27304 10124
rect 3240 9911 3292 9920
rect 3240 9877 3249 9911
rect 3249 9877 3283 9911
rect 3283 9877 3292 9911
rect 3240 9868 3292 9877
rect 4344 9911 4396 9920
rect 4344 9877 4353 9911
rect 4353 9877 4387 9911
rect 4387 9877 4396 9911
rect 4344 9868 4396 9877
rect 17960 9911 18012 9920
rect 17960 9877 17969 9911
rect 17969 9877 18003 9911
rect 18003 9877 18012 9911
rect 17960 9868 18012 9877
rect 18512 9868 18564 9920
rect 20720 9868 20772 9920
rect 21456 9868 21508 9920
rect 22376 10004 22428 10056
rect 23572 10004 23624 10056
rect 27712 10047 27764 10056
rect 27712 10013 27721 10047
rect 27721 10013 27755 10047
rect 27755 10013 27764 10047
rect 27712 10004 27764 10013
rect 27988 10004 28040 10056
rect 23480 9868 23532 9920
rect 27436 9868 27488 9920
rect 27896 9868 27948 9920
rect 28264 9911 28316 9920
rect 28264 9877 28273 9911
rect 28273 9877 28307 9911
rect 28307 9877 28316 9911
rect 28264 9868 28316 9877
rect 28724 9868 28776 9920
rect 28908 10115 28960 10124
rect 28908 10081 28917 10115
rect 28917 10081 28951 10115
rect 28951 10081 28960 10115
rect 28908 10072 28960 10081
rect 29092 10115 29144 10124
rect 29092 10081 29101 10115
rect 29101 10081 29135 10115
rect 29135 10081 29144 10115
rect 29092 10072 29144 10081
rect 31392 10115 31444 10124
rect 31392 10081 31401 10115
rect 31401 10081 31435 10115
rect 31435 10081 31444 10115
rect 31392 10072 31444 10081
rect 31484 10115 31536 10124
rect 31484 10081 31493 10115
rect 31493 10081 31527 10115
rect 31527 10081 31536 10115
rect 31484 10072 31536 10081
rect 29368 10047 29420 10056
rect 29368 10013 29377 10047
rect 29377 10013 29411 10047
rect 29411 10013 29420 10047
rect 29368 10004 29420 10013
rect 29644 10004 29696 10056
rect 30196 10004 30248 10056
rect 6286 9766 6338 9818
rect 6350 9766 6402 9818
rect 6414 9766 6466 9818
rect 6478 9766 6530 9818
rect 6542 9766 6594 9818
rect 13646 9766 13698 9818
rect 13710 9766 13762 9818
rect 13774 9766 13826 9818
rect 13838 9766 13890 9818
rect 13902 9766 13954 9818
rect 21006 9766 21058 9818
rect 21070 9766 21122 9818
rect 21134 9766 21186 9818
rect 21198 9766 21250 9818
rect 21262 9766 21314 9818
rect 28366 9766 28418 9818
rect 28430 9766 28482 9818
rect 28494 9766 28546 9818
rect 28558 9766 28610 9818
rect 28622 9766 28674 9818
rect 8668 9528 8720 9580
rect 14924 9707 14976 9716
rect 14924 9673 14933 9707
rect 14933 9673 14967 9707
rect 14967 9673 14976 9707
rect 14924 9664 14976 9673
rect 15200 9664 15252 9716
rect 15384 9664 15436 9716
rect 21824 9664 21876 9716
rect 22560 9664 22612 9716
rect 23204 9664 23256 9716
rect 15844 9596 15896 9648
rect 19156 9596 19208 9648
rect 15016 9528 15068 9580
rect 15292 9528 15344 9580
rect 16580 9571 16632 9580
rect 16580 9537 16589 9571
rect 16589 9537 16623 9571
rect 16623 9537 16632 9571
rect 16580 9528 16632 9537
rect 20260 9571 20312 9580
rect 20260 9537 20269 9571
rect 20269 9537 20303 9571
rect 20303 9537 20312 9571
rect 20260 9528 20312 9537
rect 20904 9528 20956 9580
rect 14004 9460 14056 9512
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 18052 9503 18104 9512
rect 18052 9469 18061 9503
rect 18061 9469 18095 9503
rect 18095 9469 18104 9503
rect 18052 9460 18104 9469
rect 20352 9503 20404 9512
rect 20352 9469 20361 9503
rect 20361 9469 20395 9503
rect 20395 9469 20404 9503
rect 20352 9460 20404 9469
rect 20812 9460 20864 9512
rect 18604 9435 18656 9444
rect 18604 9401 18613 9435
rect 18613 9401 18647 9435
rect 18647 9401 18656 9435
rect 18604 9392 18656 9401
rect 8300 9324 8352 9376
rect 9588 9324 9640 9376
rect 13544 9324 13596 9376
rect 14096 9324 14148 9376
rect 15936 9324 15988 9376
rect 17684 9324 17736 9376
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 19616 9324 19668 9376
rect 20168 9324 20220 9376
rect 21916 9596 21968 9648
rect 22468 9596 22520 9648
rect 22744 9596 22796 9648
rect 24124 9664 24176 9716
rect 24308 9664 24360 9716
rect 26608 9664 26660 9716
rect 27252 9664 27304 9716
rect 23572 9596 23624 9648
rect 25412 9596 25464 9648
rect 27804 9664 27856 9716
rect 27896 9664 27948 9716
rect 27436 9596 27488 9648
rect 21272 9503 21324 9512
rect 21272 9469 21281 9503
rect 21281 9469 21315 9503
rect 21315 9469 21324 9503
rect 21272 9460 21324 9469
rect 21916 9503 21968 9512
rect 21916 9469 21925 9503
rect 21925 9469 21959 9503
rect 21959 9469 21968 9503
rect 21916 9460 21968 9469
rect 22100 9460 22152 9512
rect 22284 9460 22336 9512
rect 23480 9460 23532 9512
rect 23664 9460 23716 9512
rect 23848 9460 23900 9512
rect 24768 9503 24820 9512
rect 21180 9324 21232 9376
rect 22928 9435 22980 9444
rect 22928 9401 22937 9435
rect 22937 9401 22971 9435
rect 22971 9401 22980 9435
rect 22928 9392 22980 9401
rect 23388 9392 23440 9444
rect 23940 9435 23992 9444
rect 23940 9401 23949 9435
rect 23949 9401 23983 9435
rect 23983 9401 23992 9435
rect 23940 9392 23992 9401
rect 24768 9469 24777 9503
rect 24777 9469 24811 9503
rect 24811 9469 24820 9503
rect 24768 9460 24820 9469
rect 25228 9460 25280 9512
rect 24584 9435 24636 9444
rect 24584 9401 24593 9435
rect 24593 9401 24627 9435
rect 24627 9401 24636 9435
rect 24584 9392 24636 9401
rect 25136 9392 25188 9444
rect 25688 9503 25740 9512
rect 25688 9469 25697 9503
rect 25697 9469 25731 9503
rect 25731 9469 25740 9503
rect 25688 9460 25740 9469
rect 24400 9367 24452 9376
rect 24400 9333 24409 9367
rect 24409 9333 24443 9367
rect 24443 9333 24452 9367
rect 24400 9324 24452 9333
rect 25412 9367 25464 9376
rect 25412 9333 25421 9367
rect 25421 9333 25455 9367
rect 25455 9333 25464 9367
rect 25412 9324 25464 9333
rect 25872 9324 25924 9376
rect 26240 9435 26292 9444
rect 26240 9401 26249 9435
rect 26249 9401 26283 9435
rect 26283 9401 26292 9435
rect 26240 9392 26292 9401
rect 26332 9392 26384 9444
rect 26608 9503 26660 9512
rect 26608 9469 26617 9503
rect 26617 9469 26651 9503
rect 26651 9469 26660 9503
rect 26608 9460 26660 9469
rect 27712 9571 27764 9580
rect 27712 9537 27721 9571
rect 27721 9537 27755 9571
rect 27755 9537 27764 9571
rect 27712 9528 27764 9537
rect 29460 9664 29512 9716
rect 29644 9664 29696 9716
rect 29000 9596 29052 9648
rect 28172 9528 28224 9580
rect 26976 9435 27028 9444
rect 26976 9401 26985 9435
rect 26985 9401 27019 9435
rect 27019 9401 27028 9435
rect 26976 9392 27028 9401
rect 26884 9324 26936 9376
rect 27068 9367 27120 9376
rect 27068 9333 27077 9367
rect 27077 9333 27111 9367
rect 27111 9333 27120 9367
rect 27068 9324 27120 9333
rect 28264 9460 28316 9512
rect 27620 9392 27672 9444
rect 28540 9528 28592 9580
rect 28448 9503 28500 9512
rect 28448 9469 28457 9503
rect 28457 9469 28491 9503
rect 28491 9469 28500 9503
rect 28448 9460 28500 9469
rect 28724 9460 28776 9512
rect 29552 9460 29604 9512
rect 30472 9528 30524 9580
rect 29184 9435 29236 9444
rect 29184 9401 29189 9435
rect 29189 9401 29223 9435
rect 29223 9401 29236 9435
rect 29184 9392 29236 9401
rect 30380 9460 30432 9512
rect 30656 9460 30708 9512
rect 31208 9503 31260 9512
rect 31208 9469 31217 9503
rect 31217 9469 31251 9503
rect 31251 9469 31260 9503
rect 31208 9460 31260 9469
rect 30288 9392 30340 9444
rect 27528 9324 27580 9376
rect 27804 9324 27856 9376
rect 28356 9324 28408 9376
rect 28908 9324 28960 9376
rect 29000 9324 29052 9376
rect 30104 9324 30156 9376
rect 6946 9222 6998 9274
rect 7010 9222 7062 9274
rect 7074 9222 7126 9274
rect 7138 9222 7190 9274
rect 7202 9222 7254 9274
rect 14306 9222 14358 9274
rect 14370 9222 14422 9274
rect 14434 9222 14486 9274
rect 14498 9222 14550 9274
rect 14562 9222 14614 9274
rect 21666 9222 21718 9274
rect 21730 9222 21782 9274
rect 21794 9222 21846 9274
rect 21858 9222 21910 9274
rect 21922 9222 21974 9274
rect 29026 9222 29078 9274
rect 29090 9222 29142 9274
rect 29154 9222 29206 9274
rect 29218 9222 29270 9274
rect 29282 9222 29334 9274
rect 6736 9120 6788 9172
rect 7472 9120 7524 9172
rect 14096 9120 14148 9172
rect 15844 9120 15896 9172
rect 16672 9120 16724 9172
rect 18604 9120 18656 9172
rect 14372 9095 14424 9104
rect 14372 9061 14381 9095
rect 14381 9061 14415 9095
rect 14415 9061 14424 9095
rect 14372 9052 14424 9061
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 14004 9027 14056 9036
rect 14004 8993 14013 9027
rect 14013 8993 14047 9027
rect 14047 8993 14056 9027
rect 14004 8984 14056 8993
rect 16672 8984 16724 9036
rect 11612 8959 11664 8968
rect 11612 8925 11621 8959
rect 11621 8925 11655 8959
rect 11655 8925 11664 8959
rect 11612 8916 11664 8925
rect 11704 8959 11756 8968
rect 11704 8925 11738 8959
rect 11738 8925 11756 8959
rect 11704 8916 11756 8925
rect 13544 8916 13596 8968
rect 14096 8916 14148 8968
rect 14648 8959 14700 8968
rect 14648 8925 14657 8959
rect 14657 8925 14691 8959
rect 14691 8925 14700 8959
rect 14648 8916 14700 8925
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 16304 8916 16356 8968
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 17960 9052 18012 9104
rect 18972 9052 19024 9104
rect 18512 9027 18564 9036
rect 18512 8993 18521 9027
rect 18521 8993 18555 9027
rect 18555 8993 18564 9027
rect 18512 8984 18564 8993
rect 19616 9052 19668 9104
rect 20720 9052 20772 9104
rect 21272 9052 21324 9104
rect 18788 8916 18840 8968
rect 19248 8959 19300 8968
rect 19248 8925 19257 8959
rect 19257 8925 19291 8959
rect 19291 8925 19300 8959
rect 19248 8916 19300 8925
rect 23940 9120 23992 9172
rect 25412 9120 25464 9172
rect 26608 9163 26660 9172
rect 24400 9052 24452 9104
rect 21456 9027 21508 9036
rect 21456 8993 21465 9027
rect 21465 8993 21499 9027
rect 21499 8993 21508 9027
rect 21456 8984 21508 8993
rect 23848 8984 23900 9036
rect 24768 9027 24820 9036
rect 24768 8993 24777 9027
rect 24777 8993 24811 9027
rect 24811 8993 24820 9027
rect 24768 8984 24820 8993
rect 24952 8984 25004 9036
rect 25688 9027 25740 9036
rect 25688 8993 25697 9027
rect 25697 8993 25731 9027
rect 25731 8993 25740 9027
rect 25688 8984 25740 8993
rect 26608 9129 26617 9163
rect 26617 9129 26651 9163
rect 26651 9129 26660 9163
rect 26608 9120 26660 9129
rect 27068 9120 27120 9172
rect 27252 9120 27304 9172
rect 27436 9163 27488 9172
rect 27436 9129 27445 9163
rect 27445 9129 27479 9163
rect 27479 9129 27488 9163
rect 27436 9120 27488 9129
rect 27804 9163 27856 9172
rect 27804 9129 27813 9163
rect 27813 9129 27847 9163
rect 27847 9129 27856 9163
rect 27804 9120 27856 9129
rect 27896 9120 27948 9172
rect 28356 9120 28408 9172
rect 28448 9120 28500 9172
rect 29552 9120 29604 9172
rect 29460 9052 29512 9104
rect 30104 9120 30156 9172
rect 31208 9120 31260 9172
rect 31116 9052 31168 9104
rect 26424 9027 26476 9036
rect 26424 8993 26433 9027
rect 26433 8993 26467 9027
rect 26467 8993 26476 9027
rect 26424 8984 26476 8993
rect 26608 8984 26660 9036
rect 14004 8780 14056 8832
rect 14648 8780 14700 8832
rect 17960 8848 18012 8900
rect 18880 8848 18932 8900
rect 24308 8916 24360 8968
rect 24676 8916 24728 8968
rect 25872 8959 25924 8968
rect 25872 8925 25881 8959
rect 25881 8925 25915 8959
rect 25915 8925 25924 8959
rect 25872 8916 25924 8925
rect 33140 9052 33192 9104
rect 28080 8916 28132 8968
rect 28632 8959 28684 8968
rect 28632 8925 28641 8959
rect 28641 8925 28675 8959
rect 28675 8925 28684 8959
rect 28632 8916 28684 8925
rect 28908 8916 28960 8968
rect 15016 8780 15068 8832
rect 15384 8780 15436 8832
rect 16120 8780 16172 8832
rect 16488 8823 16540 8832
rect 16488 8789 16497 8823
rect 16497 8789 16531 8823
rect 16531 8789 16540 8823
rect 16488 8780 16540 8789
rect 16948 8780 17000 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 18696 8823 18748 8832
rect 18696 8789 18705 8823
rect 18705 8789 18739 8823
rect 18739 8789 18748 8823
rect 18696 8780 18748 8789
rect 21180 8780 21232 8832
rect 21732 8780 21784 8832
rect 21916 8780 21968 8832
rect 23756 8780 23808 8832
rect 25228 8780 25280 8832
rect 25780 8780 25832 8832
rect 27068 8848 27120 8900
rect 28448 8848 28500 8900
rect 29368 8916 29420 8968
rect 29460 8848 29512 8900
rect 31668 8891 31720 8900
rect 31668 8857 31677 8891
rect 31677 8857 31711 8891
rect 31711 8857 31720 8891
rect 31668 8848 31720 8857
rect 26148 8823 26200 8832
rect 26148 8789 26157 8823
rect 26157 8789 26191 8823
rect 26191 8789 26200 8823
rect 26148 8780 26200 8789
rect 26332 8780 26384 8832
rect 27528 8780 27580 8832
rect 27620 8780 27672 8832
rect 29276 8823 29328 8832
rect 29276 8789 29285 8823
rect 29285 8789 29319 8823
rect 29319 8789 29328 8823
rect 29276 8780 29328 8789
rect 29644 8780 29696 8832
rect 30288 8780 30340 8832
rect 31484 8823 31536 8832
rect 31484 8789 31493 8823
rect 31493 8789 31527 8823
rect 31527 8789 31536 8823
rect 31484 8780 31536 8789
rect 6286 8678 6338 8730
rect 6350 8678 6402 8730
rect 6414 8678 6466 8730
rect 6478 8678 6530 8730
rect 6542 8678 6594 8730
rect 13646 8678 13698 8730
rect 13710 8678 13762 8730
rect 13774 8678 13826 8730
rect 13838 8678 13890 8730
rect 13902 8678 13954 8730
rect 21006 8678 21058 8730
rect 21070 8678 21122 8730
rect 21134 8678 21186 8730
rect 21198 8678 21250 8730
rect 21262 8678 21314 8730
rect 28366 8678 28418 8730
rect 28430 8678 28482 8730
rect 28494 8678 28546 8730
rect 28558 8678 28610 8730
rect 28622 8678 28674 8730
rect 3332 8576 3384 8628
rect 6736 8440 6788 8492
rect 14372 8576 14424 8628
rect 14740 8576 14792 8628
rect 14924 8619 14976 8628
rect 14924 8585 14933 8619
rect 14933 8585 14967 8619
rect 14967 8585 14976 8619
rect 14924 8576 14976 8585
rect 15844 8576 15896 8628
rect 16488 8576 16540 8628
rect 16948 8576 17000 8628
rect 18328 8576 18380 8628
rect 18696 8576 18748 8628
rect 19248 8576 19300 8628
rect 21364 8576 21416 8628
rect 21916 8576 21968 8628
rect 22008 8576 22060 8628
rect 14004 8508 14056 8560
rect 8300 8372 8352 8424
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 13820 8415 13872 8424
rect 13820 8381 13829 8415
rect 13829 8381 13863 8415
rect 13863 8381 13872 8415
rect 13820 8372 13872 8381
rect 14924 8372 14976 8424
rect 16028 8372 16080 8424
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 18972 8508 19024 8560
rect 18880 8440 18932 8492
rect 18788 8415 18840 8424
rect 18788 8381 18797 8415
rect 18797 8381 18831 8415
rect 18831 8381 18840 8415
rect 18788 8372 18840 8381
rect 4252 8236 4304 8288
rect 6184 8236 6236 8288
rect 13544 8236 13596 8288
rect 14832 8236 14884 8288
rect 15752 8279 15804 8288
rect 15752 8245 15761 8279
rect 15761 8245 15795 8279
rect 15795 8245 15804 8279
rect 15752 8236 15804 8245
rect 16580 8304 16632 8356
rect 18236 8304 18288 8356
rect 19708 8304 19760 8356
rect 19248 8279 19300 8288
rect 19248 8245 19257 8279
rect 19257 8245 19291 8279
rect 19291 8245 19300 8279
rect 19248 8236 19300 8245
rect 20352 8372 20404 8424
rect 22192 8440 22244 8492
rect 21732 8415 21784 8424
rect 21732 8381 21741 8415
rect 21741 8381 21775 8415
rect 21775 8381 21784 8415
rect 21732 8372 21784 8381
rect 25136 8576 25188 8628
rect 25688 8576 25740 8628
rect 27896 8619 27948 8628
rect 27896 8585 27905 8619
rect 27905 8585 27939 8619
rect 27939 8585 27948 8619
rect 27896 8576 27948 8585
rect 27988 8576 28040 8628
rect 28816 8576 28868 8628
rect 29736 8576 29788 8628
rect 30656 8576 30708 8628
rect 31116 8576 31168 8628
rect 26884 8508 26936 8560
rect 27528 8508 27580 8560
rect 29644 8551 29696 8560
rect 29644 8517 29653 8551
rect 29653 8517 29687 8551
rect 29687 8517 29696 8551
rect 29644 8508 29696 8517
rect 20904 8304 20956 8356
rect 20444 8236 20496 8288
rect 21548 8304 21600 8356
rect 22008 8304 22060 8356
rect 24676 8440 24728 8492
rect 26148 8483 26200 8492
rect 26148 8449 26157 8483
rect 26157 8449 26191 8483
rect 26191 8449 26200 8483
rect 26148 8440 26200 8449
rect 27068 8483 27120 8492
rect 27068 8449 27077 8483
rect 27077 8449 27111 8483
rect 27111 8449 27120 8483
rect 27068 8440 27120 8449
rect 23296 8415 23348 8424
rect 23296 8381 23305 8415
rect 23305 8381 23339 8415
rect 23339 8381 23348 8415
rect 23296 8372 23348 8381
rect 24308 8372 24360 8424
rect 24584 8372 24636 8424
rect 22192 8236 22244 8288
rect 23112 8279 23164 8288
rect 23112 8245 23121 8279
rect 23121 8245 23155 8279
rect 23155 8245 23164 8279
rect 23112 8236 23164 8245
rect 23388 8236 23440 8288
rect 25320 8415 25372 8424
rect 25320 8381 25329 8415
rect 25329 8381 25363 8415
rect 25363 8381 25372 8415
rect 25320 8372 25372 8381
rect 25872 8415 25924 8424
rect 25872 8381 25881 8415
rect 25881 8381 25915 8415
rect 25915 8381 25924 8415
rect 25872 8372 25924 8381
rect 26976 8415 27028 8424
rect 26976 8381 26985 8415
rect 26985 8381 27019 8415
rect 27019 8381 27028 8415
rect 26976 8372 27028 8381
rect 26608 8304 26660 8356
rect 27528 8372 27580 8424
rect 28080 8415 28132 8424
rect 28080 8381 28089 8415
rect 28089 8381 28123 8415
rect 28123 8381 28132 8415
rect 28080 8372 28132 8381
rect 28448 8372 28500 8424
rect 28724 8372 28776 8424
rect 29276 8372 29328 8424
rect 29460 8372 29512 8424
rect 29828 8372 29880 8424
rect 30288 8372 30340 8424
rect 29644 8304 29696 8356
rect 30656 8415 30708 8424
rect 30656 8381 30665 8415
rect 30665 8381 30699 8415
rect 30699 8381 30708 8415
rect 30656 8372 30708 8381
rect 30840 8415 30892 8424
rect 30840 8381 30849 8415
rect 30849 8381 30883 8415
rect 30883 8381 30892 8415
rect 30840 8372 30892 8381
rect 31116 8372 31168 8424
rect 31208 8372 31260 8424
rect 31392 8415 31444 8424
rect 31392 8381 31401 8415
rect 31401 8381 31435 8415
rect 31435 8381 31444 8415
rect 31392 8372 31444 8381
rect 31484 8372 31536 8424
rect 25780 8279 25832 8288
rect 25780 8245 25789 8279
rect 25789 8245 25823 8279
rect 25823 8245 25832 8279
rect 25780 8236 25832 8245
rect 26700 8279 26752 8288
rect 26700 8245 26709 8279
rect 26709 8245 26743 8279
rect 26743 8245 26752 8279
rect 26700 8236 26752 8245
rect 27436 8236 27488 8288
rect 28264 8236 28316 8288
rect 28724 8279 28776 8288
rect 28724 8245 28733 8279
rect 28733 8245 28767 8279
rect 28767 8245 28776 8279
rect 28724 8236 28776 8245
rect 28816 8236 28868 8288
rect 29460 8279 29512 8288
rect 29460 8245 29469 8279
rect 29469 8245 29503 8279
rect 29503 8245 29512 8279
rect 29460 8236 29512 8245
rect 30472 8236 30524 8288
rect 30564 8236 30616 8288
rect 6946 8134 6998 8186
rect 7010 8134 7062 8186
rect 7074 8134 7126 8186
rect 7138 8134 7190 8186
rect 7202 8134 7254 8186
rect 14306 8134 14358 8186
rect 14370 8134 14422 8186
rect 14434 8134 14486 8186
rect 14498 8134 14550 8186
rect 14562 8134 14614 8186
rect 21666 8134 21718 8186
rect 21730 8134 21782 8186
rect 21794 8134 21846 8186
rect 21858 8134 21910 8186
rect 21922 8134 21974 8186
rect 29026 8134 29078 8186
rect 29090 8134 29142 8186
rect 29154 8134 29206 8186
rect 29218 8134 29270 8186
rect 29282 8134 29334 8186
rect 3240 8032 3292 8084
rect 14188 8032 14240 8084
rect 1308 7896 1360 7948
rect 6092 7828 6144 7880
rect 6184 7828 6236 7880
rect 14188 7939 14240 7948
rect 14188 7905 14222 7939
rect 14222 7905 14240 7939
rect 14188 7896 14240 7905
rect 15752 7896 15804 7948
rect 18052 8032 18104 8084
rect 19248 8032 19300 8084
rect 16580 7964 16632 8016
rect 16764 7964 16816 8016
rect 18420 7964 18472 8016
rect 22100 7964 22152 8016
rect 23296 8032 23348 8084
rect 26424 8032 26476 8084
rect 18328 7939 18380 7948
rect 18328 7905 18337 7939
rect 18337 7905 18371 7939
rect 18371 7905 18380 7939
rect 18328 7896 18380 7905
rect 20168 7939 20220 7948
rect 20168 7905 20202 7939
rect 20202 7905 20220 7939
rect 20168 7896 20220 7905
rect 20352 7939 20404 7948
rect 20352 7905 20361 7939
rect 20361 7905 20395 7939
rect 20395 7905 20404 7939
rect 20352 7896 20404 7905
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 13912 7828 13964 7880
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 6828 7760 6880 7812
rect 13728 7692 13780 7744
rect 15200 7828 15252 7880
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 19340 7871 19392 7880
rect 19340 7837 19349 7871
rect 19349 7837 19383 7871
rect 19383 7837 19392 7871
rect 19340 7828 19392 7837
rect 20076 7871 20128 7880
rect 20076 7837 20085 7871
rect 20085 7837 20119 7871
rect 20119 7837 20128 7871
rect 20076 7828 20128 7837
rect 21916 7828 21968 7880
rect 15568 7760 15620 7812
rect 14188 7692 14240 7744
rect 14740 7692 14792 7744
rect 14832 7692 14884 7744
rect 15292 7735 15344 7744
rect 15292 7701 15301 7735
rect 15301 7701 15335 7735
rect 15335 7701 15344 7735
rect 15292 7692 15344 7701
rect 20904 7692 20956 7744
rect 22560 7939 22612 7948
rect 22560 7905 22569 7939
rect 22569 7905 22603 7939
rect 22603 7905 22612 7939
rect 22560 7896 22612 7905
rect 25780 7964 25832 8016
rect 26700 8032 26752 8084
rect 28080 8032 28132 8084
rect 28724 8032 28776 8084
rect 23020 7896 23072 7948
rect 23112 7896 23164 7948
rect 23480 7828 23532 7880
rect 22928 7760 22980 7812
rect 24768 7896 24820 7948
rect 27620 7896 27672 7948
rect 28172 7896 28224 7948
rect 29920 8032 29972 8084
rect 30564 8032 30616 8084
rect 29460 7964 29512 8016
rect 30380 7964 30432 8016
rect 31116 8032 31168 8084
rect 22468 7735 22520 7744
rect 22468 7701 22477 7735
rect 22477 7701 22511 7735
rect 22511 7701 22520 7735
rect 22468 7692 22520 7701
rect 24124 7692 24176 7744
rect 24492 7735 24544 7744
rect 24492 7701 24501 7735
rect 24501 7701 24535 7735
rect 24535 7701 24544 7735
rect 24492 7692 24544 7701
rect 26332 7692 26384 7744
rect 27436 7871 27488 7880
rect 27436 7837 27445 7871
rect 27445 7837 27479 7871
rect 27479 7837 27488 7871
rect 27436 7828 27488 7837
rect 27712 7871 27764 7880
rect 27712 7837 27721 7871
rect 27721 7837 27755 7871
rect 27755 7837 27764 7871
rect 27712 7828 27764 7837
rect 27804 7828 27856 7880
rect 29736 7896 29788 7948
rect 30748 7896 30800 7948
rect 30840 7939 30892 7948
rect 30840 7905 30849 7939
rect 30849 7905 30883 7939
rect 30883 7905 30892 7939
rect 30840 7896 30892 7905
rect 33140 7896 33192 7948
rect 26976 7760 27028 7812
rect 26884 7735 26936 7744
rect 26884 7701 26893 7735
rect 26893 7701 26927 7735
rect 26927 7701 26936 7735
rect 26884 7692 26936 7701
rect 28724 7735 28776 7744
rect 28724 7701 28733 7735
rect 28733 7701 28767 7735
rect 28767 7701 28776 7735
rect 28724 7692 28776 7701
rect 29460 7692 29512 7744
rect 29644 7692 29696 7744
rect 30104 7735 30156 7744
rect 30104 7701 30113 7735
rect 30113 7701 30147 7735
rect 30147 7701 30156 7735
rect 30104 7692 30156 7701
rect 31668 7735 31720 7744
rect 31668 7701 31677 7735
rect 31677 7701 31711 7735
rect 31711 7701 31720 7735
rect 31668 7692 31720 7701
rect 6286 7590 6338 7642
rect 6350 7590 6402 7642
rect 6414 7590 6466 7642
rect 6478 7590 6530 7642
rect 6542 7590 6594 7642
rect 13646 7590 13698 7642
rect 13710 7590 13762 7642
rect 13774 7590 13826 7642
rect 13838 7590 13890 7642
rect 13902 7590 13954 7642
rect 21006 7590 21058 7642
rect 21070 7590 21122 7642
rect 21134 7590 21186 7642
rect 21198 7590 21250 7642
rect 21262 7590 21314 7642
rect 28366 7590 28418 7642
rect 28430 7590 28482 7642
rect 28494 7590 28546 7642
rect 28558 7590 28610 7642
rect 28622 7590 28674 7642
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 9404 7488 9456 7540
rect 13268 7531 13320 7540
rect 13268 7497 13277 7531
rect 13277 7497 13311 7531
rect 13311 7497 13320 7531
rect 13268 7488 13320 7497
rect 13636 7488 13688 7540
rect 15292 7488 15344 7540
rect 15108 7420 15160 7472
rect 16672 7488 16724 7540
rect 17960 7488 18012 7540
rect 18236 7488 18288 7540
rect 22560 7488 22612 7540
rect 23388 7531 23440 7540
rect 23388 7497 23397 7531
rect 23397 7497 23431 7531
rect 23431 7497 23440 7531
rect 23388 7488 23440 7497
rect 27712 7488 27764 7540
rect 28724 7488 28776 7540
rect 15200 7284 15252 7336
rect 14096 7216 14148 7268
rect 13176 7148 13228 7200
rect 21456 7352 21508 7404
rect 21916 7352 21968 7404
rect 15660 7216 15712 7268
rect 16764 7284 16816 7336
rect 17040 7284 17092 7336
rect 17316 7327 17368 7336
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 18512 7327 18564 7336
rect 18512 7293 18521 7327
rect 18521 7293 18555 7327
rect 18555 7293 18564 7327
rect 18512 7284 18564 7293
rect 24124 7327 24176 7336
rect 24124 7293 24133 7327
rect 24133 7293 24167 7327
rect 24167 7293 24176 7327
rect 24124 7284 24176 7293
rect 18236 7216 18288 7268
rect 22192 7216 22244 7268
rect 22652 7216 22704 7268
rect 24492 7216 24544 7268
rect 28264 7284 28316 7336
rect 16764 7191 16816 7200
rect 16764 7157 16773 7191
rect 16773 7157 16807 7191
rect 16807 7157 16816 7191
rect 16764 7148 16816 7157
rect 20444 7148 20496 7200
rect 22560 7148 22612 7200
rect 25320 7148 25372 7200
rect 25780 7148 25832 7200
rect 26240 7216 26292 7268
rect 26332 7259 26384 7268
rect 26332 7225 26341 7259
rect 26341 7225 26375 7259
rect 26375 7225 26384 7259
rect 26332 7216 26384 7225
rect 27620 7216 27672 7268
rect 28448 7327 28500 7336
rect 28448 7293 28457 7327
rect 28457 7293 28491 7327
rect 28491 7293 28500 7327
rect 28448 7284 28500 7293
rect 28908 7488 28960 7540
rect 30104 7488 30156 7540
rect 30840 7531 30892 7540
rect 30840 7497 30849 7531
rect 30849 7497 30883 7531
rect 30883 7497 30892 7531
rect 30840 7488 30892 7497
rect 29000 7284 29052 7336
rect 29368 7352 29420 7404
rect 30472 7284 30524 7336
rect 26976 7148 27028 7200
rect 27252 7148 27304 7200
rect 28724 7216 28776 7268
rect 29368 7148 29420 7200
rect 29736 7148 29788 7200
rect 6946 7046 6998 7098
rect 7010 7046 7062 7098
rect 7074 7046 7126 7098
rect 7138 7046 7190 7098
rect 7202 7046 7254 7098
rect 14306 7046 14358 7098
rect 14370 7046 14422 7098
rect 14434 7046 14486 7098
rect 14498 7046 14550 7098
rect 14562 7046 14614 7098
rect 21666 7046 21718 7098
rect 21730 7046 21782 7098
rect 21794 7046 21846 7098
rect 21858 7046 21910 7098
rect 21922 7046 21974 7098
rect 29026 7046 29078 7098
rect 29090 7046 29142 7098
rect 29154 7046 29206 7098
rect 29218 7046 29270 7098
rect 29282 7046 29334 7098
rect 7656 6876 7708 6928
rect 7196 6851 7248 6860
rect 7196 6817 7205 6851
rect 7205 6817 7239 6851
rect 7239 6817 7248 6851
rect 7196 6808 7248 6817
rect 11888 6808 11940 6860
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 9404 6740 9456 6792
rect 13544 6944 13596 6996
rect 15476 6944 15528 6996
rect 15568 6944 15620 6996
rect 16304 6987 16356 6996
rect 16304 6953 16313 6987
rect 16313 6953 16347 6987
rect 16347 6953 16356 6987
rect 16304 6944 16356 6953
rect 19340 6944 19392 6996
rect 22652 6944 22704 6996
rect 23480 6987 23532 6996
rect 23480 6953 23489 6987
rect 23489 6953 23523 6987
rect 23523 6953 23532 6987
rect 23480 6944 23532 6953
rect 26332 6944 26384 6996
rect 26884 6944 26936 6996
rect 27620 6987 27672 6996
rect 27620 6953 27629 6987
rect 27629 6953 27663 6987
rect 27663 6953 27672 6987
rect 27620 6944 27672 6953
rect 27804 6944 27856 6996
rect 28356 6944 28408 6996
rect 12532 6876 12584 6928
rect 15200 6876 15252 6928
rect 15384 6919 15436 6928
rect 15384 6885 15393 6919
rect 15393 6885 15427 6919
rect 15427 6885 15436 6919
rect 15384 6876 15436 6885
rect 16764 6876 16816 6928
rect 20076 6876 20128 6928
rect 13268 6808 13320 6860
rect 13452 6851 13504 6860
rect 13452 6817 13461 6851
rect 13461 6817 13495 6851
rect 13495 6817 13504 6851
rect 13452 6808 13504 6817
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 13636 6808 13688 6860
rect 14648 6808 14700 6860
rect 14924 6851 14976 6860
rect 14924 6817 14933 6851
rect 14933 6817 14967 6851
rect 14967 6817 14976 6851
rect 14924 6808 14976 6817
rect 15016 6851 15068 6860
rect 15016 6817 15025 6851
rect 15025 6817 15059 6851
rect 15059 6817 15068 6851
rect 15016 6808 15068 6817
rect 16396 6851 16448 6860
rect 16396 6817 16405 6851
rect 16405 6817 16439 6851
rect 16439 6817 16448 6851
rect 16396 6808 16448 6817
rect 18420 6808 18472 6860
rect 15016 6672 15068 6724
rect 16672 6740 16724 6792
rect 13176 6647 13228 6656
rect 13176 6613 13185 6647
rect 13185 6613 13219 6647
rect 13219 6613 13228 6647
rect 13176 6604 13228 6613
rect 14832 6604 14884 6656
rect 15292 6604 15344 6656
rect 15936 6672 15988 6724
rect 16212 6604 16264 6656
rect 17960 6672 18012 6724
rect 20628 6808 20680 6860
rect 21548 6808 21600 6860
rect 22928 6876 22980 6928
rect 23848 6851 23900 6860
rect 23848 6817 23857 6851
rect 23857 6817 23891 6851
rect 23891 6817 23900 6851
rect 23848 6808 23900 6817
rect 20444 6783 20496 6792
rect 20444 6749 20453 6783
rect 20453 6749 20487 6783
rect 20487 6749 20496 6783
rect 20444 6740 20496 6749
rect 20720 6740 20772 6792
rect 23388 6740 23440 6792
rect 20260 6672 20312 6724
rect 28724 6944 28776 6996
rect 27620 6808 27672 6860
rect 28264 6851 28316 6860
rect 28264 6817 28273 6851
rect 28273 6817 28307 6851
rect 28307 6817 28316 6851
rect 28264 6808 28316 6817
rect 27896 6740 27948 6792
rect 17684 6604 17736 6656
rect 19064 6647 19116 6656
rect 19064 6613 19073 6647
rect 19073 6613 19107 6647
rect 19107 6613 19116 6647
rect 19064 6604 19116 6613
rect 24676 6647 24728 6656
rect 24676 6613 24685 6647
rect 24685 6613 24719 6647
rect 24719 6613 24728 6647
rect 24676 6604 24728 6613
rect 24952 6647 25004 6656
rect 24952 6613 24961 6647
rect 24961 6613 24995 6647
rect 24995 6613 25004 6647
rect 24952 6604 25004 6613
rect 25044 6604 25096 6656
rect 28724 6740 28776 6792
rect 29828 6740 29880 6792
rect 30656 6783 30708 6792
rect 30656 6749 30665 6783
rect 30665 6749 30699 6783
rect 30699 6749 30708 6783
rect 30656 6740 30708 6749
rect 28816 6604 28868 6656
rect 30104 6647 30156 6656
rect 30104 6613 30113 6647
rect 30113 6613 30147 6647
rect 30147 6613 30156 6647
rect 30104 6604 30156 6613
rect 6286 6502 6338 6554
rect 6350 6502 6402 6554
rect 6414 6502 6466 6554
rect 6478 6502 6530 6554
rect 6542 6502 6594 6554
rect 13646 6502 13698 6554
rect 13710 6502 13762 6554
rect 13774 6502 13826 6554
rect 13838 6502 13890 6554
rect 13902 6502 13954 6554
rect 21006 6502 21058 6554
rect 21070 6502 21122 6554
rect 21134 6502 21186 6554
rect 21198 6502 21250 6554
rect 21262 6502 21314 6554
rect 28366 6502 28418 6554
rect 28430 6502 28482 6554
rect 28494 6502 28546 6554
rect 28558 6502 28610 6554
rect 28622 6502 28674 6554
rect 6920 6400 6972 6452
rect 13176 6400 13228 6452
rect 15016 6400 15068 6452
rect 15936 6400 15988 6452
rect 17316 6400 17368 6452
rect 18420 6443 18472 6452
rect 18420 6409 18429 6443
rect 18429 6409 18463 6443
rect 18463 6409 18472 6443
rect 18420 6400 18472 6409
rect 19064 6400 19116 6452
rect 20720 6443 20772 6452
rect 20720 6409 20729 6443
rect 20729 6409 20763 6443
rect 20763 6409 20772 6443
rect 20720 6400 20772 6409
rect 24676 6400 24728 6452
rect 28264 6400 28316 6452
rect 30104 6400 30156 6452
rect 30472 6443 30524 6452
rect 30472 6409 30481 6443
rect 30481 6409 30515 6443
rect 30515 6409 30524 6443
rect 30472 6400 30524 6409
rect 13268 6332 13320 6384
rect 16856 6332 16908 6384
rect 17684 6332 17736 6384
rect 18236 6332 18288 6384
rect 1308 6196 1360 6248
rect 5356 6196 5408 6248
rect 7840 6196 7892 6248
rect 9772 6239 9824 6248
rect 9772 6205 9781 6239
rect 9781 6205 9815 6239
rect 9815 6205 9824 6239
rect 9772 6196 9824 6205
rect 11612 6196 11664 6248
rect 6644 6103 6696 6112
rect 6644 6069 6653 6103
rect 6653 6069 6687 6103
rect 6687 6069 6696 6103
rect 6644 6060 6696 6069
rect 7196 6060 7248 6112
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 9036 6060 9088 6112
rect 14188 6196 14240 6248
rect 15292 6196 15344 6248
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 17316 6196 17368 6248
rect 17960 6196 18012 6248
rect 13912 6128 13964 6180
rect 14280 6128 14332 6180
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 12900 6103 12952 6112
rect 12900 6069 12909 6103
rect 12909 6069 12943 6103
rect 12943 6069 12952 6103
rect 12900 6060 12952 6069
rect 13544 6060 13596 6112
rect 14648 6060 14700 6112
rect 15752 6103 15804 6112
rect 15752 6069 15761 6103
rect 15761 6069 15795 6103
rect 15795 6069 15804 6103
rect 15752 6060 15804 6069
rect 16856 6128 16908 6180
rect 16580 6060 16632 6112
rect 18788 6196 18840 6248
rect 21548 6264 21600 6316
rect 22100 6264 22152 6316
rect 29828 6332 29880 6384
rect 26240 6264 26292 6316
rect 27620 6264 27672 6316
rect 28908 6264 28960 6316
rect 30012 6264 30064 6316
rect 23572 6196 23624 6248
rect 24584 6239 24636 6248
rect 24584 6205 24593 6239
rect 24593 6205 24627 6239
rect 24627 6205 24636 6239
rect 24584 6196 24636 6205
rect 27252 6128 27304 6180
rect 27712 6128 27764 6180
rect 29552 6128 29604 6180
rect 20260 6060 20312 6112
rect 23940 6103 23992 6112
rect 23940 6069 23949 6103
rect 23949 6069 23983 6103
rect 23983 6069 23992 6103
rect 23940 6060 23992 6069
rect 24032 6060 24084 6112
rect 29460 6060 29512 6112
rect 31208 6196 31260 6248
rect 33140 6196 33192 6248
rect 6946 5958 6998 6010
rect 7010 5958 7062 6010
rect 7074 5958 7126 6010
rect 7138 5958 7190 6010
rect 7202 5958 7254 6010
rect 14306 5958 14358 6010
rect 14370 5958 14422 6010
rect 14434 5958 14486 6010
rect 14498 5958 14550 6010
rect 14562 5958 14614 6010
rect 21666 5958 21718 6010
rect 21730 5958 21782 6010
rect 21794 5958 21846 6010
rect 21858 5958 21910 6010
rect 21922 5958 21974 6010
rect 29026 5958 29078 6010
rect 29090 5958 29142 6010
rect 29154 5958 29206 6010
rect 29218 5958 29270 6010
rect 29282 5958 29334 6010
rect 6644 5856 6696 5908
rect 7840 5899 7892 5908
rect 7840 5865 7849 5899
rect 7849 5865 7883 5899
rect 7883 5865 7892 5899
rect 7840 5856 7892 5865
rect 9772 5856 9824 5908
rect 9956 5856 10008 5908
rect 12992 5899 13044 5908
rect 12992 5865 13001 5899
rect 13001 5865 13035 5899
rect 13035 5865 13044 5899
rect 12992 5856 13044 5865
rect 14832 5856 14884 5908
rect 15384 5856 15436 5908
rect 15752 5856 15804 5908
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 17684 5899 17736 5908
rect 17684 5865 17693 5899
rect 17693 5865 17727 5899
rect 17727 5865 17736 5899
rect 17684 5856 17736 5865
rect 18604 5899 18656 5908
rect 18604 5865 18613 5899
rect 18613 5865 18647 5899
rect 18647 5865 18656 5899
rect 18604 5856 18656 5865
rect 19064 5856 19116 5908
rect 20628 5899 20680 5908
rect 20628 5865 20637 5899
rect 20637 5865 20671 5899
rect 20671 5865 20680 5899
rect 20628 5856 20680 5865
rect 21548 5856 21600 5908
rect 23756 5899 23808 5908
rect 23756 5865 23765 5899
rect 23765 5865 23799 5899
rect 23799 5865 23808 5899
rect 23756 5856 23808 5865
rect 23848 5899 23900 5908
rect 23848 5865 23857 5899
rect 23857 5865 23891 5899
rect 23891 5865 23900 5899
rect 23848 5856 23900 5865
rect 23940 5856 23992 5908
rect 24584 5856 24636 5908
rect 25044 5899 25096 5908
rect 25044 5865 25053 5899
rect 25053 5865 25087 5899
rect 25087 5865 25096 5899
rect 25044 5856 25096 5865
rect 27712 5856 27764 5908
rect 28816 5856 28868 5908
rect 17132 5788 17184 5840
rect 18696 5788 18748 5840
rect 8208 5763 8260 5772
rect 8208 5729 8217 5763
rect 8217 5729 8251 5763
rect 8251 5729 8260 5763
rect 8208 5720 8260 5729
rect 10416 5720 10468 5772
rect 12808 5720 12860 5772
rect 14832 5763 14884 5772
rect 14832 5729 14841 5763
rect 14841 5729 14875 5763
rect 14875 5729 14884 5763
rect 14832 5720 14884 5729
rect 22560 5788 22612 5840
rect 22744 5831 22796 5840
rect 22744 5797 22753 5831
rect 22753 5797 22787 5831
rect 22787 5797 22796 5831
rect 22744 5788 22796 5797
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 5356 5652 5408 5661
rect 6092 5695 6144 5704
rect 6092 5661 6101 5695
rect 6101 5661 6135 5695
rect 6135 5661 6144 5695
rect 6092 5652 6144 5661
rect 6000 5559 6052 5568
rect 6000 5525 6009 5559
rect 6009 5525 6043 5559
rect 6043 5525 6052 5559
rect 6000 5516 6052 5525
rect 8300 5516 8352 5568
rect 9588 5652 9640 5704
rect 12992 5652 13044 5704
rect 13912 5652 13964 5704
rect 15016 5652 15068 5704
rect 15200 5652 15252 5704
rect 18788 5695 18840 5704
rect 18788 5661 18797 5695
rect 18797 5661 18831 5695
rect 18831 5661 18840 5695
rect 18788 5652 18840 5661
rect 19524 5652 19576 5704
rect 21640 5652 21692 5704
rect 24952 5788 25004 5840
rect 15476 5584 15528 5636
rect 21364 5584 21416 5636
rect 28172 5720 28224 5772
rect 28724 5720 28776 5772
rect 29552 5899 29604 5908
rect 29552 5865 29561 5899
rect 29561 5865 29595 5899
rect 29595 5865 29604 5899
rect 29552 5856 29604 5865
rect 30656 5856 30708 5908
rect 29460 5763 29512 5772
rect 29460 5729 29469 5763
rect 29469 5729 29503 5763
rect 29503 5729 29512 5763
rect 29460 5720 29512 5729
rect 25596 5695 25648 5704
rect 25596 5661 25605 5695
rect 25605 5661 25639 5695
rect 25639 5661 25648 5695
rect 25596 5652 25648 5661
rect 29368 5652 29420 5704
rect 14832 5516 14884 5568
rect 16028 5516 16080 5568
rect 18420 5516 18472 5568
rect 22376 5516 22428 5568
rect 22560 5559 22612 5568
rect 22560 5525 22569 5559
rect 22569 5525 22603 5559
rect 22603 5525 22612 5559
rect 22560 5516 22612 5525
rect 23664 5516 23716 5568
rect 24492 5516 24544 5568
rect 28724 5516 28776 5568
rect 29920 5516 29972 5568
rect 6286 5414 6338 5466
rect 6350 5414 6402 5466
rect 6414 5414 6466 5466
rect 6478 5414 6530 5466
rect 6542 5414 6594 5466
rect 13646 5414 13698 5466
rect 13710 5414 13762 5466
rect 13774 5414 13826 5466
rect 13838 5414 13890 5466
rect 13902 5414 13954 5466
rect 21006 5414 21058 5466
rect 21070 5414 21122 5466
rect 21134 5414 21186 5466
rect 21198 5414 21250 5466
rect 21262 5414 21314 5466
rect 28366 5414 28418 5466
rect 28430 5414 28482 5466
rect 28494 5414 28546 5466
rect 28558 5414 28610 5466
rect 28622 5414 28674 5466
rect 6736 5312 6788 5364
rect 8300 5312 8352 5364
rect 12992 5312 13044 5364
rect 7564 5244 7616 5296
rect 6092 5176 6144 5228
rect 9036 5176 9088 5228
rect 9588 5176 9640 5228
rect 12256 5176 12308 5228
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 12900 5176 12952 5228
rect 14188 5312 14240 5364
rect 16396 5312 16448 5364
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 17960 5312 18012 5364
rect 18052 5312 18104 5364
rect 19524 5355 19576 5364
rect 19524 5321 19533 5355
rect 19533 5321 19567 5355
rect 19567 5321 19576 5355
rect 19524 5312 19576 5321
rect 15200 5176 15252 5228
rect 4344 5151 4396 5160
rect 4344 5117 4353 5151
rect 4353 5117 4387 5151
rect 4387 5117 4396 5151
rect 4344 5108 4396 5117
rect 6000 5151 6052 5160
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 6920 5108 6972 5160
rect 1308 5040 1360 5092
rect 6828 5040 6880 5092
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 8208 5108 8260 5160
rect 14924 5108 14976 5160
rect 15752 5176 15804 5228
rect 15936 5176 15988 5228
rect 16304 5151 16356 5160
rect 16304 5117 16313 5151
rect 16313 5117 16347 5151
rect 16347 5117 16356 5151
rect 16304 5108 16356 5117
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 16856 5151 16908 5160
rect 16856 5117 16865 5151
rect 16865 5117 16899 5151
rect 16899 5117 16908 5151
rect 16856 5108 16908 5117
rect 18512 5176 18564 5228
rect 17040 5108 17092 5160
rect 18052 5151 18104 5160
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 18144 5108 18196 5160
rect 18328 5151 18380 5160
rect 18328 5117 18337 5151
rect 18337 5117 18371 5151
rect 18371 5117 18380 5151
rect 18328 5108 18380 5117
rect 18880 5108 18932 5160
rect 20076 5244 20128 5296
rect 19064 5219 19116 5228
rect 19064 5185 19073 5219
rect 19073 5185 19107 5219
rect 19107 5185 19116 5219
rect 19064 5176 19116 5185
rect 19248 5219 19300 5228
rect 19248 5185 19257 5219
rect 19257 5185 19291 5219
rect 19291 5185 19300 5219
rect 19248 5176 19300 5185
rect 21272 5312 21324 5364
rect 23940 5312 23992 5364
rect 24032 5312 24084 5364
rect 25596 5312 25648 5364
rect 20628 5151 20680 5160
rect 20628 5117 20637 5151
rect 20637 5117 20671 5151
rect 20671 5117 20680 5151
rect 20628 5108 20680 5117
rect 20720 5151 20772 5160
rect 20720 5117 20729 5151
rect 20729 5117 20763 5151
rect 20763 5117 20772 5151
rect 21640 5244 21692 5296
rect 21548 5176 21600 5228
rect 22100 5176 22152 5228
rect 24768 5244 24820 5296
rect 24216 5176 24268 5228
rect 20720 5108 20772 5117
rect 22008 5108 22060 5160
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 24124 5108 24176 5160
rect 9680 5040 9732 5092
rect 13544 5040 13596 5092
rect 6000 4972 6052 5024
rect 6644 4972 6696 5024
rect 10416 5015 10468 5024
rect 10416 4981 10425 5015
rect 10425 4981 10459 5015
rect 10459 4981 10468 5015
rect 10416 4972 10468 4981
rect 13452 4972 13504 5024
rect 21180 5040 21232 5092
rect 24676 5040 24728 5092
rect 23664 4972 23716 5024
rect 23756 4972 23808 5024
rect 24952 5151 25004 5160
rect 24952 5117 24961 5151
rect 24961 5117 24995 5151
rect 24995 5117 25004 5151
rect 24952 5108 25004 5117
rect 30012 5151 30064 5160
rect 30012 5117 30021 5151
rect 30021 5117 30055 5151
rect 30055 5117 30064 5151
rect 30012 5108 30064 5117
rect 24860 5040 24912 5092
rect 28540 5015 28592 5024
rect 28540 4981 28549 5015
rect 28549 4981 28583 5015
rect 28583 4981 28592 5015
rect 28540 4972 28592 4981
rect 29460 5015 29512 5024
rect 29460 4981 29469 5015
rect 29469 4981 29503 5015
rect 29503 4981 29512 5015
rect 29460 4972 29512 4981
rect 6946 4870 6998 4922
rect 7010 4870 7062 4922
rect 7074 4870 7126 4922
rect 7138 4870 7190 4922
rect 7202 4870 7254 4922
rect 14306 4870 14358 4922
rect 14370 4870 14422 4922
rect 14434 4870 14486 4922
rect 14498 4870 14550 4922
rect 14562 4870 14614 4922
rect 21666 4870 21718 4922
rect 21730 4870 21782 4922
rect 21794 4870 21846 4922
rect 21858 4870 21910 4922
rect 21922 4870 21974 4922
rect 29026 4870 29078 4922
rect 29090 4870 29142 4922
rect 29154 4870 29206 4922
rect 29218 4870 29270 4922
rect 29282 4870 29334 4922
rect 4436 4768 4488 4820
rect 5356 4768 5408 4820
rect 6828 4811 6880 4820
rect 6828 4777 6837 4811
rect 6837 4777 6871 4811
rect 6871 4777 6880 4811
rect 6828 4768 6880 4777
rect 9680 4768 9732 4820
rect 10232 4768 10284 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 12992 4811 13044 4820
rect 12992 4777 13001 4811
rect 13001 4777 13035 4811
rect 13035 4777 13044 4811
rect 12992 4768 13044 4777
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 13636 4768 13688 4820
rect 15292 4768 15344 4820
rect 17500 4768 17552 4820
rect 8208 4632 8260 4684
rect 6000 4564 6052 4616
rect 6092 4428 6144 4480
rect 6736 4564 6788 4616
rect 13544 4564 13596 4616
rect 14004 4564 14056 4616
rect 14188 4564 14240 4616
rect 15568 4632 15620 4684
rect 15108 4607 15160 4616
rect 15108 4573 15117 4607
rect 15117 4573 15151 4607
rect 15151 4573 15160 4607
rect 15108 4564 15160 4573
rect 15200 4607 15252 4616
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 16396 4632 16448 4684
rect 15200 4564 15252 4573
rect 16120 4607 16172 4616
rect 16120 4573 16129 4607
rect 16129 4573 16163 4607
rect 16163 4573 16172 4607
rect 16120 4564 16172 4573
rect 18052 4632 18104 4684
rect 18236 4632 18288 4684
rect 19064 4768 19116 4820
rect 21180 4768 21232 4820
rect 21456 4768 21508 4820
rect 22008 4768 22060 4820
rect 18420 4700 18472 4752
rect 18972 4700 19024 4752
rect 19800 4700 19852 4752
rect 18696 4675 18748 4684
rect 18696 4641 18705 4675
rect 18705 4641 18739 4675
rect 18739 4641 18748 4675
rect 18696 4632 18748 4641
rect 20720 4632 20772 4684
rect 23112 4700 23164 4752
rect 23572 4811 23624 4820
rect 23572 4777 23581 4811
rect 23581 4777 23615 4811
rect 23615 4777 23624 4811
rect 23572 4768 23624 4777
rect 23940 4768 23992 4820
rect 24952 4700 25004 4752
rect 29460 4768 29512 4820
rect 29736 4768 29788 4820
rect 21548 4675 21600 4684
rect 21548 4641 21557 4675
rect 21557 4641 21591 4675
rect 21591 4641 21600 4675
rect 21548 4632 21600 4641
rect 23480 4632 23532 4684
rect 24124 4632 24176 4684
rect 19432 4564 19484 4616
rect 20352 4564 20404 4616
rect 24032 4607 24084 4616
rect 24032 4573 24041 4607
rect 24041 4573 24075 4607
rect 24075 4573 24084 4607
rect 24032 4564 24084 4573
rect 19248 4496 19300 4548
rect 6736 4428 6788 4480
rect 14004 4428 14056 4480
rect 16212 4471 16264 4480
rect 16212 4437 16221 4471
rect 16221 4437 16255 4471
rect 16255 4437 16264 4471
rect 16212 4428 16264 4437
rect 19524 4428 19576 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 20260 4428 20312 4480
rect 20444 4471 20496 4480
rect 20444 4437 20453 4471
rect 20453 4437 20487 4471
rect 20487 4437 20496 4471
rect 20444 4428 20496 4437
rect 23388 4428 23440 4480
rect 23572 4428 23624 4480
rect 24492 4632 24544 4684
rect 28540 4632 28592 4684
rect 30840 4675 30892 4684
rect 30840 4641 30858 4675
rect 30858 4641 30892 4675
rect 30840 4632 30892 4641
rect 25412 4471 25464 4480
rect 25412 4437 25421 4471
rect 25421 4437 25455 4471
rect 25455 4437 25464 4471
rect 25412 4428 25464 4437
rect 28264 4428 28316 4480
rect 30472 4564 30524 4616
rect 30932 4607 30984 4616
rect 30932 4573 30941 4607
rect 30941 4573 30975 4607
rect 30975 4573 30984 4607
rect 30932 4564 30984 4573
rect 31668 4607 31720 4616
rect 31668 4573 31677 4607
rect 31677 4573 31711 4607
rect 31711 4573 31720 4607
rect 31668 4564 31720 4573
rect 31852 4607 31904 4616
rect 31852 4573 31861 4607
rect 31861 4573 31895 4607
rect 31895 4573 31904 4607
rect 31852 4564 31904 4573
rect 6286 4326 6338 4378
rect 6350 4326 6402 4378
rect 6414 4326 6466 4378
rect 6478 4326 6530 4378
rect 6542 4326 6594 4378
rect 13646 4326 13698 4378
rect 13710 4326 13762 4378
rect 13774 4326 13826 4378
rect 13838 4326 13890 4378
rect 13902 4326 13954 4378
rect 21006 4326 21058 4378
rect 21070 4326 21122 4378
rect 21134 4326 21186 4378
rect 21198 4326 21250 4378
rect 21262 4326 21314 4378
rect 28366 4326 28418 4378
rect 28430 4326 28482 4378
rect 28494 4326 28546 4378
rect 28558 4326 28610 4378
rect 28622 4326 28674 4378
rect 6736 4224 6788 4276
rect 7656 4224 7708 4276
rect 13452 4224 13504 4276
rect 14648 4224 14700 4276
rect 6092 4088 6144 4140
rect 12624 4088 12676 4140
rect 14096 4088 14148 4140
rect 16212 4224 16264 4276
rect 18052 4267 18104 4276
rect 18052 4233 18061 4267
rect 18061 4233 18095 4267
rect 18095 4233 18104 4267
rect 18052 4224 18104 4233
rect 17592 4156 17644 4208
rect 18880 4224 18932 4276
rect 19616 4224 19668 4276
rect 20076 4224 20128 4276
rect 3056 4063 3108 4072
rect 3056 4029 3065 4063
rect 3065 4029 3099 4063
rect 3099 4029 3108 4063
rect 3056 4020 3108 4029
rect 2596 3952 2648 4004
rect 15476 4020 15528 4072
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 6736 3952 6788 4004
rect 13544 3952 13596 4004
rect 17960 4020 18012 4072
rect 18236 4020 18288 4072
rect 18420 4156 18472 4208
rect 23388 4267 23440 4276
rect 23388 4233 23397 4267
rect 23397 4233 23431 4267
rect 23431 4233 23440 4267
rect 23388 4224 23440 4233
rect 25412 4224 25464 4276
rect 30012 4224 30064 4276
rect 31668 4224 31720 4276
rect 18788 4131 18840 4140
rect 18788 4097 18797 4131
rect 18797 4097 18831 4131
rect 18831 4097 18840 4131
rect 18788 4088 18840 4097
rect 20260 4088 20312 4140
rect 20904 4131 20956 4140
rect 20904 4097 20913 4131
rect 20913 4097 20947 4131
rect 20947 4097 20956 4131
rect 20904 4088 20956 4097
rect 21548 4088 21600 4140
rect 21824 4088 21876 4140
rect 27620 4088 27672 4140
rect 30472 4156 30524 4208
rect 18696 4020 18748 4072
rect 33048 4088 33100 4140
rect 17868 3952 17920 4004
rect 19524 3952 19576 4004
rect 20352 3952 20404 4004
rect 21180 3995 21232 4004
rect 21180 3961 21189 3995
rect 21189 3961 21223 3995
rect 21223 3961 21232 3995
rect 21180 3952 21232 3961
rect 11704 3884 11756 3936
rect 15384 3884 15436 3936
rect 15568 3927 15620 3936
rect 15568 3893 15577 3927
rect 15577 3893 15611 3927
rect 15611 3893 15620 3927
rect 15568 3884 15620 3893
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16948 3884 17000 3936
rect 21824 3884 21876 3936
rect 22192 3884 22244 3936
rect 23480 3884 23532 3936
rect 23572 3927 23624 3936
rect 23572 3893 23581 3927
rect 23581 3893 23615 3927
rect 23615 3893 23624 3927
rect 23572 3884 23624 3893
rect 28264 3952 28316 4004
rect 28172 3884 28224 3936
rect 33508 3952 33560 4004
rect 31300 3884 31352 3936
rect 6946 3782 6998 3834
rect 7010 3782 7062 3834
rect 7074 3782 7126 3834
rect 7138 3782 7190 3834
rect 7202 3782 7254 3834
rect 14306 3782 14358 3834
rect 14370 3782 14422 3834
rect 14434 3782 14486 3834
rect 14498 3782 14550 3834
rect 14562 3782 14614 3834
rect 21666 3782 21718 3834
rect 21730 3782 21782 3834
rect 21794 3782 21846 3834
rect 21858 3782 21910 3834
rect 21922 3782 21974 3834
rect 29026 3782 29078 3834
rect 29090 3782 29142 3834
rect 29154 3782 29206 3834
rect 29218 3782 29270 3834
rect 29282 3782 29334 3834
rect 3516 3680 3568 3732
rect 13360 3680 13412 3732
rect 13544 3680 13596 3732
rect 14004 3680 14056 3732
rect 6828 3612 6880 3664
rect 16028 3680 16080 3732
rect 16580 3680 16632 3732
rect 17592 3680 17644 3732
rect 17868 3680 17920 3732
rect 19432 3680 19484 3732
rect 4252 3587 4304 3596
rect 4252 3553 4261 3587
rect 4261 3553 4295 3587
rect 4295 3553 4304 3587
rect 4252 3544 4304 3553
rect 5724 3544 5776 3596
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 12624 3544 12676 3596
rect 13636 3544 13688 3596
rect 1308 3476 1360 3528
rect 4528 3476 4580 3528
rect 10324 3476 10376 3528
rect 15844 3612 15896 3664
rect 19800 3612 19852 3664
rect 20444 3680 20496 3732
rect 21180 3680 21232 3732
rect 22192 3680 22244 3732
rect 23112 3723 23164 3732
rect 23112 3689 23121 3723
rect 23121 3689 23155 3723
rect 23155 3689 23164 3723
rect 23112 3680 23164 3689
rect 23388 3680 23440 3732
rect 15476 3544 15528 3596
rect 16120 3544 16172 3596
rect 17040 3544 17092 3596
rect 20904 3544 20956 3596
rect 16948 3476 17000 3528
rect 20260 3476 20312 3528
rect 20720 3408 20772 3460
rect 23480 3476 23532 3528
rect 24032 3680 24084 3732
rect 31668 3612 31720 3664
rect 25780 3587 25832 3596
rect 25780 3553 25789 3587
rect 25789 3553 25823 3587
rect 25823 3553 25832 3587
rect 25780 3544 25832 3553
rect 30012 3544 30064 3596
rect 24492 3476 24544 3528
rect 20628 3340 20680 3392
rect 30288 3476 30340 3528
rect 6286 3238 6338 3290
rect 6350 3238 6402 3290
rect 6414 3238 6466 3290
rect 6478 3238 6530 3290
rect 6542 3238 6594 3290
rect 13646 3238 13698 3290
rect 13710 3238 13762 3290
rect 13774 3238 13826 3290
rect 13838 3238 13890 3290
rect 13902 3238 13954 3290
rect 21006 3238 21058 3290
rect 21070 3238 21122 3290
rect 21134 3238 21186 3290
rect 21198 3238 21250 3290
rect 21262 3238 21314 3290
rect 28366 3238 28418 3290
rect 28430 3238 28482 3290
rect 28494 3238 28546 3290
rect 28558 3238 28610 3290
rect 28622 3238 28674 3290
rect 14188 3136 14240 3188
rect 14832 3136 14884 3188
rect 15016 3136 15068 3188
rect 15568 3068 15620 3120
rect 20904 3136 20956 3188
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 16396 3000 16448 3052
rect 18052 3000 18104 3052
rect 18236 3000 18288 3052
rect 19064 3043 19116 3052
rect 19064 3009 19073 3043
rect 19073 3009 19107 3043
rect 19107 3009 19116 3043
rect 19064 3000 19116 3009
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 20 2864 72 2916
rect 3608 2864 3660 2916
rect 7656 2932 7708 2984
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 5816 2864 5868 2916
rect 7288 2864 7340 2916
rect 9036 2864 9088 2916
rect 11520 2932 11572 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 15384 2932 15436 2984
rect 16304 2932 16356 2984
rect 17960 2975 18012 2984
rect 17960 2941 17969 2975
rect 17969 2941 18003 2975
rect 18003 2941 18012 2975
rect 17960 2932 18012 2941
rect 19432 3000 19484 3052
rect 22560 3000 22612 3052
rect 25780 3000 25832 3052
rect 21272 2932 21324 2984
rect 23480 2975 23532 2984
rect 23480 2941 23489 2975
rect 23489 2941 23523 2975
rect 23523 2941 23532 2975
rect 23480 2932 23532 2941
rect 23572 2932 23624 2984
rect 18144 2864 18196 2916
rect 18328 2864 18380 2916
rect 30932 3136 30984 3188
rect 31852 3136 31904 3188
rect 27068 2932 27120 2984
rect 29368 2932 29420 2984
rect 32220 3000 32272 3052
rect 18696 2796 18748 2848
rect 19708 2796 19760 2848
rect 33140 2864 33192 2916
rect 34796 2796 34848 2848
rect 6946 2694 6998 2746
rect 7010 2694 7062 2746
rect 7074 2694 7126 2746
rect 7138 2694 7190 2746
rect 7202 2694 7254 2746
rect 14306 2694 14358 2746
rect 14370 2694 14422 2746
rect 14434 2694 14486 2746
rect 14498 2694 14550 2746
rect 14562 2694 14614 2746
rect 21666 2694 21718 2746
rect 21730 2694 21782 2746
rect 21794 2694 21846 2746
rect 21858 2694 21910 2746
rect 21922 2694 21974 2746
rect 29026 2694 29078 2746
rect 29090 2694 29142 2746
rect 29154 2694 29206 2746
rect 29218 2694 29270 2746
rect 29282 2694 29334 2746
<< metal2 >>
rect 662 33674 718 34344
rect 1950 33674 2006 34344
rect 3882 33674 3938 34344
rect 4526 34096 4582 34105
rect 4526 34031 4582 34040
rect 662 33646 1072 33674
rect 662 33544 718 33646
rect 1044 31958 1072 33646
rect 1950 33646 2360 33674
rect 1950 33544 2006 33646
rect 1032 31952 1084 31958
rect 1032 31894 1084 31900
rect 2332 31346 2360 33646
rect 3882 33646 4200 33674
rect 3882 33544 3938 33646
rect 2778 32056 2834 32065
rect 2778 31991 2834 32000
rect 2320 31340 2372 31346
rect 2320 31282 2372 31288
rect 1308 30728 1360 30734
rect 1306 30696 1308 30705
rect 1360 30696 1362 30705
rect 1306 30631 1362 30640
rect 2792 30258 2820 31991
rect 4172 31958 4200 33646
rect 4160 31952 4212 31958
rect 4160 31894 4212 31900
rect 3884 31884 3936 31890
rect 3884 31826 3936 31832
rect 2780 30252 2832 30258
rect 2780 30194 2832 30200
rect 3148 29708 3200 29714
rect 3148 29650 3200 29656
rect 1308 27464 1360 27470
rect 1308 27406 1360 27412
rect 1320 27305 1348 27406
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 1308 24812 1360 24818
rect 1308 24754 1360 24760
rect 1320 23905 1348 24754
rect 1306 23896 1362 23905
rect 1306 23831 1362 23840
rect 1306 22536 1362 22545
rect 1306 22471 1308 22480
rect 1360 22471 1362 22480
rect 1308 22442 1360 22448
rect 3160 22094 3188 29650
rect 3516 29640 3568 29646
rect 3516 29582 3568 29588
rect 3528 28665 3556 29582
rect 3896 29306 3924 31826
rect 4160 31272 4212 31278
rect 4160 31214 4212 31220
rect 3884 29300 3936 29306
rect 3884 29242 3936 29248
rect 3514 28656 3570 28665
rect 3514 28591 3570 28600
rect 3896 28082 3924 29242
rect 3884 28076 3936 28082
rect 3884 28018 3936 28024
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3252 25945 3280 26318
rect 3238 25936 3294 25945
rect 3238 25871 3294 25880
rect 3424 25288 3476 25294
rect 3424 25230 3476 25236
rect 3240 24744 3292 24750
rect 3240 24686 3292 24692
rect 3252 24274 3280 24686
rect 3436 24410 3464 25230
rect 3884 24676 3936 24682
rect 3884 24618 3936 24624
rect 3896 24410 3924 24618
rect 3424 24404 3476 24410
rect 3424 24346 3476 24352
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 3240 24268 3292 24274
rect 3240 24210 3292 24216
rect 3252 23866 3280 24210
rect 4172 23866 4200 31214
rect 4540 30802 4568 34031
rect 5170 33544 5226 34344
rect 6458 33544 6514 34344
rect 8390 33674 8446 34344
rect 8390 33646 8708 33674
rect 8390 33544 8446 33646
rect 5184 31958 5212 33544
rect 6472 31958 6500 33544
rect 6946 32124 7254 32133
rect 6946 32122 6952 32124
rect 7008 32122 7032 32124
rect 7088 32122 7112 32124
rect 7168 32122 7192 32124
rect 7248 32122 7254 32124
rect 7008 32070 7010 32122
rect 7190 32070 7192 32122
rect 6946 32068 6952 32070
rect 7008 32068 7032 32070
rect 7088 32068 7112 32070
rect 7168 32068 7192 32070
rect 7248 32068 7254 32070
rect 6946 32059 7254 32068
rect 7564 32020 7616 32026
rect 7564 31962 7616 31968
rect 5172 31952 5224 31958
rect 5172 31894 5224 31900
rect 6460 31952 6512 31958
rect 6460 31894 6512 31900
rect 6644 31884 6696 31890
rect 6644 31826 6696 31832
rect 6286 31580 6594 31589
rect 6286 31578 6292 31580
rect 6348 31578 6372 31580
rect 6428 31578 6452 31580
rect 6508 31578 6532 31580
rect 6588 31578 6594 31580
rect 6348 31526 6350 31578
rect 6530 31526 6532 31578
rect 6286 31524 6292 31526
rect 6348 31524 6372 31526
rect 6428 31524 6452 31526
rect 6508 31524 6532 31526
rect 6588 31524 6594 31526
rect 6286 31515 6594 31524
rect 4436 30796 4488 30802
rect 4436 30738 4488 30744
rect 4528 30796 4580 30802
rect 4528 30738 4580 30744
rect 4448 29850 4476 30738
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 4528 30184 4580 30190
rect 4528 30126 4580 30132
rect 4436 29844 4488 29850
rect 4436 29786 4488 29792
rect 4252 28960 4304 28966
rect 4252 28902 4304 28908
rect 4264 28422 4292 28902
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4264 25906 4292 28358
rect 4540 26450 4568 30126
rect 4988 29028 5040 29034
rect 4988 28970 5040 28976
rect 5000 28218 5028 28970
rect 5264 28688 5316 28694
rect 5264 28630 5316 28636
rect 4988 28212 5040 28218
rect 4988 28154 5040 28160
rect 5276 27674 5304 28630
rect 5264 27668 5316 27674
rect 5264 27610 5316 27616
rect 4528 26444 4580 26450
rect 4528 26386 4580 26392
rect 4540 26042 4568 26386
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 4528 26036 4580 26042
rect 4528 25978 4580 25984
rect 4252 25900 4304 25906
rect 4252 25842 4304 25848
rect 4264 24818 4292 25842
rect 4988 25764 5040 25770
rect 4988 25706 5040 25712
rect 5000 25498 5028 25706
rect 5184 25498 5212 26182
rect 5264 25696 5316 25702
rect 5264 25638 5316 25644
rect 5276 25498 5304 25638
rect 4988 25492 5040 25498
rect 4988 25434 5040 25440
rect 5172 25492 5224 25498
rect 5172 25434 5224 25440
rect 5264 25492 5316 25498
rect 5264 25434 5316 25440
rect 4528 25152 4580 25158
rect 4528 25094 4580 25100
rect 4252 24812 4304 24818
rect 4252 24754 4304 24760
rect 4264 24274 4292 24754
rect 4252 24268 4304 24274
rect 4252 24210 4304 24216
rect 4252 24132 4304 24138
rect 4252 24074 4304 24080
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 4160 23860 4212 23866
rect 4160 23802 4212 23808
rect 4172 23322 4200 23802
rect 4264 23338 4292 24074
rect 4540 23730 4568 25094
rect 4620 24608 4672 24614
rect 4620 24550 4672 24556
rect 5264 24608 5316 24614
rect 5264 24550 5316 24556
rect 4632 24410 4660 24550
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4528 23724 4580 23730
rect 4528 23666 4580 23672
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 4264 23322 4476 23338
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 4264 23316 4488 23322
rect 4264 23310 4436 23316
rect 3160 22066 3280 22094
rect 3252 22030 3280 22066
rect 3240 22024 3292 22030
rect 3240 21966 3292 21972
rect 3252 21690 3280 21966
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 3240 21684 3292 21690
rect 3240 21626 3292 21632
rect 4172 21146 4200 21830
rect 4160 21140 4212 21146
rect 4160 21082 4212 21088
rect 3330 21040 3386 21049
rect 3330 20975 3332 20984
rect 3384 20975 3386 20984
rect 3332 20946 3384 20952
rect 4264 20942 4292 23310
rect 4436 23258 4488 23264
rect 4988 23248 5040 23254
rect 4988 23190 5040 23196
rect 5000 22778 5028 23190
rect 4988 22772 5040 22778
rect 4988 22714 5040 22720
rect 5184 22574 5212 23462
rect 5276 23322 5304 24550
rect 5264 23316 5316 23322
rect 5264 23258 5316 23264
rect 5172 22568 5224 22574
rect 5172 22510 5224 22516
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4632 21146 4660 21354
rect 4712 21344 4764 21350
rect 4712 21286 4764 21292
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 3068 20505 3096 20878
rect 4264 20602 4292 20878
rect 4252 20596 4304 20602
rect 4252 20538 4304 20544
rect 3054 20496 3110 20505
rect 3054 20431 3110 20440
rect 4724 19854 4752 21286
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 5276 19990 5304 20742
rect 5264 19984 5316 19990
rect 5264 19926 5316 19932
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 1308 19304 1360 19310
rect 1308 19246 1360 19252
rect 1320 19145 1348 19246
rect 3240 19168 3292 19174
rect 1306 19136 1362 19145
rect 3240 19110 3292 19116
rect 1306 19071 1362 19080
rect 1308 15972 1360 15978
rect 1308 15914 1360 15920
rect 1320 15745 1348 15914
rect 1306 15736 1362 15745
rect 1306 15671 1362 15680
rect 1306 14376 1362 14385
rect 1306 14311 1362 14320
rect 1320 13938 1348 14311
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1320 13025 1348 13262
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 3252 12434 3280 19110
rect 4724 18766 4752 19790
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5000 18426 5028 18702
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 5184 18358 5212 18566
rect 5172 18352 5224 18358
rect 5172 18294 5224 18300
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4080 17785 4108 18090
rect 4066 17776 4122 17785
rect 4066 17711 4122 17720
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 3424 15904 3476 15910
rect 3424 15846 3476 15852
rect 3436 15706 3464 15846
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 5276 15638 5304 16390
rect 5264 15632 5316 15638
rect 5264 15574 5316 15580
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4264 14278 4292 14758
rect 4448 14414 4476 14758
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4252 14272 4304 14278
rect 4252 14214 4304 14220
rect 4264 13870 4292 14214
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 3252 12406 3372 12434
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3252 10985 3280 11086
rect 3238 10976 3294 10985
rect 3238 10911 3294 10920
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 3068 9625 3096 10066
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3054 9616 3110 9625
rect 3054 9551 3110 9560
rect 3252 8090 3280 9862
rect 3344 8634 3372 12406
rect 4344 12368 4396 12374
rect 4344 12310 4396 12316
rect 4356 11898 4384 12310
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11898 4752 12038
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4436 11552 4488 11558
rect 4436 11494 4488 11500
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 4448 11218 4476 11494
rect 5276 11286 5304 11494
rect 5264 11280 5316 11286
rect 5264 11222 5316 11228
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4344 10600 4396 10606
rect 4344 10542 4396 10548
rect 4356 9926 4384 10542
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 1308 7948 1360 7954
rect 1308 7890 1360 7896
rect 1320 7585 1348 7890
rect 4264 7750 4292 8230
rect 4252 7744 4304 7750
rect 4252 7686 4304 7692
rect 1306 7576 1362 7585
rect 1306 7511 1362 7520
rect 1308 6248 1360 6254
rect 1306 6216 1308 6225
rect 1360 6216 1362 6225
rect 1306 6151 1362 6160
rect 1308 5092 1360 5098
rect 1308 5034 1360 5040
rect 1320 4865 1348 5034
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 2596 4004 2648 4010
rect 2596 3946 2648 3952
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 20 2916 72 2922
rect 20 2858 72 2864
rect 32 800 60 2858
rect 1320 800 1348 3470
rect 2608 800 2636 3946
rect 3068 1465 3096 4014
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3528 3738 3556 3878
rect 3516 3732 3568 3738
rect 3516 3674 3568 3680
rect 4264 3602 4292 7686
rect 4356 5166 4384 9862
rect 5368 6254 5396 30670
rect 6286 30492 6594 30501
rect 6286 30490 6292 30492
rect 6348 30490 6372 30492
rect 6428 30490 6452 30492
rect 6508 30490 6532 30492
rect 6588 30490 6594 30492
rect 6348 30438 6350 30490
rect 6530 30438 6532 30490
rect 6286 30436 6292 30438
rect 6348 30436 6372 30438
rect 6428 30436 6452 30438
rect 6508 30436 6532 30438
rect 6588 30436 6594 30438
rect 6286 30427 6594 30436
rect 6286 29404 6594 29413
rect 6286 29402 6292 29404
rect 6348 29402 6372 29404
rect 6428 29402 6452 29404
rect 6508 29402 6532 29404
rect 6588 29402 6594 29404
rect 6348 29350 6350 29402
rect 6530 29350 6532 29402
rect 6286 29348 6292 29350
rect 6348 29348 6372 29350
rect 6428 29348 6452 29350
rect 6508 29348 6532 29350
rect 6588 29348 6594 29350
rect 6286 29339 6594 29348
rect 6184 29028 6236 29034
rect 6184 28970 6236 28976
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5460 28218 5488 28494
rect 5816 28416 5868 28422
rect 5816 28358 5868 28364
rect 5828 28218 5856 28358
rect 5448 28212 5500 28218
rect 5448 28154 5500 28160
rect 5816 28212 5868 28218
rect 5816 28154 5868 28160
rect 5540 27940 5592 27946
rect 5540 27882 5592 27888
rect 5552 27334 5580 27882
rect 6196 27538 6224 28970
rect 6656 28626 6684 31826
rect 6946 31036 7254 31045
rect 6946 31034 6952 31036
rect 7008 31034 7032 31036
rect 7088 31034 7112 31036
rect 7168 31034 7192 31036
rect 7248 31034 7254 31036
rect 7008 30982 7010 31034
rect 7190 30982 7192 31034
rect 6946 30980 6952 30982
rect 7008 30980 7032 30982
rect 7088 30980 7112 30982
rect 7168 30980 7192 30982
rect 7248 30980 7254 30982
rect 6946 30971 7254 30980
rect 6946 29948 7254 29957
rect 6946 29946 6952 29948
rect 7008 29946 7032 29948
rect 7088 29946 7112 29948
rect 7168 29946 7192 29948
rect 7248 29946 7254 29948
rect 7008 29894 7010 29946
rect 7190 29894 7192 29946
rect 6946 29892 6952 29894
rect 7008 29892 7032 29894
rect 7088 29892 7112 29894
rect 7168 29892 7192 29894
rect 7248 29892 7254 29894
rect 6946 29883 7254 29892
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 6828 28960 6880 28966
rect 6828 28902 6880 28908
rect 6644 28620 6696 28626
rect 6644 28562 6696 28568
rect 6644 28484 6696 28490
rect 6644 28426 6696 28432
rect 6286 28316 6594 28325
rect 6286 28314 6292 28316
rect 6348 28314 6372 28316
rect 6428 28314 6452 28316
rect 6508 28314 6532 28316
rect 6588 28314 6594 28316
rect 6348 28262 6350 28314
rect 6530 28262 6532 28314
rect 6286 28260 6292 28262
rect 6348 28260 6372 28262
rect 6428 28260 6452 28262
rect 6508 28260 6532 28262
rect 6588 28260 6594 28262
rect 6286 28251 6594 28260
rect 6552 27872 6604 27878
rect 6552 27814 6604 27820
rect 6564 27606 6592 27814
rect 6656 27674 6684 28426
rect 6840 27946 6868 28902
rect 6946 28860 7254 28869
rect 6946 28858 6952 28860
rect 7008 28858 7032 28860
rect 7088 28858 7112 28860
rect 7168 28858 7192 28860
rect 7248 28858 7254 28860
rect 7008 28806 7010 28858
rect 7190 28806 7192 28858
rect 6946 28804 6952 28806
rect 7008 28804 7032 28806
rect 7088 28804 7112 28806
rect 7168 28804 7192 28806
rect 7248 28804 7254 28806
rect 6946 28795 7254 28804
rect 6828 27940 6880 27946
rect 6828 27882 6880 27888
rect 7392 27878 7420 29582
rect 7288 27872 7340 27878
rect 7288 27814 7340 27820
rect 7380 27872 7432 27878
rect 7380 27814 7432 27820
rect 6946 27772 7254 27781
rect 6946 27770 6952 27772
rect 7008 27770 7032 27772
rect 7088 27770 7112 27772
rect 7168 27770 7192 27772
rect 7248 27770 7254 27772
rect 7008 27718 7010 27770
rect 7190 27718 7192 27770
rect 6946 27716 6952 27718
rect 7008 27716 7032 27718
rect 7088 27716 7112 27718
rect 7168 27716 7192 27718
rect 7248 27716 7254 27718
rect 6946 27707 7254 27716
rect 7300 27674 7328 27814
rect 6644 27668 6696 27674
rect 6644 27610 6696 27616
rect 7288 27668 7340 27674
rect 7288 27610 7340 27616
rect 6552 27600 6604 27606
rect 6920 27600 6972 27606
rect 6552 27542 6604 27548
rect 6826 27568 6882 27577
rect 6184 27532 6236 27538
rect 7196 27600 7248 27606
rect 6972 27560 7196 27588
rect 6920 27542 6972 27548
rect 7196 27542 7248 27548
rect 6826 27503 6828 27512
rect 6184 27474 6236 27480
rect 6880 27503 6882 27512
rect 6828 27474 6880 27480
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 5552 26234 5580 27270
rect 6196 26926 6224 27474
rect 6828 27396 6880 27402
rect 6828 27338 6880 27344
rect 6644 27328 6696 27334
rect 6840 27282 6868 27338
rect 6696 27276 6868 27282
rect 6644 27270 6868 27276
rect 6656 27254 6868 27270
rect 6286 27228 6594 27237
rect 6286 27226 6292 27228
rect 6348 27226 6372 27228
rect 6428 27226 6452 27228
rect 6508 27226 6532 27228
rect 6588 27226 6594 27228
rect 6348 27174 6350 27226
rect 6530 27174 6532 27226
rect 6286 27172 6292 27174
rect 6348 27172 6372 27174
rect 6428 27172 6452 27174
rect 6508 27172 6532 27174
rect 6588 27172 6594 27174
rect 6286 27163 6594 27172
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6644 26784 6696 26790
rect 6644 26726 6696 26732
rect 6656 26518 6684 26726
rect 6840 26586 6868 27254
rect 6946 26684 7254 26693
rect 6946 26682 6952 26684
rect 7008 26682 7032 26684
rect 7088 26682 7112 26684
rect 7168 26682 7192 26684
rect 7248 26682 7254 26684
rect 7008 26630 7010 26682
rect 7190 26630 7192 26682
rect 6946 26628 6952 26630
rect 7008 26628 7032 26630
rect 7088 26628 7112 26630
rect 7168 26628 7192 26630
rect 7248 26628 7254 26630
rect 6946 26619 7254 26628
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6644 26512 6696 26518
rect 6644 26454 6696 26460
rect 5816 26444 5868 26450
rect 5816 26386 5868 26392
rect 5460 26206 5580 26234
rect 5460 24614 5488 26206
rect 5828 25906 5856 26386
rect 7392 26382 7420 27814
rect 7380 26376 7432 26382
rect 7380 26318 7432 26324
rect 6286 26140 6594 26149
rect 6286 26138 6292 26140
rect 6348 26138 6372 26140
rect 6428 26138 6452 26140
rect 6508 26138 6532 26140
rect 6588 26138 6594 26140
rect 6348 26086 6350 26138
rect 6530 26086 6532 26138
rect 6286 26084 6292 26086
rect 6348 26084 6372 26086
rect 6428 26084 6452 26086
rect 6508 26084 6532 26086
rect 6588 26084 6594 26086
rect 6286 26075 6594 26084
rect 5816 25900 5868 25906
rect 5816 25842 5868 25848
rect 5632 25696 5684 25702
rect 5632 25638 5684 25644
rect 6184 25696 6236 25702
rect 6184 25638 6236 25644
rect 7288 25696 7340 25702
rect 7288 25638 7340 25644
rect 5644 25158 5672 25638
rect 6196 25430 6224 25638
rect 6946 25596 7254 25605
rect 6946 25594 6952 25596
rect 7008 25594 7032 25596
rect 7088 25594 7112 25596
rect 7168 25594 7192 25596
rect 7248 25594 7254 25596
rect 7008 25542 7010 25594
rect 7190 25542 7192 25594
rect 6946 25540 6952 25542
rect 7008 25540 7032 25542
rect 7088 25540 7112 25542
rect 7168 25540 7192 25542
rect 7248 25540 7254 25542
rect 6946 25531 7254 25540
rect 5816 25424 5868 25430
rect 5816 25366 5868 25372
rect 6184 25424 6236 25430
rect 6184 25366 6236 25372
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5552 24750 5580 25094
rect 5644 24834 5672 25094
rect 5828 24954 5856 25366
rect 7300 25362 7328 25638
rect 6276 25356 6328 25362
rect 6276 25298 6328 25304
rect 7288 25356 7340 25362
rect 7288 25298 7340 25304
rect 5908 25288 5960 25294
rect 6288 25242 6316 25298
rect 5908 25230 5960 25236
rect 5816 24948 5868 24954
rect 5816 24890 5868 24896
rect 5920 24834 5948 25230
rect 5644 24806 5948 24834
rect 5540 24744 5592 24750
rect 5540 24686 5592 24692
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5644 24274 5672 24550
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 5920 24070 5948 24806
rect 6196 25214 6316 25242
rect 6196 24750 6224 25214
rect 6286 25052 6594 25061
rect 6286 25050 6292 25052
rect 6348 25050 6372 25052
rect 6428 25050 6452 25052
rect 6508 25050 6532 25052
rect 6588 25050 6594 25052
rect 6348 24998 6350 25050
rect 6530 24998 6532 25050
rect 6286 24996 6292 24998
rect 6348 24996 6372 24998
rect 6428 24996 6452 24998
rect 6508 24996 6532 24998
rect 6588 24996 6594 24998
rect 6286 24987 6594 24996
rect 7392 24818 7420 26318
rect 7472 25356 7524 25362
rect 7472 25298 7524 25304
rect 7380 24812 7432 24818
rect 7380 24754 7432 24760
rect 6184 24744 6236 24750
rect 6184 24686 6236 24692
rect 6460 24744 6512 24750
rect 6460 24686 6512 24692
rect 7288 24744 7340 24750
rect 7484 24698 7512 25298
rect 7288 24686 7340 24692
rect 6472 24410 6500 24686
rect 6946 24508 7254 24517
rect 6946 24506 6952 24508
rect 7008 24506 7032 24508
rect 7088 24506 7112 24508
rect 7168 24506 7192 24508
rect 7248 24506 7254 24508
rect 7008 24454 7010 24506
rect 7190 24454 7192 24506
rect 6946 24452 6952 24454
rect 7008 24452 7032 24454
rect 7088 24452 7112 24454
rect 7168 24452 7192 24454
rect 7248 24452 7254 24454
rect 6946 24443 7254 24452
rect 7300 24410 7328 24686
rect 7392 24670 7512 24698
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 7288 24404 7340 24410
rect 7288 24346 7340 24352
rect 5908 24064 5960 24070
rect 5908 24006 5960 24012
rect 5724 23724 5776 23730
rect 5724 23666 5776 23672
rect 5540 23520 5592 23526
rect 5540 23462 5592 23468
rect 5552 23254 5580 23462
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5736 23186 5764 23666
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5448 22432 5500 22438
rect 5448 22374 5500 22380
rect 5460 22234 5488 22374
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5644 18290 5672 22918
rect 5736 22778 5764 23122
rect 5920 23118 5948 24006
rect 6286 23964 6594 23973
rect 6286 23962 6292 23964
rect 6348 23962 6372 23964
rect 6428 23962 6452 23964
rect 6508 23962 6532 23964
rect 6588 23962 6594 23964
rect 6348 23910 6350 23962
rect 6530 23910 6532 23962
rect 6286 23908 6292 23910
rect 6348 23908 6372 23910
rect 6428 23908 6452 23910
rect 6508 23908 6532 23910
rect 6588 23908 6594 23910
rect 6286 23899 6594 23908
rect 6552 23656 6604 23662
rect 6552 23598 6604 23604
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 6472 23322 6500 23462
rect 6564 23322 6592 23598
rect 6946 23420 7254 23429
rect 6946 23418 6952 23420
rect 7008 23418 7032 23420
rect 7088 23418 7112 23420
rect 7168 23418 7192 23420
rect 7248 23418 7254 23420
rect 7008 23366 7010 23418
rect 7190 23366 7192 23418
rect 6946 23364 6952 23366
rect 7008 23364 7032 23366
rect 7088 23364 7112 23366
rect 7168 23364 7192 23366
rect 7248 23364 7254 23366
rect 6946 23355 7254 23364
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 6552 23316 6604 23322
rect 6552 23258 6604 23264
rect 7104 23248 7156 23254
rect 7104 23190 7156 23196
rect 5908 23112 5960 23118
rect 5908 23054 5960 23060
rect 6736 23112 6788 23118
rect 6736 23054 6788 23060
rect 6286 22876 6594 22885
rect 6286 22874 6292 22876
rect 6348 22874 6372 22876
rect 6428 22874 6452 22876
rect 6508 22874 6532 22876
rect 6588 22874 6594 22876
rect 6348 22822 6350 22874
rect 6530 22822 6532 22874
rect 6286 22820 6292 22822
rect 6348 22820 6372 22822
rect 6428 22820 6452 22822
rect 6508 22820 6532 22822
rect 6588 22820 6594 22822
rect 6286 22811 6594 22820
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5736 22094 5764 22714
rect 6092 22568 6144 22574
rect 6144 22528 6224 22556
rect 6092 22510 6144 22516
rect 5736 22066 6132 22094
rect 6104 22030 6132 22066
rect 6092 22024 6144 22030
rect 6092 21966 6144 21972
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 6012 21554 6040 21830
rect 6000 21548 6052 21554
rect 6000 21490 6052 21496
rect 5724 21344 5776 21350
rect 5724 21286 5776 21292
rect 5736 19990 5764 21286
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5828 20602 5856 20878
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 5724 19848 5776 19854
rect 5828 19802 5856 20402
rect 5920 20398 5948 20946
rect 6104 20466 6132 21966
rect 6196 21690 6224 22528
rect 6644 22500 6696 22506
rect 6644 22442 6696 22448
rect 6276 22432 6328 22438
rect 6276 22374 6328 22380
rect 6552 22432 6604 22438
rect 6552 22374 6604 22380
rect 6288 22234 6316 22374
rect 6564 22234 6592 22374
rect 6656 22234 6684 22442
rect 6276 22228 6328 22234
rect 6276 22170 6328 22176
rect 6552 22228 6604 22234
rect 6552 22170 6604 22176
rect 6644 22228 6696 22234
rect 6644 22170 6696 22176
rect 6460 22024 6512 22030
rect 6512 21972 6684 21978
rect 6460 21966 6684 21972
rect 6472 21950 6684 21966
rect 6286 21788 6594 21797
rect 6286 21786 6292 21788
rect 6348 21786 6372 21788
rect 6428 21786 6452 21788
rect 6508 21786 6532 21788
rect 6588 21786 6594 21788
rect 6348 21734 6350 21786
rect 6530 21734 6532 21786
rect 6286 21732 6292 21734
rect 6348 21732 6372 21734
rect 6428 21732 6452 21734
rect 6508 21732 6532 21734
rect 6588 21732 6594 21734
rect 6286 21723 6594 21732
rect 6184 21684 6236 21690
rect 6184 21626 6236 21632
rect 6286 20700 6594 20709
rect 6286 20698 6292 20700
rect 6348 20698 6372 20700
rect 6428 20698 6452 20700
rect 6508 20698 6532 20700
rect 6588 20698 6594 20700
rect 6348 20646 6350 20698
rect 6530 20646 6532 20698
rect 6286 20644 6292 20646
rect 6348 20644 6372 20646
rect 6428 20644 6452 20646
rect 6508 20644 6532 20646
rect 6588 20644 6594 20646
rect 6286 20635 6594 20644
rect 6092 20460 6144 20466
rect 6092 20402 6144 20408
rect 5908 20392 5960 20398
rect 5908 20334 5960 20340
rect 6368 20324 6420 20330
rect 6368 20266 6420 20272
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5776 19796 5856 19802
rect 5724 19790 5856 19796
rect 5736 19774 5856 19790
rect 6012 19786 6040 20198
rect 6380 20058 6408 20266
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6000 19780 6052 19786
rect 6000 19722 6052 19728
rect 6286 19612 6594 19621
rect 6286 19610 6292 19612
rect 6348 19610 6372 19612
rect 6428 19610 6452 19612
rect 6508 19610 6532 19612
rect 6588 19610 6594 19612
rect 6348 19558 6350 19610
rect 6530 19558 6532 19610
rect 6286 19556 6292 19558
rect 6348 19556 6372 19558
rect 6428 19556 6452 19558
rect 6508 19556 6532 19558
rect 6588 19556 6594 19558
rect 6286 19547 6594 19556
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6000 18624 6052 18630
rect 6000 18566 6052 18572
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5908 16652 5960 16658
rect 5908 16594 5960 16600
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15706 5488 15846
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5460 14414 5488 15438
rect 5644 15026 5672 16050
rect 5816 15972 5868 15978
rect 5816 15914 5868 15920
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15026 5764 15302
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5460 13938 5488 14350
rect 5644 14074 5672 14962
rect 5828 14958 5856 15914
rect 5920 15162 5948 16594
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5816 14952 5868 14958
rect 5816 14894 5868 14900
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 6012 13394 6040 18566
rect 6104 18426 6132 18770
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6092 18284 6144 18290
rect 6092 18226 6144 18232
rect 6104 14958 6132 18226
rect 6196 18222 6224 18634
rect 6286 18524 6594 18533
rect 6286 18522 6292 18524
rect 6348 18522 6372 18524
rect 6428 18522 6452 18524
rect 6508 18522 6532 18524
rect 6588 18522 6594 18524
rect 6348 18470 6350 18522
rect 6530 18470 6532 18522
rect 6286 18468 6292 18470
rect 6348 18468 6372 18470
rect 6428 18468 6452 18470
rect 6508 18468 6532 18470
rect 6588 18468 6594 18470
rect 6286 18459 6594 18468
rect 6460 18420 6512 18426
rect 6460 18362 6512 18368
rect 6472 18306 6500 18362
rect 6380 18290 6500 18306
rect 6368 18284 6500 18290
rect 6420 18278 6500 18284
rect 6368 18226 6420 18232
rect 6184 18216 6236 18222
rect 6184 18158 6236 18164
rect 6286 17436 6594 17445
rect 6286 17434 6292 17436
rect 6348 17434 6372 17436
rect 6428 17434 6452 17436
rect 6508 17434 6532 17436
rect 6588 17434 6594 17436
rect 6348 17382 6350 17434
rect 6530 17382 6532 17434
rect 6286 17380 6292 17382
rect 6348 17380 6372 17382
rect 6428 17380 6452 17382
rect 6508 17380 6532 17382
rect 6588 17380 6594 17382
rect 6286 17371 6594 17380
rect 6286 16348 6594 16357
rect 6286 16346 6292 16348
rect 6348 16346 6372 16348
rect 6428 16346 6452 16348
rect 6508 16346 6532 16348
rect 6588 16346 6594 16348
rect 6348 16294 6350 16346
rect 6530 16294 6532 16346
rect 6286 16292 6292 16294
rect 6348 16292 6372 16294
rect 6428 16292 6452 16294
rect 6508 16292 6532 16294
rect 6588 16292 6594 16294
rect 6286 16283 6594 16292
rect 6656 16114 6684 21950
rect 6748 21554 6776 23054
rect 7116 22642 7144 23190
rect 7196 22976 7248 22982
rect 7196 22918 7248 22924
rect 7208 22778 7236 22918
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 6828 22432 6880 22438
rect 6828 22374 6880 22380
rect 6840 21622 6868 22374
rect 6946 22332 7254 22341
rect 6946 22330 6952 22332
rect 7008 22330 7032 22332
rect 7088 22330 7112 22332
rect 7168 22330 7192 22332
rect 7248 22330 7254 22332
rect 7008 22278 7010 22330
rect 7190 22278 7192 22330
rect 6946 22276 6952 22278
rect 7008 22276 7032 22278
rect 7088 22276 7112 22278
rect 7168 22276 7192 22278
rect 7248 22276 7254 22278
rect 6946 22267 7254 22276
rect 7392 22094 7420 24670
rect 7116 22066 7420 22094
rect 7472 22092 7524 22098
rect 7116 21894 7144 22066
rect 7472 22034 7524 22040
rect 7104 21888 7156 21894
rect 7104 21830 7156 21836
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20058 6776 20878
rect 6736 20052 6788 20058
rect 6736 19994 6788 20000
rect 6840 19904 6868 21558
rect 7116 21486 7144 21830
rect 7484 21690 7512 22034
rect 7472 21684 7524 21690
rect 7472 21626 7524 21632
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7288 21480 7340 21486
rect 7288 21422 7340 21428
rect 6946 21244 7254 21253
rect 6946 21242 6952 21244
rect 7008 21242 7032 21244
rect 7088 21242 7112 21244
rect 7168 21242 7192 21244
rect 7248 21242 7254 21244
rect 7008 21190 7010 21242
rect 7190 21190 7192 21242
rect 6946 21188 6952 21190
rect 7008 21188 7032 21190
rect 7088 21188 7112 21190
rect 7168 21188 7192 21190
rect 7248 21188 7254 21190
rect 6946 21179 7254 21188
rect 7300 20262 7328 21422
rect 7380 20324 7432 20330
rect 7380 20266 7432 20272
rect 7288 20256 7340 20262
rect 7288 20198 7340 20204
rect 6946 20156 7254 20165
rect 6946 20154 6952 20156
rect 7008 20154 7032 20156
rect 7088 20154 7112 20156
rect 7168 20154 7192 20156
rect 7248 20154 7254 20156
rect 7008 20102 7010 20154
rect 7190 20102 7192 20154
rect 6946 20100 6952 20102
rect 7008 20100 7032 20102
rect 7088 20100 7112 20102
rect 7168 20100 7192 20102
rect 7248 20100 7254 20102
rect 6946 20091 7254 20100
rect 7300 19922 7328 20198
rect 7392 20058 7420 20266
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 6920 19916 6972 19922
rect 6840 19876 6920 19904
rect 6920 19858 6972 19864
rect 7288 19916 7340 19922
rect 7288 19858 7340 19864
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 6932 19224 6960 19858
rect 7392 19768 7420 19858
rect 6840 19196 6960 19224
rect 7300 19740 7420 19768
rect 6840 18952 6868 19196
rect 6946 19068 7254 19077
rect 6946 19066 6952 19068
rect 7008 19066 7032 19068
rect 7088 19066 7112 19068
rect 7168 19066 7192 19068
rect 7248 19066 7254 19068
rect 7008 19014 7010 19066
rect 7190 19014 7192 19066
rect 6946 19012 6952 19014
rect 7008 19012 7032 19014
rect 7088 19012 7112 19014
rect 7168 19012 7192 19014
rect 7248 19012 7254 19014
rect 6946 19003 7254 19012
rect 6840 18924 6960 18952
rect 6932 18426 6960 18924
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 6932 18290 6960 18362
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 7196 18080 7248 18086
rect 7300 18068 7328 19740
rect 7248 18040 7328 18068
rect 7380 18080 7432 18086
rect 7196 18022 7248 18028
rect 7380 18022 7432 18028
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 6946 17980 7254 17989
rect 6946 17978 6952 17980
rect 7008 17978 7032 17980
rect 7088 17978 7112 17980
rect 7168 17978 7192 17980
rect 7248 17978 7254 17980
rect 7008 17926 7010 17978
rect 7190 17926 7192 17978
rect 6946 17924 6952 17926
rect 7008 17924 7032 17926
rect 7088 17924 7112 17926
rect 7168 17924 7192 17926
rect 7248 17924 7254 17926
rect 6946 17915 7254 17924
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7300 17134 7328 17818
rect 7392 17746 7420 18022
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7484 17626 7512 18022
rect 7392 17598 7512 17626
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 6946 16892 7254 16901
rect 6946 16890 6952 16892
rect 7008 16890 7032 16892
rect 7088 16890 7112 16892
rect 7168 16890 7192 16892
rect 7248 16890 7254 16892
rect 7008 16838 7010 16890
rect 7190 16838 7192 16890
rect 6946 16836 6952 16838
rect 7008 16836 7032 16838
rect 7088 16836 7112 16838
rect 7168 16836 7192 16838
rect 7248 16836 7254 16838
rect 6946 16827 7254 16836
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6748 16046 6776 16458
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6184 15972 6236 15978
rect 6184 15914 6236 15920
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6000 13388 6052 13394
rect 6000 13330 6052 13336
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5644 12374 5672 12582
rect 5736 12442 5764 12718
rect 5724 12436 5776 12442
rect 6104 12434 6132 14894
rect 6196 14550 6224 15914
rect 6828 15904 6880 15910
rect 6828 15846 6880 15852
rect 6840 15706 6868 15846
rect 6946 15804 7254 15813
rect 6946 15802 6952 15804
rect 7008 15802 7032 15804
rect 7088 15802 7112 15804
rect 7168 15802 7192 15804
rect 7248 15802 7254 15804
rect 7008 15750 7010 15802
rect 7190 15750 7192 15802
rect 6946 15748 6952 15750
rect 7008 15748 7032 15750
rect 7088 15748 7112 15750
rect 7168 15748 7192 15750
rect 7248 15748 7254 15750
rect 6946 15739 7254 15748
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 7300 15502 7328 17070
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 6286 15260 6594 15269
rect 6286 15258 6292 15260
rect 6348 15258 6372 15260
rect 6428 15258 6452 15260
rect 6508 15258 6532 15260
rect 6588 15258 6594 15260
rect 6348 15206 6350 15258
rect 6530 15206 6532 15258
rect 6286 15204 6292 15206
rect 6348 15204 6372 15206
rect 6428 15204 6452 15206
rect 6508 15204 6532 15206
rect 6588 15204 6594 15206
rect 6286 15195 6594 15204
rect 7300 15026 7328 15438
rect 7392 15162 7420 17598
rect 7576 17218 7604 31962
rect 8680 31958 8708 33646
rect 9678 33544 9734 34344
rect 11610 33544 11666 34344
rect 12898 33544 12954 34344
rect 14186 33544 14242 34344
rect 16118 33544 16174 34344
rect 17406 33544 17462 34344
rect 18694 33544 18750 34344
rect 20626 33544 20682 34344
rect 21914 33544 21970 34344
rect 23846 33544 23902 34344
rect 25134 33544 25190 34344
rect 26422 33544 26478 34344
rect 28354 33544 28410 34344
rect 29642 33674 29698 34344
rect 29642 33646 29960 33674
rect 29642 33544 29698 33646
rect 9692 32026 9720 33544
rect 11624 32026 11652 33544
rect 9680 32020 9732 32026
rect 9680 31962 9732 31968
rect 11612 32020 11664 32026
rect 11612 31962 11664 31968
rect 8668 31952 8720 31958
rect 8668 31894 8720 31900
rect 9680 31884 9732 31890
rect 9680 31826 9732 31832
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 9692 30258 9720 31826
rect 11888 31680 11940 31686
rect 11888 31622 11940 31628
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11796 31136 11848 31142
rect 11796 31078 11848 31084
rect 9680 30252 9732 30258
rect 9680 30194 9732 30200
rect 7656 30048 7708 30054
rect 7656 29990 7708 29996
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8760 30048 8812 30054
rect 8760 29990 8812 29996
rect 7668 29102 7696 29990
rect 8312 29782 8340 29990
rect 8300 29776 8352 29782
rect 8300 29718 8352 29724
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8312 29306 8340 29582
rect 8300 29300 8352 29306
rect 8300 29242 8352 29248
rect 8392 29232 8444 29238
rect 8392 29174 8444 29180
rect 7656 29096 7708 29102
rect 7656 29038 7708 29044
rect 8404 28626 8432 29174
rect 8772 29102 8800 29990
rect 9692 29850 9720 30194
rect 10324 30116 10376 30122
rect 10324 30058 10376 30064
rect 10336 29850 10364 30058
rect 9680 29844 9732 29850
rect 9680 29786 9732 29792
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10796 29170 10824 31078
rect 10876 30728 10928 30734
rect 10876 30670 10928 30676
rect 10888 30258 10916 30670
rect 10876 30252 10928 30258
rect 10876 30194 10928 30200
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 8760 29096 8812 29102
rect 8760 29038 8812 29044
rect 8852 29096 8904 29102
rect 8852 29038 8904 29044
rect 8864 28762 8892 29038
rect 9956 29028 10008 29034
rect 9956 28970 10008 28976
rect 8852 28756 8904 28762
rect 8852 28698 8904 28704
rect 8392 28620 8444 28626
rect 8392 28562 8444 28568
rect 9496 28552 9548 28558
rect 9496 28494 9548 28500
rect 7840 28416 7892 28422
rect 7840 28358 7892 28364
rect 7852 27946 7880 28358
rect 9508 28218 9536 28494
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 7840 27940 7892 27946
rect 7840 27882 7892 27888
rect 9036 27872 9088 27878
rect 9036 27814 9088 27820
rect 8944 27668 8996 27674
rect 8944 27610 8996 27616
rect 8116 27464 8168 27470
rect 8116 27406 8168 27412
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7668 24274 7696 27270
rect 8128 27130 8156 27406
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8116 27124 8168 27130
rect 8116 27066 8168 27072
rect 7748 26852 7800 26858
rect 7748 26794 7800 26800
rect 7760 26586 7788 26794
rect 7840 26784 7892 26790
rect 7840 26726 7892 26732
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7852 26450 7880 26726
rect 8404 26586 8432 27270
rect 8484 26852 8536 26858
rect 8484 26794 8536 26800
rect 8392 26580 8444 26586
rect 8392 26522 8444 26528
rect 7840 26444 7892 26450
rect 7840 26386 7892 26392
rect 7748 25764 7800 25770
rect 7748 25706 7800 25712
rect 7760 25498 7788 25706
rect 7852 25702 7880 26386
rect 8496 26382 8524 26794
rect 8772 26586 8800 27270
rect 8956 27062 8984 27610
rect 9048 27538 9076 27814
rect 9692 27606 9720 28358
rect 9864 28008 9916 28014
rect 9864 27950 9916 27956
rect 9772 27940 9824 27946
rect 9772 27882 9824 27888
rect 9680 27600 9732 27606
rect 9218 27568 9274 27577
rect 9036 27532 9088 27538
rect 9600 27560 9680 27588
rect 9274 27526 9352 27554
rect 9218 27503 9274 27512
rect 9036 27474 9088 27480
rect 8944 27056 8996 27062
rect 8944 26998 8996 27004
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8484 26376 8536 26382
rect 8484 26318 8536 26324
rect 8116 26240 8168 26246
rect 8116 26182 8168 26188
rect 7840 25696 7892 25702
rect 7840 25638 7892 25644
rect 7748 25492 7800 25498
rect 7748 25434 7800 25440
rect 7852 25362 7880 25638
rect 7840 25356 7892 25362
rect 7840 25298 7892 25304
rect 8128 25226 8156 26182
rect 8496 25838 8524 26318
rect 8484 25832 8536 25838
rect 8484 25774 8536 25780
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8220 25498 8248 25706
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8208 25492 8260 25498
rect 8208 25434 8260 25440
rect 8116 25220 8168 25226
rect 8116 25162 8168 25168
rect 8588 24954 8616 25638
rect 8576 24948 8628 24954
rect 8576 24890 8628 24896
rect 8956 24410 8984 26998
rect 9324 26518 9352 27526
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9416 26586 9444 26862
rect 9600 26858 9628 27560
rect 9680 27542 9732 27548
rect 9784 27402 9812 27882
rect 9772 27396 9824 27402
rect 9772 27338 9824 27344
rect 9876 27130 9904 27950
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 9968 26994 9996 28970
rect 10888 28626 10916 30194
rect 11244 29640 11296 29646
rect 11244 29582 11296 29588
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 10876 28620 10928 28626
rect 10876 28562 10928 28568
rect 10232 28552 10284 28558
rect 10232 28494 10284 28500
rect 10244 28218 10272 28494
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 10888 28150 10916 28562
rect 10876 28144 10928 28150
rect 10876 28086 10928 28092
rect 10600 28008 10652 28014
rect 10600 27950 10652 27956
rect 10508 27940 10560 27946
rect 10508 27882 10560 27888
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 10336 27674 10364 27814
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 10324 27464 10376 27470
rect 10324 27406 10376 27412
rect 10048 27328 10100 27334
rect 10048 27270 10100 27276
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 9680 26920 9732 26926
rect 9680 26862 9732 26868
rect 9588 26852 9640 26858
rect 9588 26794 9640 26800
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9312 26512 9364 26518
rect 9312 26454 9364 26460
rect 9036 26444 9088 26450
rect 9036 26386 9088 26392
rect 9048 26042 9076 26386
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 9128 24676 9180 24682
rect 9128 24618 9180 24624
rect 7748 24404 7800 24410
rect 7748 24346 7800 24352
rect 8944 24404 8996 24410
rect 8944 24346 8996 24352
rect 7656 24268 7708 24274
rect 7656 24210 7708 24216
rect 7668 23746 7696 24210
rect 7760 23866 7788 24346
rect 9140 24342 9168 24618
rect 9128 24336 9180 24342
rect 9128 24278 9180 24284
rect 9036 24268 9088 24274
rect 9036 24210 9088 24216
rect 8760 24064 8812 24070
rect 8760 24006 8812 24012
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 7840 23860 7892 23866
rect 7840 23802 7892 23808
rect 7668 23718 7788 23746
rect 7760 23662 7788 23718
rect 7748 23656 7800 23662
rect 7748 23598 7800 23604
rect 7656 23588 7708 23594
rect 7656 23530 7708 23536
rect 7668 22982 7696 23530
rect 7748 23520 7800 23526
rect 7748 23462 7800 23468
rect 7760 23186 7788 23462
rect 7748 23180 7800 23186
rect 7748 23122 7800 23128
rect 7656 22976 7708 22982
rect 7656 22918 7708 22924
rect 7668 22438 7696 22918
rect 7656 22432 7708 22438
rect 7656 22374 7708 22380
rect 7852 22094 7880 23802
rect 8772 23730 8800 24006
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 8760 23724 8812 23730
rect 8760 23666 8812 23672
rect 8116 23588 8168 23594
rect 8116 23530 8168 23536
rect 8128 23050 8156 23530
rect 8208 23248 8260 23254
rect 8208 23190 8260 23196
rect 8116 23044 8168 23050
rect 8116 22986 8168 22992
rect 7760 22066 7880 22094
rect 7656 18080 7708 18086
rect 7760 18068 7788 22066
rect 8220 22030 8248 23190
rect 8404 23118 8432 23666
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8668 23112 8720 23118
rect 8668 23054 8720 23060
rect 8404 22642 8432 23054
rect 8680 22778 8708 23054
rect 8668 22772 8720 22778
rect 8668 22714 8720 22720
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21690 7972 21830
rect 8128 21690 8156 21966
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 8116 21684 8168 21690
rect 8116 21626 8168 21632
rect 7944 21486 7972 21626
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 8024 21344 8076 21350
rect 8024 21286 8076 21292
rect 8036 20534 8064 21286
rect 8220 20942 8248 21966
rect 8404 21554 8432 22578
rect 9048 22094 9076 24210
rect 9232 22094 9260 26250
rect 9588 26240 9640 26246
rect 9692 26234 9720 26862
rect 10060 26790 10088 27270
rect 10336 27130 10364 27406
rect 10324 27124 10376 27130
rect 10324 27066 10376 27072
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 10048 26784 10100 26790
rect 10048 26726 10100 26732
rect 9640 26206 9720 26234
rect 9588 26182 9640 26188
rect 9600 26042 9628 26182
rect 9588 26036 9640 26042
rect 9588 25978 9640 25984
rect 9404 25832 9456 25838
rect 9404 25774 9456 25780
rect 9312 25696 9364 25702
rect 9312 25638 9364 25644
rect 9324 25498 9352 25638
rect 9312 25492 9364 25498
rect 9312 25434 9364 25440
rect 9312 25288 9364 25294
rect 9312 25230 9364 25236
rect 9324 24954 9352 25230
rect 9416 24954 9444 25774
rect 9600 25702 9628 25978
rect 9588 25696 9640 25702
rect 9588 25638 9640 25644
rect 9600 25158 9628 25638
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9312 24948 9364 24954
rect 9312 24890 9364 24896
rect 9404 24948 9456 24954
rect 9404 24890 9456 24896
rect 9600 24750 9628 25094
rect 9692 24750 9720 25298
rect 9588 24744 9640 24750
rect 9588 24686 9640 24692
rect 9680 24744 9732 24750
rect 9876 24721 9904 26726
rect 10060 26246 10088 26726
rect 10324 26580 10376 26586
rect 10324 26522 10376 26528
rect 10048 26240 10100 26246
rect 10048 26182 10100 26188
rect 10060 25362 10088 26182
rect 10336 26042 10364 26522
rect 10520 26246 10548 27882
rect 10612 27062 10640 27950
rect 10888 27690 10916 28086
rect 11164 28014 11192 29106
rect 11256 29034 11284 29582
rect 11244 29028 11296 29034
rect 11244 28970 11296 28976
rect 11152 28008 11204 28014
rect 11152 27950 11204 27956
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 11072 27713 11100 27882
rect 11058 27704 11114 27713
rect 10888 27662 11008 27690
rect 10980 27588 11008 27662
rect 11058 27639 11114 27648
rect 10980 27560 11100 27588
rect 10600 27056 10652 27062
rect 10600 26998 10652 27004
rect 10612 26586 10640 26998
rect 10968 26920 11020 26926
rect 10968 26862 11020 26868
rect 10600 26580 10652 26586
rect 10600 26522 10652 26528
rect 10876 26512 10928 26518
rect 10876 26454 10928 26460
rect 10600 26444 10652 26450
rect 10600 26386 10652 26392
rect 10508 26240 10560 26246
rect 10508 26182 10560 26188
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10520 25786 10548 26182
rect 10612 25838 10640 26386
rect 10888 26042 10916 26454
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10428 25758 10548 25786
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10784 25832 10836 25838
rect 10784 25774 10836 25780
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 10324 25356 10376 25362
rect 10324 25298 10376 25304
rect 10060 24954 10088 25298
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 10048 24948 10100 24954
rect 10048 24890 10100 24896
rect 10152 24750 10180 25094
rect 9956 24744 10008 24750
rect 9680 24686 9732 24692
rect 9862 24712 9918 24721
rect 9600 24562 9628 24686
rect 9956 24686 10008 24692
rect 10140 24744 10192 24750
rect 10336 24698 10364 25298
rect 10140 24686 10192 24692
rect 9862 24647 9918 24656
rect 9600 24534 9720 24562
rect 9692 23322 9720 24534
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9784 22234 9812 22510
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9048 22066 9168 22094
rect 9232 22066 9352 22094
rect 8484 22024 8536 22030
rect 8484 21966 8536 21972
rect 8496 21622 8524 21966
rect 8484 21616 8536 21622
rect 8484 21558 8536 21564
rect 8392 21548 8444 21554
rect 8392 21490 8444 21496
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 8036 19854 8064 20470
rect 8404 20466 8432 21490
rect 8392 20460 8444 20466
rect 8392 20402 8444 20408
rect 8944 20324 8996 20330
rect 8944 20266 8996 20272
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8128 19990 8156 20198
rect 8956 20058 8984 20266
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 8024 19848 8076 19854
rect 8024 19790 8076 19796
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7708 18040 7788 18068
rect 7656 18022 7708 18028
rect 7852 17610 7880 19246
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7944 18290 7972 18702
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7932 17808 7984 17814
rect 7932 17750 7984 17756
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7484 17190 7604 17218
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6564 14618 6592 14758
rect 6946 14716 7254 14725
rect 6946 14714 6952 14716
rect 7008 14714 7032 14716
rect 7088 14714 7112 14716
rect 7168 14714 7192 14716
rect 7248 14714 7254 14716
rect 7008 14662 7010 14714
rect 7190 14662 7192 14714
rect 6946 14660 6952 14662
rect 7008 14660 7032 14662
rect 7088 14660 7112 14662
rect 7168 14660 7192 14662
rect 7248 14660 7254 14662
rect 6946 14651 7254 14660
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6184 14544 6236 14550
rect 6184 14486 6236 14492
rect 6286 14172 6594 14181
rect 6286 14170 6292 14172
rect 6348 14170 6372 14172
rect 6428 14170 6452 14172
rect 6508 14170 6532 14172
rect 6588 14170 6594 14172
rect 6348 14118 6350 14170
rect 6530 14118 6532 14170
rect 6286 14116 6292 14118
rect 6348 14116 6372 14118
rect 6428 14116 6452 14118
rect 6508 14116 6532 14118
rect 6588 14116 6594 14118
rect 6286 14107 6594 14116
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6286 13084 6594 13093
rect 6286 13082 6292 13084
rect 6348 13082 6372 13084
rect 6428 13082 6452 13084
rect 6508 13082 6532 13084
rect 6588 13082 6594 13084
rect 6348 13030 6350 13082
rect 6530 13030 6532 13082
rect 6286 13028 6292 13030
rect 6348 13028 6372 13030
rect 6428 13028 6452 13030
rect 6508 13028 6532 13030
rect 6588 13028 6594 13030
rect 6286 13019 6594 13028
rect 6656 12986 6684 14010
rect 7300 13938 7328 14962
rect 7380 14544 7432 14550
rect 7380 14486 7432 14492
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 6946 13628 7254 13637
rect 6946 13626 6952 13628
rect 7008 13626 7032 13628
rect 7088 13626 7112 13628
rect 7168 13626 7192 13628
rect 7248 13626 7254 13628
rect 7008 13574 7010 13626
rect 7190 13574 7192 13626
rect 6946 13572 6952 13574
rect 7008 13572 7032 13574
rect 7088 13572 7112 13574
rect 7168 13572 7192 13574
rect 7248 13572 7254 13574
rect 6946 13563 7254 13572
rect 7288 13252 7340 13258
rect 7288 13194 7340 13200
rect 6644 12980 6696 12986
rect 6644 12922 6696 12928
rect 5724 12378 5776 12384
rect 5920 12406 6132 12434
rect 5632 12368 5684 12374
rect 5632 12310 5684 12316
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 10198 5580 11494
rect 5644 11354 5672 12174
rect 5632 11348 5684 11354
rect 5632 11290 5684 11296
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5356 6248 5408 6254
rect 5356 6190 5408 6196
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 4344 5160 4396 5166
rect 4344 5102 4396 5108
rect 5368 4826 5396 5646
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4448 2990 4476 4762
rect 5736 3602 5764 12242
rect 5816 11552 5868 11558
rect 5816 11494 5868 11500
rect 5828 11286 5856 11494
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5920 10810 5948 12406
rect 6656 12238 6684 12922
rect 6840 12702 6960 12730
rect 6840 12434 6868 12702
rect 6932 12646 6960 12702
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6946 12540 7254 12549
rect 6946 12538 6952 12540
rect 7008 12538 7032 12540
rect 7088 12538 7112 12540
rect 7168 12538 7192 12540
rect 7248 12538 7254 12540
rect 7008 12486 7010 12538
rect 7190 12486 7192 12538
rect 6946 12484 6952 12486
rect 7008 12484 7032 12486
rect 7088 12484 7112 12486
rect 7168 12484 7192 12486
rect 7248 12484 7254 12486
rect 6946 12475 7254 12484
rect 7300 12434 7328 13194
rect 7392 12986 7420 14486
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 6840 12406 6960 12434
rect 6932 12374 6960 12406
rect 7116 12406 7328 12434
rect 6920 12368 6972 12374
rect 6918 12336 6920 12345
rect 6972 12336 6974 12345
rect 6828 12300 6880 12306
rect 7116 12306 7144 12406
rect 7392 12306 7420 12922
rect 6918 12271 6974 12280
rect 7104 12300 7156 12306
rect 6828 12242 6880 12248
rect 7104 12242 7156 12248
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6286 11996 6594 12005
rect 6286 11994 6292 11996
rect 6348 11994 6372 11996
rect 6428 11994 6452 11996
rect 6508 11994 6532 11996
rect 6588 11994 6594 11996
rect 6348 11942 6350 11994
rect 6530 11942 6532 11994
rect 6286 11940 6292 11942
rect 6348 11940 6372 11942
rect 6428 11940 6452 11942
rect 6508 11940 6532 11942
rect 6588 11940 6594 11942
rect 6286 11931 6594 11940
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6012 10674 6040 11834
rect 6656 11778 6684 12174
rect 6840 11898 6868 12242
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6656 11750 6776 11778
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6104 11354 6132 11630
rect 6656 11354 6684 11630
rect 6092 11348 6144 11354
rect 6092 11290 6144 11296
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 6104 10062 6132 11290
rect 6748 11218 6776 11750
rect 6946 11452 7254 11461
rect 6946 11450 6952 11452
rect 7008 11450 7032 11452
rect 7088 11450 7112 11452
rect 7168 11450 7192 11452
rect 7248 11450 7254 11452
rect 7008 11398 7010 11450
rect 7190 11398 7192 11450
rect 6946 11396 6952 11398
rect 7008 11396 7032 11398
rect 7088 11396 7112 11398
rect 7168 11396 7192 11398
rect 7248 11396 7254 11398
rect 6946 11387 7254 11396
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6286 10908 6594 10917
rect 6286 10906 6292 10908
rect 6348 10906 6372 10908
rect 6428 10906 6452 10908
rect 6508 10906 6532 10908
rect 6588 10906 6594 10908
rect 6348 10854 6350 10906
rect 6530 10854 6532 10906
rect 6286 10852 6292 10854
rect 6348 10852 6372 10854
rect 6428 10852 6452 10854
rect 6508 10852 6532 10854
rect 6588 10852 6594 10854
rect 6286 10843 6594 10852
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6288 10266 6316 10406
rect 6380 10266 6408 10746
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6104 7886 6132 9998
rect 6286 9820 6594 9829
rect 6286 9818 6292 9820
rect 6348 9818 6372 9820
rect 6428 9818 6452 9820
rect 6508 9818 6532 9820
rect 6588 9818 6594 9820
rect 6348 9766 6350 9818
rect 6530 9766 6532 9818
rect 6286 9764 6292 9766
rect 6348 9764 6372 9766
rect 6428 9764 6452 9766
rect 6508 9764 6532 9766
rect 6588 9764 6594 9766
rect 6286 9755 6594 9764
rect 6748 9178 6776 11154
rect 6946 10364 7254 10373
rect 6946 10362 6952 10364
rect 7008 10362 7032 10364
rect 7088 10362 7112 10364
rect 7168 10362 7192 10364
rect 7248 10362 7254 10364
rect 7008 10310 7010 10362
rect 7190 10310 7192 10362
rect 6946 10308 6952 10310
rect 7008 10308 7032 10310
rect 7088 10308 7112 10310
rect 7168 10308 7192 10310
rect 7248 10308 7254 10310
rect 6946 10299 7254 10308
rect 6946 9276 7254 9285
rect 6946 9274 6952 9276
rect 7008 9274 7032 9276
rect 7088 9274 7112 9276
rect 7168 9274 7192 9276
rect 7248 9274 7254 9276
rect 7008 9222 7010 9274
rect 7190 9222 7192 9274
rect 6946 9220 6952 9222
rect 7008 9220 7032 9222
rect 7088 9220 7112 9222
rect 7168 9220 7192 9222
rect 7248 9220 7254 9222
rect 6946 9211 7254 9220
rect 7484 9178 7512 17190
rect 7944 16794 7972 17750
rect 8128 17202 8156 18566
rect 8772 18426 8800 19110
rect 8864 18698 8892 19110
rect 8956 18902 8984 19110
rect 8944 18896 8996 18902
rect 8944 18838 8996 18844
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8208 18420 8260 18426
rect 8208 18362 8260 18368
rect 8760 18420 8812 18426
rect 8760 18362 8812 18368
rect 8116 17196 8168 17202
rect 8116 17138 8168 17144
rect 8220 16810 8248 18362
rect 9140 18306 9168 22066
rect 9324 20262 9352 22066
rect 9588 21956 9640 21962
rect 9588 21898 9640 21904
rect 9600 21554 9628 21898
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 21554 9720 21830
rect 9588 21548 9640 21554
rect 9588 21490 9640 21496
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9600 21010 9628 21490
rect 9680 21344 9732 21350
rect 9680 21286 9732 21292
rect 9588 21004 9640 21010
rect 9588 20946 9640 20952
rect 9692 20602 9720 21286
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9678 20496 9734 20505
rect 9588 20460 9640 20466
rect 9678 20431 9734 20440
rect 9588 20402 9640 20408
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9324 19922 9352 20198
rect 9600 19922 9628 20402
rect 9692 19922 9720 20431
rect 9876 19990 9904 24647
rect 9968 23225 9996 24686
rect 10244 24670 10364 24698
rect 9954 23216 10010 23225
rect 9954 23151 10010 23160
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10152 22012 10180 22374
rect 10244 22094 10272 24670
rect 10428 22234 10456 25758
rect 10508 25696 10560 25702
rect 10508 25638 10560 25644
rect 10416 22228 10468 22234
rect 10416 22170 10468 22176
rect 10244 22066 10364 22094
rect 10232 22024 10284 22030
rect 10152 21984 10232 22012
rect 10232 21966 10284 21972
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9968 21486 9996 21830
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 10060 21078 10088 21830
rect 10244 21418 10272 21966
rect 10232 21412 10284 21418
rect 10232 21354 10284 21360
rect 10048 21072 10100 21078
rect 10048 21014 10100 21020
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10060 20058 10088 20334
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9864 19984 9916 19990
rect 9864 19926 9916 19932
rect 10244 19922 10272 21354
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9680 19916 9732 19922
rect 9680 19858 9732 19864
rect 9772 19916 9824 19922
rect 9772 19858 9824 19864
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 9232 19310 9260 19654
rect 9600 19378 9628 19858
rect 9784 19786 9812 19858
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9220 19304 9272 19310
rect 9272 19264 9444 19292
rect 9220 19246 9272 19252
rect 9416 19174 9444 19264
rect 9784 19174 9812 19722
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10048 19372 10100 19378
rect 10048 19314 10100 19320
rect 9862 19272 9918 19281
rect 9862 19207 9918 19216
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9876 18902 9904 19207
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 9864 18896 9916 18902
rect 9864 18838 9916 18844
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18358 9720 18770
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9864 18760 9916 18766
rect 9864 18702 9916 18708
rect 9680 18352 9732 18358
rect 8392 18284 8444 18290
rect 9140 18278 9260 18306
rect 9680 18294 9732 18300
rect 8392 18226 8444 18232
rect 8404 18154 8432 18226
rect 8392 18148 8444 18154
rect 8392 18090 8444 18096
rect 9128 18148 9180 18154
rect 9128 18090 9180 18096
rect 8852 17808 8904 17814
rect 8852 17750 8904 17756
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8312 17338 8340 17614
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8220 16794 8340 16810
rect 8496 16794 8524 17002
rect 8864 16794 8892 17750
rect 9140 16794 9168 18090
rect 7932 16788 7984 16794
rect 8220 16788 8352 16794
rect 8220 16782 8300 16788
rect 7932 16730 7984 16736
rect 8300 16730 8352 16736
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 7564 15904 7616 15910
rect 7564 15846 7616 15852
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7576 14890 7604 15846
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7668 14618 7696 15438
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7944 14498 7972 15846
rect 8024 14884 8076 14890
rect 8024 14826 8076 14832
rect 8036 14618 8064 14826
rect 8496 14618 8524 15982
rect 8576 15972 8628 15978
rect 8576 15914 8628 15920
rect 8588 15366 8616 15914
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 14618 8984 15302
rect 9048 15162 9076 15438
rect 9232 15162 9260 18278
rect 9692 17746 9720 18294
rect 9784 17882 9812 18702
rect 9876 18426 9904 18702
rect 9864 18420 9916 18426
rect 9864 18362 9916 18368
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9784 17202 9812 17818
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9036 15156 9088 15162
rect 9036 15098 9088 15104
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 8484 14612 8536 14618
rect 8484 14554 8536 14560
rect 8944 14612 8996 14618
rect 8944 14554 8996 14560
rect 7944 14482 8064 14498
rect 7944 14476 8076 14482
rect 7944 14470 8024 14476
rect 8024 14418 8076 14424
rect 7746 14376 7802 14385
rect 7746 14311 7748 14320
rect 7800 14311 7802 14320
rect 7748 14282 7800 14288
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7668 13530 7696 13738
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 8036 13326 8064 14418
rect 9048 14414 9076 14758
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8496 14074 8524 14214
rect 9140 14074 9168 14350
rect 9692 14346 9720 17070
rect 9968 17066 9996 19110
rect 10060 18766 10088 19314
rect 10048 18760 10100 18766
rect 10048 18702 10100 18708
rect 10060 18222 10088 18702
rect 10140 18692 10192 18698
rect 10140 18634 10192 18640
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10060 17202 10088 18158
rect 10152 18086 10180 18634
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10152 17814 10180 18022
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 10048 17196 10100 17202
rect 10048 17138 10100 17144
rect 9956 17060 10008 17066
rect 9956 17002 10008 17008
rect 10152 16658 10180 17614
rect 10244 16998 10272 19654
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12714 8064 13262
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7944 12442 7972 12582
rect 8036 12458 8064 12650
rect 8114 12472 8170 12481
rect 7932 12436 7984 12442
rect 8036 12430 8114 12458
rect 8114 12407 8116 12416
rect 7932 12378 7984 12384
rect 8168 12407 8170 12416
rect 8116 12378 8168 12384
rect 7840 12368 7892 12374
rect 8220 12322 8248 13874
rect 8300 13184 8352 13190
rect 8300 13126 8352 13132
rect 8312 12986 8340 13126
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8484 12708 8536 12714
rect 8484 12650 8536 12656
rect 7840 12310 7892 12316
rect 7852 11898 7880 12310
rect 8036 12306 8248 12322
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 8024 12300 8248 12306
rect 8076 12294 8248 12300
rect 8024 12242 8076 12248
rect 7840 11892 7892 11898
rect 7944 11880 7972 12242
rect 8024 11892 8076 11898
rect 7944 11852 8024 11880
rect 7840 11834 7892 11840
rect 8024 11834 8076 11840
rect 7748 11620 7800 11626
rect 7748 11562 7800 11568
rect 7760 11354 7788 11562
rect 7852 11354 7880 11834
rect 8496 11762 8524 12650
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8588 12442 8616 12582
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8772 12374 8800 12718
rect 9140 12434 9168 14010
rect 9692 12434 9720 14282
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9784 13462 9812 13670
rect 9772 13456 9824 13462
rect 9772 13398 9824 13404
rect 9772 13320 9824 13326
rect 9772 13262 9824 13268
rect 9784 12442 9812 13262
rect 9140 12406 9260 12434
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8484 11756 8536 11762
rect 8484 11698 8536 11704
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11354 8432 11494
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8036 10674 8064 10950
rect 8588 10810 8616 11562
rect 8680 11286 8708 11698
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8864 11150 8892 12038
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9140 11354 9168 11494
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9140 11218 9168 11290
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8024 10668 8076 10674
rect 8024 10610 8076 10616
rect 8668 10464 8720 10470
rect 8668 10406 8720 10412
rect 8680 9586 8708 10406
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 6286 8732 6594 8741
rect 6286 8730 6292 8732
rect 6348 8730 6372 8732
rect 6428 8730 6452 8732
rect 6508 8730 6532 8732
rect 6588 8730 6594 8732
rect 6348 8678 6350 8730
rect 6530 8678 6532 8730
rect 6286 8676 6292 8678
rect 6348 8676 6372 8678
rect 6428 8676 6452 8678
rect 6508 8676 6532 8678
rect 6588 8676 6594 8678
rect 6286 8667 6594 8676
rect 6748 8498 6776 9114
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6196 7886 6224 8230
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6104 5710 6132 7822
rect 6286 7644 6594 7653
rect 6286 7642 6292 7644
rect 6348 7642 6372 7644
rect 6428 7642 6452 7644
rect 6508 7642 6532 7644
rect 6588 7642 6594 7644
rect 6348 7590 6350 7642
rect 6530 7590 6532 7642
rect 6286 7588 6292 7590
rect 6348 7588 6372 7590
rect 6428 7588 6452 7590
rect 6508 7588 6532 7590
rect 6588 7588 6594 7590
rect 6286 7579 6594 7588
rect 6286 6556 6594 6565
rect 6286 6554 6292 6556
rect 6348 6554 6372 6556
rect 6428 6554 6452 6556
rect 6508 6554 6532 6556
rect 6588 6554 6594 6556
rect 6348 6502 6350 6554
rect 6530 6502 6532 6554
rect 6286 6500 6292 6502
rect 6348 6500 6372 6502
rect 6428 6500 6452 6502
rect 6508 6500 6532 6502
rect 6588 6500 6594 6502
rect 6286 6491 6594 6500
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6656 5914 6684 6054
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6092 5704 6144 5710
rect 6092 5646 6144 5652
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6012 5166 6040 5510
rect 6104 5234 6132 5646
rect 6286 5468 6594 5477
rect 6286 5466 6292 5468
rect 6348 5466 6372 5468
rect 6428 5466 6452 5468
rect 6508 5466 6532 5468
rect 6588 5466 6594 5468
rect 6348 5414 6350 5466
rect 6530 5414 6532 5466
rect 6286 5412 6292 5414
rect 6348 5412 6372 5414
rect 6428 5412 6452 5414
rect 6508 5412 6532 5414
rect 6588 5412 6594 5414
rect 6286 5403 6594 5412
rect 6748 5370 6776 8434
rect 8312 8430 8340 9318
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 6946 8188 7254 8197
rect 6946 8186 6952 8188
rect 7008 8186 7032 8188
rect 7088 8186 7112 8188
rect 7168 8186 7192 8188
rect 7248 8186 7254 8188
rect 7008 8134 7010 8186
rect 7190 8134 7192 8186
rect 6946 8132 6952 8134
rect 7008 8132 7032 8134
rect 7088 8132 7112 8134
rect 7168 8132 7192 8134
rect 7248 8132 7254 8134
rect 6946 8123 7254 8132
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6840 5794 6868 7754
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 6946 7100 7254 7109
rect 6946 7098 6952 7100
rect 7008 7098 7032 7100
rect 7088 7098 7112 7100
rect 7168 7098 7192 7100
rect 7248 7098 7254 7100
rect 7008 7046 7010 7098
rect 7190 7046 7192 7098
rect 6946 7044 6952 7046
rect 7008 7044 7032 7046
rect 7088 7044 7112 7046
rect 7168 7044 7192 7046
rect 7248 7044 7254 7046
rect 6946 7035 7254 7044
rect 7668 6934 7696 7482
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 6920 6656 6972 6662
rect 6920 6598 6972 6604
rect 6932 6458 6960 6598
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 7208 6118 7236 6802
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 6946 6012 7254 6021
rect 6946 6010 6952 6012
rect 7008 6010 7032 6012
rect 7088 6010 7112 6012
rect 7168 6010 7192 6012
rect 7248 6010 7254 6012
rect 7008 5958 7010 6010
rect 7190 5958 7192 6010
rect 6946 5956 6952 5958
rect 7008 5956 7032 5958
rect 7088 5956 7112 5958
rect 7168 5956 7192 5958
rect 7248 5956 7254 5958
rect 6946 5947 7254 5956
rect 6840 5766 6960 5794
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 6012 4622 6040 4966
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6104 4486 6132 5170
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 6104 4146 6132 4422
rect 6286 4380 6594 4389
rect 6286 4378 6292 4380
rect 6348 4378 6372 4380
rect 6428 4378 6452 4380
rect 6508 4378 6532 4380
rect 6588 4378 6594 4380
rect 6348 4326 6350 4378
rect 6530 4326 6532 4378
rect 6286 4324 6292 4326
rect 6348 4324 6372 4326
rect 6428 4324 6452 4326
rect 6508 4324 6532 4326
rect 6588 4324 6594 4326
rect 6286 4315 6594 4324
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6656 3992 6684 4966
rect 6748 4622 6776 5306
rect 6932 5166 6960 5766
rect 7576 5302 7604 6054
rect 7852 5914 7880 6190
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 8220 5166 8248 5714
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5370 8340 5510
rect 8300 5364 8352 5370
rect 8300 5306 8352 5312
rect 9048 5234 9076 6054
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6840 4826 6868 5034
rect 6946 4924 7254 4933
rect 6946 4922 6952 4924
rect 7008 4922 7032 4924
rect 7088 4922 7112 4924
rect 7168 4922 7192 4924
rect 7248 4922 7254 4924
rect 7008 4870 7010 4922
rect 7190 4870 7192 4922
rect 6946 4868 6952 4870
rect 7008 4868 7032 4870
rect 7088 4868 7112 4870
rect 7168 4868 7192 4870
rect 7248 4868 7254 4870
rect 6946 4859 7254 4868
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6736 4616 6788 4622
rect 6788 4564 6868 4570
rect 6736 4558 6868 4564
rect 6748 4542 6868 4558
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 4282 6776 4422
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 6736 4004 6788 4010
rect 6656 3964 6736 3992
rect 6736 3946 6788 3952
rect 6840 3670 6868 4542
rect 7668 4282 7696 5102
rect 8220 4690 8248 5102
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 7656 4276 7708 4282
rect 7656 4218 7708 4224
rect 6946 3836 7254 3845
rect 6946 3834 6952 3836
rect 7008 3834 7032 3836
rect 7088 3834 7112 3836
rect 7168 3834 7192 3836
rect 7248 3834 7254 3836
rect 7008 3782 7010 3834
rect 7190 3782 7192 3834
rect 6946 3780 6952 3782
rect 7008 3780 7032 3782
rect 7088 3780 7112 3782
rect 7168 3780 7192 3782
rect 7248 3780 7254 3782
rect 6946 3771 7254 3780
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 3608 2916 3660 2922
rect 3608 2858 3660 2864
rect 3620 2825 3648 2858
rect 3606 2816 3662 2825
rect 3606 2751 3662 2760
rect 3054 1456 3110 1465
rect 3054 1391 3110 1400
rect 4540 800 4568 3470
rect 6286 3292 6594 3301
rect 6286 3290 6292 3292
rect 6348 3290 6372 3292
rect 6428 3290 6452 3292
rect 6508 3290 6532 3292
rect 6588 3290 6594 3292
rect 6348 3238 6350 3290
rect 6530 3238 6532 3290
rect 6286 3236 6292 3238
rect 6348 3236 6372 3238
rect 6428 3236 6452 3238
rect 6508 3236 6532 3238
rect 6588 3236 6594 3238
rect 6286 3227 6594 3236
rect 7668 2990 7696 4218
rect 9232 2990 9260 12406
rect 9324 12406 9720 12434
rect 9772 12436 9824 12442
rect 9324 11218 9352 12406
rect 9772 12378 9824 12384
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 9324 10266 9352 11154
rect 9508 11150 9536 11630
rect 9692 11218 9720 12106
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9784 11898 9812 12038
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9876 11218 9904 14554
rect 9680 11212 9732 11218
rect 9680 11154 9732 11160
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9588 11144 9640 11150
rect 9588 11086 9640 11092
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9324 9674 9352 10202
rect 9324 9646 9444 9674
rect 9416 7546 9444 9646
rect 9600 9382 9628 11086
rect 9692 10656 9720 11154
rect 9692 10628 9812 10656
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9692 10266 9720 10474
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9784 10198 9812 10628
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9416 6798 9444 7482
rect 9404 6792 9456 6798
rect 9404 6734 9456 6740
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9784 5914 9812 6190
rect 9968 5914 9996 15098
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10060 13394 10088 13874
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10152 12306 10180 16594
rect 10244 14278 10272 16934
rect 10336 14618 10364 22066
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10428 19922 10456 21286
rect 10520 20602 10548 25638
rect 10796 25362 10824 25774
rect 10888 25378 10916 25978
rect 10980 25974 11008 26862
rect 11072 26466 11100 27560
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 11164 26858 11192 27066
rect 11256 26994 11284 28970
rect 11244 26988 11296 26994
rect 11244 26930 11296 26936
rect 11152 26852 11204 26858
rect 11152 26794 11204 26800
rect 11244 26580 11296 26586
rect 11244 26522 11296 26528
rect 11072 26438 11192 26466
rect 10968 25968 11020 25974
rect 10968 25910 11020 25916
rect 10980 25498 11008 25910
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 10784 25356 10836 25362
rect 10888 25350 11008 25378
rect 10784 25298 10836 25304
rect 10796 24886 10824 25298
rect 10876 25152 10928 25158
rect 10876 25094 10928 25100
rect 10888 24954 10916 25094
rect 10876 24948 10928 24954
rect 10876 24890 10928 24896
rect 10692 24880 10744 24886
rect 10692 24822 10744 24828
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10600 24608 10652 24614
rect 10600 24550 10652 24556
rect 10612 24342 10640 24550
rect 10704 24410 10732 24822
rect 10980 24750 11008 25350
rect 11060 25288 11112 25294
rect 11060 25230 11112 25236
rect 10784 24744 10836 24750
rect 10784 24686 10836 24692
rect 10968 24744 11020 24750
rect 10968 24686 11020 24692
rect 10796 24410 10824 24686
rect 11072 24682 11100 25230
rect 11164 25226 11192 26438
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 11060 24676 11112 24682
rect 11060 24618 11112 24624
rect 10692 24404 10744 24410
rect 10692 24346 10744 24352
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 10600 24336 10652 24342
rect 10600 24278 10652 24284
rect 10796 24206 10824 24346
rect 11164 24274 11192 25162
rect 11256 24614 11284 26522
rect 11348 25906 11376 31078
rect 11808 30938 11836 31078
rect 11900 30938 11928 31622
rect 11796 30932 11848 30938
rect 11796 30874 11848 30880
rect 11888 30932 11940 30938
rect 11888 30874 11940 30880
rect 12360 30326 12388 31826
rect 12912 31346 12940 33544
rect 14200 31940 14228 33544
rect 14306 32124 14614 32133
rect 14306 32122 14312 32124
rect 14368 32122 14392 32124
rect 14448 32122 14472 32124
rect 14528 32122 14552 32124
rect 14608 32122 14614 32124
rect 14368 32070 14370 32122
rect 14550 32070 14552 32122
rect 14306 32068 14312 32070
rect 14368 32068 14392 32070
rect 14448 32068 14472 32070
rect 14528 32068 14552 32070
rect 14608 32068 14614 32070
rect 14306 32059 14614 32068
rect 16132 31958 16160 33544
rect 17420 32026 17448 33544
rect 17776 32292 17828 32298
rect 17776 32234 17828 32240
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 14372 31952 14424 31958
rect 14200 31912 14372 31940
rect 14372 31894 14424 31900
rect 16120 31952 16172 31958
rect 16120 31894 16172 31900
rect 15384 31884 15436 31890
rect 15384 31826 15436 31832
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 14096 31816 14148 31822
rect 14096 31758 14148 31764
rect 13646 31580 13954 31589
rect 13646 31578 13652 31580
rect 13708 31578 13732 31580
rect 13788 31578 13812 31580
rect 13868 31578 13892 31580
rect 13948 31578 13954 31580
rect 13708 31526 13710 31578
rect 13890 31526 13892 31578
rect 13646 31524 13652 31526
rect 13708 31524 13732 31526
rect 13788 31524 13812 31526
rect 13868 31524 13892 31526
rect 13948 31524 13954 31526
rect 13646 31515 13954 31524
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 12440 31272 12492 31278
rect 12440 31214 12492 31220
rect 12452 30802 12480 31214
rect 12440 30796 12492 30802
rect 12440 30738 12492 30744
rect 12624 30796 12676 30802
rect 12624 30738 12676 30744
rect 12348 30320 12400 30326
rect 12348 30262 12400 30268
rect 11980 30184 12032 30190
rect 11980 30126 12032 30132
rect 11888 30048 11940 30054
rect 11888 29990 11940 29996
rect 11612 29640 11664 29646
rect 11612 29582 11664 29588
rect 11624 29238 11652 29582
rect 11612 29232 11664 29238
rect 11612 29174 11664 29180
rect 11900 29170 11928 29990
rect 11992 29850 12020 30126
rect 12360 29850 12388 30262
rect 11980 29844 12032 29850
rect 11980 29786 12032 29792
rect 12348 29844 12400 29850
rect 12348 29786 12400 29792
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 11888 29164 11940 29170
rect 11888 29106 11940 29112
rect 11796 29096 11848 29102
rect 11796 29038 11848 29044
rect 11612 27940 11664 27946
rect 11612 27882 11664 27888
rect 11428 27872 11480 27878
rect 11428 27814 11480 27820
rect 11440 27130 11468 27814
rect 11624 27674 11652 27882
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11808 27402 11836 29038
rect 12084 28218 12112 29514
rect 12532 29096 12584 29102
rect 12532 29038 12584 29044
rect 12440 29028 12492 29034
rect 12440 28970 12492 28976
rect 12072 28212 12124 28218
rect 12072 28154 12124 28160
rect 12452 27606 12480 28970
rect 12544 28762 12572 29038
rect 12532 28756 12584 28762
rect 12532 28698 12584 28704
rect 12440 27600 12492 27606
rect 12440 27542 12492 27548
rect 12164 27532 12216 27538
rect 12164 27474 12216 27480
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 11440 26450 11468 27066
rect 12176 26518 12204 27474
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 12360 26858 12388 27338
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 12440 26852 12492 26858
rect 12440 26794 12492 26800
rect 12164 26512 12216 26518
rect 12164 26454 12216 26460
rect 11428 26444 11480 26450
rect 11428 26386 11480 26392
rect 11612 26444 11664 26450
rect 11612 26386 11664 26392
rect 11520 26240 11572 26246
rect 11520 26182 11572 26188
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 11348 25809 11376 25842
rect 11334 25800 11390 25809
rect 11334 25735 11390 25744
rect 11428 25696 11480 25702
rect 11428 25638 11480 25644
rect 11440 25430 11468 25638
rect 11428 25424 11480 25430
rect 11348 25384 11428 25412
rect 11244 24608 11296 24614
rect 11244 24550 11296 24556
rect 11152 24268 11204 24274
rect 10980 24228 11152 24256
rect 10784 24200 10836 24206
rect 10836 24148 10916 24154
rect 10784 24142 10916 24148
rect 10796 24126 10916 24142
rect 10692 23520 10744 23526
rect 10692 23462 10744 23468
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10704 19310 10732 23462
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10796 21078 10824 22374
rect 10888 22030 10916 24126
rect 10980 23118 11008 24228
rect 11152 24210 11204 24216
rect 11244 24268 11296 24274
rect 11244 24210 11296 24216
rect 11058 24168 11114 24177
rect 11058 24103 11114 24112
rect 11072 23866 11100 24103
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11152 23860 11204 23866
rect 11152 23802 11204 23808
rect 11060 23316 11112 23322
rect 11060 23258 11112 23264
rect 10968 23112 11020 23118
rect 10968 23054 11020 23060
rect 11072 22522 11100 23258
rect 10980 22494 11100 22522
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10784 21072 10836 21078
rect 10784 21014 10836 21020
rect 10888 20466 10916 21966
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10508 19304 10560 19310
rect 10508 19246 10560 19252
rect 10692 19304 10744 19310
rect 10692 19246 10744 19252
rect 10520 18630 10548 19246
rect 10980 18834 11008 22494
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22234 11100 22374
rect 11060 22228 11112 22234
rect 11060 22170 11112 22176
rect 11072 21146 11100 22170
rect 11060 21140 11112 21146
rect 11060 21082 11112 21088
rect 11164 20602 11192 23802
rect 11256 22094 11284 24210
rect 11348 23866 11376 25384
rect 11428 25366 11480 25372
rect 11532 25294 11560 26182
rect 11624 26042 11652 26386
rect 11888 26240 11940 26246
rect 11888 26182 11940 26188
rect 11612 26036 11664 26042
rect 11612 25978 11664 25984
rect 11900 25498 11928 26182
rect 11612 25492 11664 25498
rect 11612 25434 11664 25440
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11520 25288 11572 25294
rect 11520 25230 11572 25236
rect 11428 24744 11480 24750
rect 11428 24686 11480 24692
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11440 23866 11468 24686
rect 11532 24274 11560 24686
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11520 24064 11572 24070
rect 11520 24006 11572 24012
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11348 23254 11376 23666
rect 11336 23248 11388 23254
rect 11336 23190 11388 23196
rect 11256 22066 11468 22094
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 11072 19922 11100 20266
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11348 19786 11376 21626
rect 11336 19780 11388 19786
rect 11336 19722 11388 19728
rect 11440 19174 11468 22066
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 10968 18828 11020 18834
rect 10968 18770 11020 18776
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10520 17814 10548 18566
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10508 17808 10560 17814
rect 10508 17750 10560 17756
rect 10612 17338 10640 18158
rect 10980 18154 11008 18770
rect 10968 18148 11020 18154
rect 10968 18090 11020 18096
rect 10600 17332 10652 17338
rect 10600 17274 10652 17280
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10980 16794 11008 17070
rect 10968 16788 11020 16794
rect 10968 16730 11020 16736
rect 10966 16688 11022 16697
rect 10966 16623 10968 16632
rect 11020 16623 11022 16632
rect 10968 16594 11020 16600
rect 10414 16552 10470 16561
rect 10414 16487 10416 16496
rect 10468 16487 10470 16496
rect 10416 16458 10468 16464
rect 10428 15978 10456 16458
rect 10980 16046 11008 16594
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10416 15972 10468 15978
rect 10416 15914 10468 15920
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10704 15366 10732 15846
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10968 15360 11020 15366
rect 10968 15302 11020 15308
rect 10704 15026 10732 15302
rect 10876 15088 10928 15094
rect 10876 15030 10928 15036
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10324 14612 10376 14618
rect 10324 14554 10376 14560
rect 10704 14278 10732 14962
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10232 14272 10284 14278
rect 10232 14214 10284 14220
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 11150 10088 12174
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10152 10674 10180 10950
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9600 5234 9628 5646
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9692 4826 9720 5034
rect 10244 4826 10272 14214
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10428 13530 10456 13738
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10428 12986 10456 13466
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10520 11694 10548 12174
rect 10612 11898 10640 13806
rect 10796 12782 10824 14758
rect 10888 14414 10916 15030
rect 10876 14408 10928 14414
rect 10876 14350 10928 14356
rect 10888 13938 10916 14350
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10980 13326 11008 15302
rect 11072 14074 11100 15506
rect 11164 14618 11192 15506
rect 11348 14958 11376 19110
rect 11532 18086 11560 24006
rect 11624 23769 11652 25434
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 11610 23760 11666 23769
rect 11610 23695 11666 23704
rect 11716 22574 11744 24890
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11900 24750 11928 24822
rect 11888 24744 11940 24750
rect 11888 24686 11940 24692
rect 12254 24712 12310 24721
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 11808 24177 11836 24550
rect 11794 24168 11850 24177
rect 11794 24103 11850 24112
rect 11900 23594 11928 24686
rect 12254 24647 12256 24656
rect 12308 24647 12310 24656
rect 12256 24618 12308 24624
rect 12256 24064 12308 24070
rect 12256 24006 12308 24012
rect 12268 23730 12296 24006
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 11888 23588 11940 23594
rect 11888 23530 11940 23536
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11704 22568 11756 22574
rect 11704 22510 11756 22516
rect 11624 21146 11652 22510
rect 11900 22420 11928 23530
rect 11992 22522 12020 23598
rect 12162 22536 12218 22545
rect 11992 22494 12112 22522
rect 11716 22392 11928 22420
rect 11980 22432 12032 22438
rect 11612 21140 11664 21146
rect 11612 21082 11664 21088
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11624 20058 11652 20538
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11610 19952 11666 19961
rect 11610 19887 11666 19896
rect 11624 19786 11652 19887
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11532 17542 11560 18022
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11532 16590 11560 17002
rect 11624 16658 11652 19722
rect 11716 17338 11744 22392
rect 11980 22374 12032 22380
rect 11992 22234 12020 22374
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 11796 22160 11848 22166
rect 11796 22102 11848 22108
rect 11808 21690 11836 22102
rect 12084 22094 12112 22494
rect 12162 22471 12218 22480
rect 11992 22066 12112 22094
rect 11992 22030 12020 22066
rect 11980 22024 12032 22030
rect 11980 21966 12032 21972
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 12084 21350 12112 22066
rect 12072 21344 12124 21350
rect 12072 21286 12124 21292
rect 11980 21072 12032 21078
rect 11980 21014 12032 21020
rect 11992 20466 12020 21014
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11704 17332 11756 17338
rect 11704 17274 11756 17280
rect 11716 16658 11744 17274
rect 11612 16652 11664 16658
rect 11612 16594 11664 16600
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11532 15910 11560 16526
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11336 14952 11388 14958
rect 11520 14952 11572 14958
rect 11336 14894 11388 14900
rect 11518 14920 11520 14929
rect 11572 14920 11574 14929
rect 11518 14855 11574 14864
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11152 14612 11204 14618
rect 11152 14554 11204 14560
rect 11152 14476 11204 14482
rect 11256 14464 11284 14758
rect 11348 14550 11376 14758
rect 11336 14544 11388 14550
rect 11336 14486 11388 14492
rect 11624 14498 11652 16594
rect 11808 15502 11836 19246
rect 11888 19236 11940 19242
rect 11888 19178 11940 19184
rect 11900 18426 11928 19178
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11900 17882 11928 18362
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11992 17678 12020 19110
rect 12084 18834 12112 21286
rect 12176 19310 12204 22471
rect 12256 20936 12308 20942
rect 12256 20878 12308 20884
rect 12268 20466 12296 20878
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 19922 12296 20402
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 17672 12032 17678
rect 11900 17632 11980 17660
rect 11900 16046 11928 17632
rect 11980 17614 12032 17620
rect 12084 17610 12112 18022
rect 12360 17626 12388 26794
rect 12452 26586 12480 26794
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12544 26234 12572 27406
rect 12636 26790 12664 30738
rect 13544 30728 13596 30734
rect 13544 30670 13596 30676
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 12912 30122 12940 30534
rect 12900 30116 12952 30122
rect 12900 30058 12952 30064
rect 13556 29850 13584 30670
rect 13646 30492 13954 30501
rect 13646 30490 13652 30492
rect 13708 30490 13732 30492
rect 13788 30490 13812 30492
rect 13868 30490 13892 30492
rect 13948 30490 13954 30492
rect 13708 30438 13710 30490
rect 13890 30438 13892 30490
rect 13646 30436 13652 30438
rect 13708 30436 13732 30438
rect 13788 30436 13812 30438
rect 13868 30436 13892 30438
rect 13948 30436 13954 30438
rect 13646 30427 13954 30436
rect 14108 30138 14136 31758
rect 15016 31476 15068 31482
rect 15016 31418 15068 31424
rect 14554 31376 14610 31385
rect 14188 31340 14240 31346
rect 14554 31311 14556 31320
rect 14188 31282 14240 31288
rect 14608 31311 14610 31320
rect 14556 31282 14608 31288
rect 14200 30258 14228 31282
rect 14306 31036 14614 31045
rect 14306 31034 14312 31036
rect 14368 31034 14392 31036
rect 14448 31034 14472 31036
rect 14528 31034 14552 31036
rect 14608 31034 14614 31036
rect 14368 30982 14370 31034
rect 14550 30982 14552 31034
rect 14306 30980 14312 30982
rect 14368 30980 14392 30982
rect 14448 30980 14472 30982
rect 14528 30980 14552 30982
rect 14608 30980 14614 30982
rect 14306 30971 14614 30980
rect 15028 30666 15056 31418
rect 15108 31136 15160 31142
rect 15108 31078 15160 31084
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15016 30660 15068 30666
rect 15016 30602 15068 30608
rect 14280 30592 14332 30598
rect 14280 30534 14332 30540
rect 14292 30258 14320 30534
rect 14188 30252 14240 30258
rect 14188 30194 14240 30200
rect 14280 30252 14332 30258
rect 14280 30194 14332 30200
rect 14740 30252 14792 30258
rect 14740 30194 14792 30200
rect 14752 30138 14780 30194
rect 14108 30110 14780 30138
rect 13544 29844 13596 29850
rect 13544 29786 13596 29792
rect 14108 29646 14136 30110
rect 14306 29948 14614 29957
rect 14306 29946 14312 29948
rect 14368 29946 14392 29948
rect 14448 29946 14472 29948
rect 14528 29946 14552 29948
rect 14608 29946 14614 29948
rect 14368 29894 14370 29946
rect 14550 29894 14552 29946
rect 14306 29892 14312 29894
rect 14368 29892 14392 29894
rect 14448 29892 14472 29894
rect 14528 29892 14552 29894
rect 14608 29892 14614 29894
rect 14306 29883 14614 29892
rect 15028 29850 15056 30602
rect 15120 30190 15148 31078
rect 15304 30870 15332 31078
rect 15292 30864 15344 30870
rect 15292 30806 15344 30812
rect 15200 30592 15252 30598
rect 15200 30534 15252 30540
rect 15212 30258 15240 30534
rect 15200 30252 15252 30258
rect 15200 30194 15252 30200
rect 15108 30184 15160 30190
rect 15108 30126 15160 30132
rect 15212 29850 15240 30194
rect 15016 29844 15068 29850
rect 15016 29786 15068 29792
rect 15200 29844 15252 29850
rect 15200 29786 15252 29792
rect 15108 29776 15160 29782
rect 15108 29718 15160 29724
rect 14832 29708 14884 29714
rect 14832 29650 14884 29656
rect 13636 29640 13688 29646
rect 13556 29588 13636 29594
rect 13556 29582 13688 29588
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14740 29640 14792 29646
rect 14740 29582 14792 29588
rect 13556 29566 13676 29582
rect 13452 29504 13504 29510
rect 13452 29446 13504 29452
rect 13360 29096 13412 29102
rect 13360 29038 13412 29044
rect 12900 28620 12952 28626
rect 12900 28562 12952 28568
rect 12912 28218 12940 28562
rect 13372 28218 13400 29038
rect 12900 28212 12952 28218
rect 12900 28154 12952 28160
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13464 27606 13492 29446
rect 13556 29034 13584 29566
rect 13646 29404 13954 29413
rect 13646 29402 13652 29404
rect 13708 29402 13732 29404
rect 13788 29402 13812 29404
rect 13868 29402 13892 29404
rect 13948 29402 13954 29404
rect 13708 29350 13710 29402
rect 13890 29350 13892 29402
rect 13646 29348 13652 29350
rect 13708 29348 13732 29350
rect 13788 29348 13812 29350
rect 13868 29348 13892 29350
rect 13948 29348 13954 29350
rect 13646 29339 13954 29348
rect 14108 29170 14136 29582
rect 14372 29504 14424 29510
rect 14372 29446 14424 29452
rect 14384 29306 14412 29446
rect 14372 29300 14424 29306
rect 14372 29242 14424 29248
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14188 29096 14240 29102
rect 14188 29038 14240 29044
rect 13544 29028 13596 29034
rect 13544 28970 13596 28976
rect 14096 28960 14148 28966
rect 14096 28902 14148 28908
rect 14004 28552 14056 28558
rect 14004 28494 14056 28500
rect 13646 28316 13954 28325
rect 13646 28314 13652 28316
rect 13708 28314 13732 28316
rect 13788 28314 13812 28316
rect 13868 28314 13892 28316
rect 13948 28314 13954 28316
rect 13708 28262 13710 28314
rect 13890 28262 13892 28314
rect 13646 28260 13652 28262
rect 13708 28260 13732 28262
rect 13788 28260 13812 28262
rect 13868 28260 13892 28262
rect 13948 28260 13954 28262
rect 13646 28251 13954 28260
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13452 27600 13504 27606
rect 13452 27542 13504 27548
rect 12624 26784 12676 26790
rect 12624 26726 12676 26732
rect 12636 26450 12664 26726
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12452 26206 12572 26234
rect 12452 24410 12480 26206
rect 13280 25906 13308 26454
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 12808 25832 12860 25838
rect 12808 25774 12860 25780
rect 12820 25498 12848 25774
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 13188 25498 13216 25706
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 13280 24818 13308 25842
rect 13268 24812 13320 24818
rect 13268 24754 13320 24760
rect 12992 24676 13044 24682
rect 12992 24618 13044 24624
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12452 22642 12480 24346
rect 12624 24268 12676 24274
rect 12624 24210 12676 24216
rect 12636 23118 12664 24210
rect 13004 23866 13032 24618
rect 13280 24342 13308 24754
rect 13372 24410 13400 26318
rect 13452 26240 13504 26246
rect 13452 26182 13504 26188
rect 13464 25362 13492 26182
rect 13556 25430 13584 27950
rect 14016 27946 14044 28494
rect 14108 28082 14136 28902
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 14016 27674 14044 27882
rect 14004 27668 14056 27674
rect 14004 27610 14056 27616
rect 14200 27334 14228 29038
rect 14648 28960 14700 28966
rect 14648 28902 14700 28908
rect 14306 28860 14614 28869
rect 14306 28858 14312 28860
rect 14368 28858 14392 28860
rect 14448 28858 14472 28860
rect 14528 28858 14552 28860
rect 14608 28858 14614 28860
rect 14368 28806 14370 28858
rect 14550 28806 14552 28858
rect 14306 28804 14312 28806
rect 14368 28804 14392 28806
rect 14448 28804 14472 28806
rect 14528 28804 14552 28806
rect 14608 28804 14614 28806
rect 14306 28795 14614 28804
rect 14660 28762 14688 28902
rect 14648 28756 14700 28762
rect 14648 28698 14700 28704
rect 14648 28416 14700 28422
rect 14752 28404 14780 29582
rect 14700 28376 14780 28404
rect 14648 28358 14700 28364
rect 14306 27772 14614 27781
rect 14306 27770 14312 27772
rect 14368 27770 14392 27772
rect 14448 27770 14472 27772
rect 14528 27770 14552 27772
rect 14608 27770 14614 27772
rect 14368 27718 14370 27770
rect 14550 27718 14552 27770
rect 14306 27716 14312 27718
rect 14368 27716 14392 27718
rect 14448 27716 14472 27718
rect 14528 27716 14552 27718
rect 14608 27716 14614 27718
rect 14306 27707 14614 27716
rect 14660 27656 14688 28358
rect 14384 27628 14688 27656
rect 14740 27668 14792 27674
rect 14384 27470 14412 27628
rect 14740 27610 14792 27616
rect 14464 27532 14516 27538
rect 14516 27492 14688 27520
rect 14464 27474 14516 27480
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 13646 27228 13954 27237
rect 13646 27226 13652 27228
rect 13708 27226 13732 27228
rect 13788 27226 13812 27228
rect 13868 27226 13892 27228
rect 13948 27226 13954 27228
rect 13708 27174 13710 27226
rect 13890 27174 13892 27226
rect 13646 27172 13652 27174
rect 13708 27172 13732 27174
rect 13788 27172 13812 27174
rect 13868 27172 13892 27174
rect 13948 27172 13954 27174
rect 13646 27163 13954 27172
rect 14384 26994 14412 27406
rect 14372 26988 14424 26994
rect 14372 26930 14424 26936
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 13646 26140 13954 26149
rect 13646 26138 13652 26140
rect 13708 26138 13732 26140
rect 13788 26138 13812 26140
rect 13868 26138 13892 26140
rect 13948 26138 13954 26140
rect 13708 26086 13710 26138
rect 13890 26086 13892 26138
rect 13646 26084 13652 26086
rect 13708 26084 13732 26086
rect 13788 26084 13812 26086
rect 13868 26084 13892 26086
rect 13948 26084 13954 26086
rect 13646 26075 13954 26084
rect 14108 25702 14136 26862
rect 14306 26684 14614 26693
rect 14306 26682 14312 26684
rect 14368 26682 14392 26684
rect 14448 26682 14472 26684
rect 14528 26682 14552 26684
rect 14608 26682 14614 26684
rect 14368 26630 14370 26682
rect 14550 26630 14552 26682
rect 14306 26628 14312 26630
rect 14368 26628 14392 26630
rect 14448 26628 14472 26630
rect 14528 26628 14552 26630
rect 14608 26628 14614 26630
rect 14306 26619 14614 26628
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14096 25696 14148 25702
rect 14016 25644 14096 25650
rect 14016 25638 14148 25644
rect 14016 25622 14136 25638
rect 13544 25424 13596 25430
rect 13544 25366 13596 25372
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 14016 25158 14044 25622
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13646 25052 13954 25061
rect 13646 25050 13652 25052
rect 13708 25050 13732 25052
rect 13788 25050 13812 25052
rect 13868 25050 13892 25052
rect 13948 25050 13954 25052
rect 13708 24998 13710 25050
rect 13890 24998 13892 25050
rect 13646 24996 13652 24998
rect 13708 24996 13732 24998
rect 13788 24996 13812 24998
rect 13868 24996 13892 24998
rect 13948 24996 13954 24998
rect 13646 24987 13954 24996
rect 14108 24818 14136 25230
rect 14096 24812 14148 24818
rect 14096 24754 14148 24760
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 14004 24744 14056 24750
rect 14004 24686 14056 24692
rect 13360 24404 13412 24410
rect 13360 24346 13412 24352
rect 13268 24336 13320 24342
rect 13268 24278 13320 24284
rect 13924 24206 13952 24686
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13646 23964 13954 23973
rect 13646 23962 13652 23964
rect 13708 23962 13732 23964
rect 13788 23962 13812 23964
rect 13868 23962 13892 23964
rect 13948 23962 13954 23964
rect 13708 23910 13710 23962
rect 13890 23910 13892 23962
rect 13646 23908 13652 23910
rect 13708 23908 13732 23910
rect 13788 23908 13812 23910
rect 13868 23908 13892 23910
rect 13948 23908 13954 23910
rect 13646 23899 13954 23908
rect 14016 23866 14044 24686
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13452 23520 13504 23526
rect 13452 23462 13504 23468
rect 13464 23168 13492 23462
rect 13556 23322 13584 23598
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13544 23180 13596 23186
rect 13464 23140 13544 23168
rect 13544 23122 13596 23128
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12624 23112 12676 23118
rect 13556 23089 13584 23122
rect 12624 23054 12676 23060
rect 13542 23080 13598 23089
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12544 22438 12572 23054
rect 13268 23044 13320 23050
rect 13452 23044 13504 23050
rect 13320 23004 13452 23032
rect 13268 22986 13320 22992
rect 13924 23066 13952 23734
rect 14108 23254 14136 24754
rect 14096 23248 14148 23254
rect 14096 23190 14148 23196
rect 13924 23038 14136 23066
rect 13542 23015 13598 23024
rect 13452 22986 13504 22992
rect 13544 22976 13596 22982
rect 13544 22918 13596 22924
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 13360 22568 13412 22574
rect 13360 22510 13412 22516
rect 12624 22500 12676 22506
rect 12624 22442 12676 22448
rect 12532 22432 12584 22438
rect 12532 22374 12584 22380
rect 12440 21072 12492 21078
rect 12440 21014 12492 21020
rect 12452 20466 12480 21014
rect 12636 20874 12664 22442
rect 12820 21690 12848 22510
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12808 21684 12860 21690
rect 12808 21626 12860 21632
rect 12912 21418 12940 21830
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 13280 21010 13308 22374
rect 13372 22234 13400 22510
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13464 22234 13492 22374
rect 13556 22234 13584 22918
rect 13646 22876 13954 22885
rect 13646 22874 13652 22876
rect 13708 22874 13732 22876
rect 13788 22874 13812 22876
rect 13868 22874 13892 22876
rect 13948 22874 13954 22876
rect 13708 22822 13710 22874
rect 13890 22822 13892 22874
rect 13646 22820 13652 22822
rect 13708 22820 13732 22822
rect 13788 22820 13812 22822
rect 13868 22820 13892 22822
rect 13948 22820 13954 22822
rect 13646 22811 13954 22820
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13452 22228 13504 22234
rect 13452 22170 13504 22176
rect 13544 22228 13596 22234
rect 13544 22170 13596 22176
rect 13464 21536 13492 22170
rect 13372 21508 13492 21536
rect 13372 21078 13400 21508
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 13360 21072 13412 21078
rect 13360 21014 13412 21020
rect 13268 21004 13320 21010
rect 13268 20946 13320 20952
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12624 20868 12676 20874
rect 12624 20810 12676 20816
rect 12440 20460 12492 20466
rect 12440 20402 12492 20408
rect 12636 20398 12664 20810
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12624 20392 12676 20398
rect 12624 20334 12676 20340
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 12532 19304 12584 19310
rect 12532 19246 12584 19252
rect 12544 18902 12572 19246
rect 12532 18896 12584 18902
rect 12532 18838 12584 18844
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 17746 12480 18566
rect 12544 18154 12572 18838
rect 12636 18766 12664 19722
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12532 18148 12584 18154
rect 12532 18090 12584 18096
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12636 17882 12664 18090
rect 12728 18086 12756 20198
rect 12820 19922 12848 20742
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12820 18970 12848 19178
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12912 18834 12940 19858
rect 13004 19825 13032 20878
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 12990 19816 13046 19825
rect 12990 19751 13046 19760
rect 13096 19417 13124 20198
rect 13188 19910 13400 19938
rect 13082 19408 13138 19417
rect 13082 19343 13138 19352
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 13004 18426 13032 18702
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 13096 18154 13124 18566
rect 13084 18148 13136 18154
rect 13084 18090 13136 18096
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12728 17882 12756 18022
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 12176 17598 12388 17626
rect 12176 17354 12204 17598
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 12084 17326 12204 17354
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11796 15496 11848 15502
rect 11796 15438 11848 15444
rect 11796 15360 11848 15366
rect 11796 15302 11848 15308
rect 11808 15065 11836 15302
rect 11794 15056 11850 15065
rect 11794 14991 11850 15000
rect 11808 14958 11836 14991
rect 11796 14952 11848 14958
rect 11796 14894 11848 14900
rect 11900 14890 11928 15982
rect 11992 15366 12020 16934
rect 12084 16522 12112 17326
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12176 16522 12204 17138
rect 12360 17134 12388 17478
rect 13004 17338 13032 18022
rect 13188 17814 13216 19910
rect 13372 19854 13400 19910
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13280 17814 13308 19790
rect 13464 18902 13492 21354
rect 13556 21078 13584 22170
rect 14004 21888 14056 21894
rect 14004 21830 14056 21836
rect 13646 21788 13954 21797
rect 13646 21786 13652 21788
rect 13708 21786 13732 21788
rect 13788 21786 13812 21788
rect 13868 21786 13892 21788
rect 13948 21786 13954 21788
rect 13708 21734 13710 21786
rect 13890 21734 13892 21786
rect 13646 21732 13652 21734
rect 13708 21732 13732 21734
rect 13788 21732 13812 21734
rect 13868 21732 13892 21734
rect 13948 21732 13954 21734
rect 13646 21723 13954 21732
rect 14016 21690 14044 21830
rect 14004 21684 14056 21690
rect 14004 21626 14056 21632
rect 14004 21412 14056 21418
rect 14004 21354 14056 21360
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13556 20262 13584 21014
rect 14016 21010 14044 21354
rect 14108 21146 14136 23038
rect 14200 22778 14228 26318
rect 14660 26314 14688 27492
rect 14752 27470 14780 27610
rect 14740 27464 14792 27470
rect 14740 27406 14792 27412
rect 14752 26518 14780 27406
rect 14844 26586 14872 29650
rect 14924 27600 14976 27606
rect 14924 27542 14976 27548
rect 14936 26926 14964 27542
rect 15016 27464 15068 27470
rect 15016 27406 15068 27412
rect 15028 27130 15056 27406
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 14924 26920 14976 26926
rect 14924 26862 14976 26868
rect 14924 26784 14976 26790
rect 14924 26726 14976 26732
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14740 26512 14792 26518
rect 14740 26454 14792 26460
rect 14648 26308 14700 26314
rect 14648 26250 14700 26256
rect 14306 25596 14614 25605
rect 14306 25594 14312 25596
rect 14368 25594 14392 25596
rect 14448 25594 14472 25596
rect 14528 25594 14552 25596
rect 14608 25594 14614 25596
rect 14368 25542 14370 25594
rect 14550 25542 14552 25594
rect 14306 25540 14312 25542
rect 14368 25540 14392 25542
rect 14448 25540 14472 25542
rect 14528 25540 14552 25542
rect 14608 25540 14614 25542
rect 14306 25531 14614 25540
rect 14660 25412 14688 26250
rect 14740 25832 14792 25838
rect 14740 25774 14792 25780
rect 14752 25498 14780 25774
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14292 25384 14688 25412
rect 14292 24954 14320 25384
rect 14740 25356 14792 25362
rect 14740 25298 14792 25304
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14648 25288 14700 25294
rect 14648 25230 14700 25236
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14476 24886 14504 25230
rect 14556 25152 14608 25158
rect 14556 25094 14608 25100
rect 14568 24954 14596 25094
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14464 24880 14516 24886
rect 14464 24822 14516 24828
rect 14306 24508 14614 24517
rect 14306 24506 14312 24508
rect 14368 24506 14392 24508
rect 14448 24506 14472 24508
rect 14528 24506 14552 24508
rect 14608 24506 14614 24508
rect 14368 24454 14370 24506
rect 14550 24454 14552 24506
rect 14306 24452 14312 24454
rect 14368 24452 14392 24454
rect 14448 24452 14472 24454
rect 14528 24452 14552 24454
rect 14608 24452 14614 24454
rect 14306 24443 14614 24452
rect 14660 24392 14688 25230
rect 14752 24426 14780 25298
rect 14844 24614 14872 26522
rect 14936 24954 14964 26726
rect 15120 26353 15148 29718
rect 15396 29050 15424 31826
rect 16592 31770 16620 31826
rect 16592 31742 16712 31770
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 15936 31136 15988 31142
rect 15936 31078 15988 31084
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 15948 30054 15976 31078
rect 16040 30870 16068 31078
rect 16028 30864 16080 30870
rect 16028 30806 16080 30812
rect 16592 30394 16620 31214
rect 16580 30388 16632 30394
rect 16580 30330 16632 30336
rect 16684 30274 16712 31742
rect 17500 31136 17552 31142
rect 17500 31078 17552 31084
rect 16948 30864 17000 30870
rect 16948 30806 17000 30812
rect 16960 30394 16988 30806
rect 17316 30660 17368 30666
rect 17316 30602 17368 30608
rect 17040 30592 17092 30598
rect 17040 30534 17092 30540
rect 16948 30388 17000 30394
rect 16948 30330 17000 30336
rect 16684 30246 16988 30274
rect 16304 30116 16356 30122
rect 16304 30058 16356 30064
rect 15936 30048 15988 30054
rect 15936 29990 15988 29996
rect 15752 29640 15804 29646
rect 15752 29582 15804 29588
rect 15304 29022 15424 29050
rect 15200 26920 15252 26926
rect 15200 26862 15252 26868
rect 15212 26586 15240 26862
rect 15200 26580 15252 26586
rect 15200 26522 15252 26528
rect 15106 26344 15162 26353
rect 15106 26279 15162 26288
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 15120 25770 15148 26182
rect 15304 25906 15332 29022
rect 15764 28762 15792 29582
rect 15948 28966 15976 29990
rect 16316 29714 16344 30058
rect 16304 29708 16356 29714
rect 16304 29650 16356 29656
rect 16580 29640 16632 29646
rect 16580 29582 16632 29588
rect 16120 29096 16172 29102
rect 16120 29038 16172 29044
rect 15844 28960 15896 28966
rect 15844 28902 15896 28908
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 15856 28694 15884 28902
rect 15844 28688 15896 28694
rect 15844 28630 15896 28636
rect 15948 28626 15976 28902
rect 15936 28620 15988 28626
rect 15936 28562 15988 28568
rect 15948 28082 15976 28562
rect 16028 28416 16080 28422
rect 16028 28358 16080 28364
rect 15936 28076 15988 28082
rect 15936 28018 15988 28024
rect 16040 27606 16068 28358
rect 16132 28218 16160 29038
rect 16592 28422 16620 29582
rect 16856 29504 16908 29510
rect 16856 29446 16908 29452
rect 16868 29034 16896 29446
rect 16856 29028 16908 29034
rect 16856 28970 16908 28976
rect 16212 28416 16264 28422
rect 16212 28358 16264 28364
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16224 28014 16252 28358
rect 16592 28121 16620 28358
rect 16578 28112 16634 28121
rect 16578 28047 16634 28056
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16304 27872 16356 27878
rect 16304 27814 16356 27820
rect 16028 27600 16080 27606
rect 16028 27542 16080 27548
rect 16316 27538 16344 27814
rect 16304 27532 16356 27538
rect 16304 27474 16356 27480
rect 16764 27532 16816 27538
rect 16764 27474 16816 27480
rect 16672 26784 16724 26790
rect 16672 26726 16724 26732
rect 15384 26580 15436 26586
rect 15384 26522 15436 26528
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15108 25764 15160 25770
rect 15108 25706 15160 25712
rect 15396 25158 15424 26522
rect 16684 26382 16712 26726
rect 16672 26376 16724 26382
rect 16672 26318 16724 26324
rect 16776 26330 16804 27474
rect 16868 27334 16896 28970
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 15568 26308 15620 26314
rect 16776 26302 16896 26330
rect 15568 26250 15620 26256
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15488 25498 15516 25638
rect 15476 25492 15528 25498
rect 15476 25434 15528 25440
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 14832 24608 14884 24614
rect 14832 24550 14884 24556
rect 14752 24398 14872 24426
rect 14476 24364 14688 24392
rect 14372 24336 14424 24342
rect 14372 24278 14424 24284
rect 14384 23866 14412 24278
rect 14476 24206 14504 24364
rect 14740 24336 14792 24342
rect 14740 24278 14792 24284
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 14476 23594 14504 24142
rect 14648 23656 14700 23662
rect 14648 23598 14700 23604
rect 14464 23588 14516 23594
rect 14464 23530 14516 23536
rect 14660 23526 14688 23598
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14306 23420 14614 23429
rect 14306 23418 14312 23420
rect 14368 23418 14392 23420
rect 14448 23418 14472 23420
rect 14528 23418 14552 23420
rect 14608 23418 14614 23420
rect 14368 23366 14370 23418
rect 14550 23366 14552 23418
rect 14306 23364 14312 23366
rect 14368 23364 14392 23366
rect 14448 23364 14472 23366
rect 14528 23364 14552 23366
rect 14608 23364 14614 23366
rect 14306 23355 14614 23364
rect 14370 23216 14426 23225
rect 14280 23180 14332 23186
rect 14370 23151 14372 23160
rect 14280 23122 14332 23128
rect 14424 23151 14426 23160
rect 14372 23122 14424 23128
rect 14292 22982 14320 23122
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14188 22772 14240 22778
rect 14188 22714 14240 22720
rect 14384 22710 14412 23122
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14372 22704 14424 22710
rect 14372 22646 14424 22652
rect 14476 22545 14504 22714
rect 14660 22658 14688 23462
rect 14752 23322 14780 24278
rect 14844 23730 14872 24398
rect 14936 24070 14964 24890
rect 15108 24880 15160 24886
rect 15108 24822 15160 24828
rect 14924 24064 14976 24070
rect 14924 24006 14976 24012
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 15120 23610 15148 24822
rect 15198 24168 15254 24177
rect 15198 24103 15254 24112
rect 15212 23798 15240 24103
rect 15292 24064 15344 24070
rect 15292 24006 15344 24012
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15120 23582 15240 23610
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 14740 23044 14792 23050
rect 14740 22986 14792 22992
rect 14752 22778 14780 22986
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14568 22630 14688 22658
rect 14568 22574 14596 22630
rect 14556 22568 14608 22574
rect 14462 22536 14518 22545
rect 14556 22510 14608 22516
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14462 22471 14518 22480
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14200 21554 14228 22374
rect 14306 22332 14614 22341
rect 14306 22330 14312 22332
rect 14368 22330 14392 22332
rect 14448 22330 14472 22332
rect 14528 22330 14552 22332
rect 14608 22330 14614 22332
rect 14368 22278 14370 22330
rect 14550 22278 14552 22330
rect 14306 22276 14312 22278
rect 14368 22276 14392 22278
rect 14448 22276 14472 22278
rect 14528 22276 14552 22278
rect 14608 22276 14614 22278
rect 14306 22267 14614 22276
rect 14660 22166 14688 22374
rect 14648 22160 14700 22166
rect 14648 22102 14700 22108
rect 14660 21962 14688 22102
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14096 21140 14148 21146
rect 14096 21082 14148 21088
rect 14200 21010 14228 21490
rect 14306 21244 14614 21253
rect 14306 21242 14312 21244
rect 14368 21242 14392 21244
rect 14448 21242 14472 21244
rect 14528 21242 14552 21244
rect 14608 21242 14614 21244
rect 14368 21190 14370 21242
rect 14550 21190 14552 21242
rect 14306 21188 14312 21190
rect 14368 21188 14392 21190
rect 14448 21188 14472 21190
rect 14528 21188 14552 21190
rect 14608 21188 14614 21190
rect 14306 21179 14614 21188
rect 14004 21004 14056 21010
rect 14188 21004 14240 21010
rect 14056 20964 14136 20992
rect 14004 20946 14056 20952
rect 13820 20936 13872 20942
rect 13818 20904 13820 20913
rect 13872 20904 13874 20913
rect 13818 20839 13874 20848
rect 13646 20700 13954 20709
rect 13646 20698 13652 20700
rect 13708 20698 13732 20700
rect 13788 20698 13812 20700
rect 13868 20698 13892 20700
rect 13948 20698 13954 20700
rect 13708 20646 13710 20698
rect 13890 20646 13892 20698
rect 13646 20644 13652 20646
rect 13708 20644 13732 20646
rect 13788 20644 13812 20646
rect 13868 20644 13892 20646
rect 13948 20644 13954 20646
rect 13646 20635 13954 20644
rect 14108 20482 14136 20964
rect 14188 20946 14240 20952
rect 14464 21004 14516 21010
rect 14464 20946 14516 20952
rect 14200 20602 14228 20946
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14108 20454 14228 20482
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 14096 20256 14148 20262
rect 14096 20198 14148 20204
rect 14004 19712 14056 19718
rect 14004 19654 14056 19660
rect 13646 19612 13954 19621
rect 13646 19610 13652 19612
rect 13708 19610 13732 19612
rect 13788 19610 13812 19612
rect 13868 19610 13892 19612
rect 13948 19610 13954 19612
rect 13708 19558 13710 19610
rect 13890 19558 13892 19610
rect 13646 19556 13652 19558
rect 13708 19556 13732 19558
rect 13788 19556 13812 19558
rect 13868 19556 13892 19558
rect 13948 19556 13954 19558
rect 13646 19547 13954 19556
rect 13542 19408 13598 19417
rect 13542 19343 13598 19352
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13360 18828 13412 18834
rect 13360 18770 13412 18776
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13268 17808 13320 17814
rect 13268 17750 13320 17756
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13082 17232 13138 17241
rect 13082 17167 13138 17176
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12072 16516 12124 16522
rect 12072 16458 12124 16464
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12084 16114 12112 16458
rect 12176 16250 12204 16458
rect 12164 16244 12216 16250
rect 12164 16186 12216 16192
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11204 14436 11284 14464
rect 11152 14418 11204 14424
rect 11348 14396 11376 14486
rect 11428 14476 11480 14482
rect 11624 14470 11744 14498
rect 11428 14418 11480 14424
rect 11256 14368 11376 14396
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11256 13870 11284 14368
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11244 13864 11296 13870
rect 11244 13806 11296 13812
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10888 12306 10916 12786
rect 11072 12481 11100 13806
rect 11164 13462 11192 13806
rect 11348 13462 11376 13942
rect 11440 13734 11468 14418
rect 11612 14272 11664 14278
rect 11612 14214 11664 14220
rect 11428 13728 11480 13734
rect 11428 13670 11480 13676
rect 11152 13456 11204 13462
rect 11152 13398 11204 13404
rect 11336 13456 11388 13462
rect 11336 13398 11388 13404
rect 11624 12986 11652 14214
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11612 12776 11664 12782
rect 11612 12718 11664 12724
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11058 12472 11114 12481
rect 11058 12407 11114 12416
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 11072 11762 11100 12407
rect 11164 12374 11192 12582
rect 11624 12442 11652 12718
rect 11716 12646 11744 14470
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 13802 11836 14350
rect 11900 14278 11928 14826
rect 11992 14482 12020 15098
rect 11980 14476 12032 14482
rect 11980 14418 12032 14424
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11888 13796 11940 13802
rect 11888 13738 11940 13744
rect 11900 12986 11928 13738
rect 11992 13734 12020 14418
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 12084 12850 12112 16050
rect 12176 15638 12204 16186
rect 12268 15706 12296 17070
rect 12360 16182 12388 17070
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 12544 16454 12572 16487
rect 12636 16454 12664 16934
rect 12820 16658 12848 16934
rect 13096 16794 13124 17167
rect 13084 16788 13136 16794
rect 13084 16730 13136 16736
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 12544 16182 12572 16390
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 12636 16046 12664 16390
rect 13096 16250 13124 16730
rect 13188 16250 13216 17750
rect 13280 17338 13308 17750
rect 13372 17490 13400 18770
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13464 17610 13492 18702
rect 13556 17746 13584 19343
rect 14016 19224 14044 19654
rect 14108 19242 14136 20198
rect 14200 19514 14228 20454
rect 14476 20346 14504 20946
rect 14556 20800 14608 20806
rect 14556 20742 14608 20748
rect 14568 20602 14596 20742
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14660 20466 14688 21898
rect 14752 21894 14780 22510
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14752 20777 14780 21830
rect 14844 21690 14872 22918
rect 14936 22098 14964 23122
rect 15016 22704 15068 22710
rect 15016 22646 15068 22652
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 14924 21888 14976 21894
rect 15028 21876 15056 22646
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15120 22273 15148 22510
rect 15106 22264 15162 22273
rect 15106 22199 15162 22208
rect 15212 22098 15240 23582
rect 15304 23254 15332 24006
rect 15396 23662 15424 25094
rect 15580 24954 15608 26250
rect 15936 26240 15988 26246
rect 15936 26182 15988 26188
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 15948 25430 15976 26182
rect 16304 25832 16356 25838
rect 16304 25774 16356 25780
rect 15936 25424 15988 25430
rect 15936 25366 15988 25372
rect 16316 24954 16344 25774
rect 16488 25696 16540 25702
rect 16488 25638 16540 25644
rect 15568 24948 15620 24954
rect 15568 24890 15620 24896
rect 16304 24948 16356 24954
rect 16304 24890 16356 24896
rect 16500 24750 16528 25638
rect 16776 25430 16804 26182
rect 16764 25424 16816 25430
rect 16764 25366 16816 25372
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16212 24608 16264 24614
rect 16212 24550 16264 24556
rect 15844 24268 15896 24274
rect 15844 24210 15896 24216
rect 15856 23866 15884 24210
rect 16028 24132 16080 24138
rect 16028 24074 16080 24080
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15660 23792 15712 23798
rect 15660 23734 15712 23740
rect 15384 23656 15436 23662
rect 15384 23598 15436 23604
rect 15476 23520 15528 23526
rect 15476 23462 15528 23468
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 15292 23248 15344 23254
rect 15292 23190 15344 23196
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15396 22098 15424 22918
rect 15488 22506 15516 23462
rect 15580 22574 15608 23462
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15476 22500 15528 22506
rect 15476 22442 15528 22448
rect 15200 22092 15252 22098
rect 15200 22034 15252 22040
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 14976 21848 15056 21876
rect 15292 21888 15344 21894
rect 14924 21830 14976 21836
rect 15292 21830 15344 21836
rect 14832 21684 14884 21690
rect 14832 21626 14884 21632
rect 14936 20890 14964 21830
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15028 21010 15056 21286
rect 15120 21146 15148 21422
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 14936 20862 15056 20890
rect 14924 20800 14976 20806
rect 14738 20768 14794 20777
rect 14924 20742 14976 20748
rect 14738 20703 14794 20712
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14740 20392 14792 20398
rect 14476 20340 14740 20346
rect 14476 20334 14792 20340
rect 14476 20318 14780 20334
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14306 20156 14614 20165
rect 14306 20154 14312 20156
rect 14368 20154 14392 20156
rect 14448 20154 14472 20156
rect 14528 20154 14552 20156
rect 14608 20154 14614 20156
rect 14368 20102 14370 20154
rect 14550 20102 14552 20154
rect 14306 20100 14312 20102
rect 14368 20100 14392 20102
rect 14448 20100 14472 20102
rect 14528 20100 14552 20102
rect 14608 20100 14614 20102
rect 14306 20091 14614 20100
rect 14660 20040 14688 20198
rect 14752 20058 14780 20198
rect 14568 20012 14688 20040
rect 14740 20052 14792 20058
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14188 19508 14240 19514
rect 14188 19450 14240 19456
rect 13832 19196 14044 19224
rect 14096 19236 14148 19242
rect 13832 18970 13860 19196
rect 14096 19178 14148 19184
rect 14292 19156 14320 19926
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 14200 19128 14320 19156
rect 14476 19156 14504 19314
rect 14568 19281 14596 20012
rect 14740 19994 14792 20000
rect 14740 19916 14792 19922
rect 14792 19876 14872 19904
rect 14740 19858 14792 19864
rect 14740 19780 14792 19786
rect 14740 19722 14792 19728
rect 14752 19417 14780 19722
rect 14738 19408 14794 19417
rect 14738 19343 14794 19352
rect 14740 19304 14792 19310
rect 14554 19272 14610 19281
rect 14554 19207 14610 19216
rect 14738 19272 14740 19281
rect 14792 19272 14794 19281
rect 14738 19207 14794 19216
rect 14728 19168 14780 19174
rect 14476 19128 14688 19156
rect 14200 19122 14228 19128
rect 14108 19094 14228 19122
rect 14108 18970 14136 19094
rect 14306 19068 14614 19077
rect 14306 19066 14312 19068
rect 14368 19066 14392 19068
rect 14448 19066 14472 19068
rect 14528 19066 14552 19068
rect 14608 19066 14614 19068
rect 14368 19014 14370 19066
rect 14550 19014 14552 19066
rect 14306 19012 14312 19014
rect 14368 19012 14392 19014
rect 14448 19012 14472 19014
rect 14528 19012 14552 19014
rect 14608 19012 14614 19014
rect 14306 19003 14614 19012
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14096 18964 14148 18970
rect 14556 18964 14608 18970
rect 14096 18906 14148 18912
rect 14200 18924 14556 18952
rect 14200 18834 14228 18924
rect 14556 18906 14608 18912
rect 14370 18864 14426 18873
rect 14188 18828 14240 18834
rect 14370 18799 14426 18808
rect 14188 18770 14240 18776
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 13646 18524 13954 18533
rect 13646 18522 13652 18524
rect 13708 18522 13732 18524
rect 13788 18522 13812 18524
rect 13868 18522 13892 18524
rect 13948 18522 13954 18524
rect 13708 18470 13710 18522
rect 13890 18470 13892 18522
rect 13646 18468 13652 18470
rect 13708 18468 13732 18470
rect 13788 18468 13812 18470
rect 13868 18468 13892 18470
rect 13948 18468 13954 18470
rect 13646 18459 13954 18468
rect 14002 17776 14058 17785
rect 13544 17740 13596 17746
rect 14002 17711 14058 17720
rect 13544 17682 13596 17688
rect 14016 17678 14044 17711
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 13452 17604 13504 17610
rect 13452 17546 13504 17552
rect 14108 17542 14136 18566
rect 14200 17796 14228 18770
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14292 18170 14320 18634
rect 14384 18426 14412 18799
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14660 18222 14688 19128
rect 14728 19110 14780 19116
rect 14740 18970 14768 19110
rect 14740 18964 14792 18970
rect 14740 18906 14792 18912
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14648 18216 14700 18222
rect 14370 18184 14426 18193
rect 14292 18142 14370 18170
rect 14648 18158 14700 18164
rect 14370 18119 14426 18128
rect 14306 17980 14614 17989
rect 14306 17978 14312 17980
rect 14368 17978 14392 17980
rect 14448 17978 14472 17980
rect 14528 17978 14552 17980
rect 14608 17978 14614 17980
rect 14368 17926 14370 17978
rect 14550 17926 14552 17978
rect 14306 17924 14312 17926
rect 14368 17924 14392 17926
rect 14448 17924 14472 17926
rect 14528 17924 14552 17926
rect 14608 17924 14614 17926
rect 14306 17915 14614 17924
rect 14648 17808 14700 17814
rect 14200 17768 14320 17796
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 13544 17536 13596 17542
rect 13372 17462 13492 17490
rect 13544 17478 13596 17484
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 13268 17332 13320 17338
rect 13268 17274 13320 17280
rect 13360 17128 13412 17134
rect 13358 17096 13360 17105
rect 13464 17116 13492 17462
rect 13556 17338 13584 17478
rect 13646 17436 13954 17445
rect 13646 17434 13652 17436
rect 13708 17434 13732 17436
rect 13788 17434 13812 17436
rect 13868 17434 13892 17436
rect 13948 17434 13954 17436
rect 13708 17382 13710 17434
rect 13890 17382 13892 17434
rect 13646 17380 13652 17382
rect 13708 17380 13732 17382
rect 13788 17380 13812 17382
rect 13868 17380 13892 17382
rect 13948 17380 13954 17382
rect 13646 17371 13954 17380
rect 14016 17338 14044 17478
rect 14094 17368 14150 17377
rect 13544 17332 13596 17338
rect 13544 17274 13596 17280
rect 14004 17332 14056 17338
rect 14094 17303 14150 17312
rect 14004 17274 14056 17280
rect 13544 17128 13596 17134
rect 13412 17096 13414 17105
rect 13358 17031 13414 17040
rect 13464 17088 13544 17116
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12624 16040 12676 16046
rect 12624 15982 12676 15988
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12360 15706 12388 15846
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12176 12714 12204 15302
rect 12360 14822 12388 15506
rect 12348 14816 12400 14822
rect 12348 14758 12400 14764
rect 12254 14240 12310 14249
rect 12254 14175 12310 14184
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 12268 12374 12296 14175
rect 12360 12918 12388 14758
rect 12452 14074 12480 15982
rect 13188 15706 13216 16186
rect 13372 16046 13400 16594
rect 13464 16114 13492 17088
rect 13544 17070 13596 17076
rect 14004 17128 14056 17134
rect 14004 17070 14056 17076
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13452 16108 13504 16114
rect 13452 16050 13504 16056
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13556 15978 13584 16934
rect 14016 16726 14044 17070
rect 14108 16794 14136 17303
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13646 16348 13954 16357
rect 13646 16346 13652 16348
rect 13708 16346 13732 16348
rect 13788 16346 13812 16348
rect 13868 16346 13892 16348
rect 13948 16346 13954 16348
rect 13708 16294 13710 16346
rect 13890 16294 13892 16346
rect 13646 16292 13652 16294
rect 13708 16292 13732 16294
rect 13788 16292 13812 16294
rect 13868 16292 13892 16294
rect 13948 16292 13954 16294
rect 13646 16283 13954 16292
rect 14108 16232 14136 16730
rect 14200 16250 14228 17614
rect 14292 17202 14320 17768
rect 14648 17750 14700 17756
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14384 17338 14412 17478
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14292 16980 14320 17138
rect 14476 17134 14504 17478
rect 14554 17368 14610 17377
rect 14554 17303 14610 17312
rect 14568 17270 14596 17303
rect 14556 17264 14608 17270
rect 14556 17206 14608 17212
rect 14660 17184 14688 17750
rect 14752 17746 14780 18362
rect 14844 17882 14872 19876
rect 14936 19854 14964 20742
rect 14924 19848 14976 19854
rect 14924 19790 14976 19796
rect 15028 19334 15056 20862
rect 15212 20466 15240 21626
rect 15304 21486 15332 21830
rect 15292 21480 15344 21486
rect 15292 21422 15344 21428
rect 15304 21185 15332 21422
rect 15290 21176 15346 21185
rect 15290 21111 15346 21120
rect 15304 20602 15332 21111
rect 15396 20602 15424 22034
rect 15488 21486 15516 22442
rect 15580 22234 15608 22510
rect 15568 22228 15620 22234
rect 15568 22170 15620 22176
rect 15568 22024 15620 22030
rect 15568 21966 15620 21972
rect 15580 21622 15608 21966
rect 15568 21616 15620 21622
rect 15568 21558 15620 21564
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15672 21350 15700 23734
rect 15752 23588 15804 23594
rect 15752 23530 15804 23536
rect 15764 23118 15792 23530
rect 16040 23526 16068 24074
rect 16132 23769 16160 24550
rect 16224 24070 16252 24550
rect 16212 24064 16264 24070
rect 16212 24006 16264 24012
rect 16118 23760 16174 23769
rect 16118 23695 16174 23704
rect 16132 23662 16160 23695
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16028 23520 16080 23526
rect 16028 23462 16080 23468
rect 15844 23248 15896 23254
rect 15844 23190 15896 23196
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15764 22420 15792 23054
rect 15856 22710 15884 23190
rect 16120 23112 16172 23118
rect 16120 23054 16172 23060
rect 16132 22778 16160 23054
rect 16120 22772 16172 22778
rect 16120 22714 16172 22720
rect 15844 22704 15896 22710
rect 15844 22646 15896 22652
rect 15844 22432 15896 22438
rect 15764 22392 15844 22420
rect 15764 22030 15792 22392
rect 15844 22374 15896 22380
rect 16500 22392 16620 22420
rect 16394 22264 16450 22273
rect 16500 22234 16528 22392
rect 16394 22199 16450 22208
rect 16488 22228 16540 22234
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15672 21010 15700 21286
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 14936 19306 15056 19334
rect 14936 18170 14964 19306
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 15028 18834 15056 19110
rect 15016 18828 15068 18834
rect 15016 18770 15068 18776
rect 15120 18329 15148 19994
rect 15198 19952 15254 19961
rect 15198 19887 15254 19896
rect 15212 19854 15240 19887
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15292 19712 15344 19718
rect 15292 19654 15344 19660
rect 15200 19236 15252 19242
rect 15200 19178 15252 19184
rect 15212 18834 15240 19178
rect 15304 19174 15332 19654
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15304 18970 15332 19110
rect 15292 18964 15344 18970
rect 15292 18906 15344 18912
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15106 18320 15162 18329
rect 15106 18255 15162 18264
rect 14936 18142 15056 18170
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14740 17740 14792 17746
rect 14740 17682 14792 17688
rect 14660 17156 14780 17184
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14292 16952 14688 16980
rect 14306 16892 14614 16901
rect 14306 16890 14312 16892
rect 14368 16890 14392 16892
rect 14448 16890 14472 16892
rect 14528 16890 14552 16892
rect 14608 16890 14614 16892
rect 14368 16838 14370 16890
rect 14550 16838 14552 16890
rect 14306 16836 14312 16838
rect 14368 16836 14392 16838
rect 14448 16836 14472 16838
rect 14528 16836 14552 16838
rect 14608 16836 14614 16838
rect 14306 16827 14614 16836
rect 13832 16204 14136 16232
rect 14188 16244 14240 16250
rect 13544 15972 13596 15978
rect 13544 15914 13596 15920
rect 13176 15700 13228 15706
rect 13004 15660 13176 15688
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 15026 12572 15438
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12544 13326 12572 14962
rect 12636 14482 12664 15506
rect 12820 15162 12848 15506
rect 12912 15162 12940 15506
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12808 14816 12860 14822
rect 12806 14784 12808 14793
rect 12860 14784 12862 14793
rect 12806 14719 12862 14728
rect 12912 14618 12940 15098
rect 13004 15094 13032 15660
rect 13176 15642 13228 15648
rect 13268 15632 13320 15638
rect 13268 15574 13320 15580
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 13096 14822 13124 14894
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13280 14618 13308 15574
rect 13832 15348 13860 16204
rect 14188 16186 14240 16192
rect 14094 16144 14150 16153
rect 14016 16102 14094 16130
rect 14016 16046 14044 16102
rect 14094 16079 14150 16088
rect 14004 16040 14056 16046
rect 14004 15982 14056 15988
rect 14016 15570 14044 15982
rect 14200 15706 14228 16186
rect 14660 16114 14688 16952
rect 14648 16108 14700 16114
rect 14648 16050 14700 16056
rect 14648 15972 14700 15978
rect 14648 15914 14700 15920
rect 14306 15804 14614 15813
rect 14306 15802 14312 15804
rect 14368 15802 14392 15804
rect 14448 15802 14472 15804
rect 14528 15802 14552 15804
rect 14608 15802 14614 15804
rect 14368 15750 14370 15802
rect 14550 15750 14552 15802
rect 14306 15748 14312 15750
rect 14368 15748 14392 15750
rect 14448 15748 14472 15750
rect 14528 15748 14552 15750
rect 14608 15748 14614 15750
rect 14306 15739 14614 15748
rect 14660 15706 14688 15914
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14004 15564 14056 15570
rect 14004 15506 14056 15512
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 13556 15320 13860 15348
rect 14004 15360 14056 15366
rect 13452 15156 13504 15162
rect 13452 15098 13504 15104
rect 13358 15056 13414 15065
rect 13358 14991 13414 15000
rect 13372 14958 13400 14991
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13358 14784 13414 14793
rect 13358 14719 13414 14728
rect 13372 14618 13400 14719
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13464 14482 13492 15098
rect 13556 15042 13584 15320
rect 14004 15302 14056 15308
rect 13646 15260 13954 15269
rect 13646 15258 13652 15260
rect 13708 15258 13732 15260
rect 13788 15258 13812 15260
rect 13868 15258 13892 15260
rect 13948 15258 13954 15260
rect 13708 15206 13710 15258
rect 13890 15206 13892 15258
rect 13646 15204 13652 15206
rect 13708 15204 13732 15206
rect 13788 15204 13812 15206
rect 13868 15204 13892 15206
rect 13948 15204 13954 15206
rect 13646 15195 13954 15204
rect 13556 15014 13952 15042
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13096 14074 13124 14418
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13556 13870 13584 14758
rect 13924 14328 13952 15014
rect 14016 14618 14044 15302
rect 14108 14929 14136 15506
rect 14200 15366 14228 15506
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14094 14920 14150 14929
rect 14094 14855 14150 14864
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 14108 14414 14136 14855
rect 14200 14532 14228 15302
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14306 14716 14614 14725
rect 14306 14714 14312 14716
rect 14368 14714 14392 14716
rect 14448 14714 14472 14716
rect 14528 14714 14552 14716
rect 14608 14714 14614 14716
rect 14368 14662 14370 14714
rect 14550 14662 14552 14714
rect 14306 14660 14312 14662
rect 14368 14660 14392 14662
rect 14448 14660 14472 14662
rect 14528 14660 14552 14662
rect 14608 14660 14614 14662
rect 14306 14651 14614 14660
rect 14660 14618 14688 14894
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14200 14504 14320 14532
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 13924 14300 14044 14328
rect 13646 14172 13954 14181
rect 13646 14170 13652 14172
rect 13708 14170 13732 14172
rect 13788 14170 13812 14172
rect 13868 14170 13892 14172
rect 13948 14170 13954 14172
rect 13708 14118 13710 14170
rect 13890 14118 13892 14170
rect 13646 14116 13652 14118
rect 13708 14116 13732 14118
rect 13788 14116 13812 14118
rect 13868 14116 13892 14118
rect 13948 14116 13954 14118
rect 13646 14107 13954 14116
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 12624 13796 12676 13802
rect 12624 13738 12676 13744
rect 12636 13462 12664 13738
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12348 12912 12400 12918
rect 12348 12854 12400 12860
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 11152 12368 11204 12374
rect 11150 12336 11152 12345
rect 11704 12368 11756 12374
rect 11204 12336 11206 12345
rect 12256 12368 12308 12374
rect 11704 12310 11756 12316
rect 12084 12328 12256 12356
rect 11150 12271 11206 12280
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 11716 11626 11744 12310
rect 12084 11694 12112 12328
rect 12256 12310 12308 12316
rect 12072 11688 12124 11694
rect 11900 11648 12072 11676
rect 11704 11620 11756 11626
rect 11704 11562 11756 11568
rect 10600 11552 10652 11558
rect 10600 11494 10652 11500
rect 10612 11286 10640 11494
rect 10416 11280 10468 11286
rect 10416 11222 10468 11228
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10428 10674 10456 11222
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 10416 10668 10468 10674
rect 10416 10610 10468 10616
rect 10520 10266 10548 11086
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11532 10470 11560 10950
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10874 9072 10930 9081
rect 10874 9007 10876 9016
rect 10928 9007 10930 9016
rect 10876 8978 10928 8984
rect 10416 5772 10468 5778
rect 10416 5714 10468 5720
rect 10428 5030 10456 5714
rect 10416 5024 10468 5030
rect 10416 4966 10468 4972
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 10428 3602 10456 4966
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10324 3528 10376 3534
rect 10324 3470 10376 3476
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 5816 2916 5868 2922
rect 5816 2858 5868 2864
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 5828 800 5856 2858
rect 6946 2748 7254 2757
rect 6946 2746 6952 2748
rect 7008 2746 7032 2748
rect 7088 2746 7112 2748
rect 7168 2746 7192 2748
rect 7248 2746 7254 2748
rect 7008 2694 7010 2746
rect 7190 2694 7192 2746
rect 6946 2692 6952 2694
rect 7008 2692 7032 2694
rect 7088 2692 7112 2694
rect 7168 2692 7192 2694
rect 7248 2692 7254 2694
rect 6946 2683 7254 2692
rect 7300 1442 7328 2858
rect 7116 1414 7328 1442
rect 7116 800 7144 1414
rect 9048 800 9076 2858
rect 10336 800 10364 3470
rect 11532 2990 11560 10406
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11624 6254 11652 8910
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11716 3942 11744 8910
rect 11900 6866 11928 11648
rect 12072 11630 12124 11636
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12072 11552 12124 11558
rect 12072 11494 12124 11500
rect 12084 11286 12112 11494
rect 12268 11354 12296 11630
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11354 12388 11494
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12452 11082 12480 12378
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12636 12102 12664 12174
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12636 11150 12664 12038
rect 12912 11762 12940 13330
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13004 12442 13032 12786
rect 13188 12714 13216 12922
rect 13556 12918 13584 13806
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 13924 13530 13952 13670
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 14016 13258 14044 14300
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 13802 14136 14214
rect 14292 14006 14320 14504
rect 14648 14476 14700 14482
rect 14752 14464 14780 17156
rect 14844 16998 14872 17818
rect 14936 17134 14964 18022
rect 15028 17814 15056 18142
rect 15016 17808 15068 17814
rect 15016 17750 15068 17756
rect 15014 17368 15070 17377
rect 15014 17303 15070 17312
rect 15028 17202 15056 17303
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15120 17134 15148 18255
rect 15290 17232 15346 17241
rect 15396 17218 15424 20334
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15672 19990 15700 20198
rect 15476 19984 15528 19990
rect 15660 19984 15712 19990
rect 15476 19926 15528 19932
rect 15658 19952 15660 19961
rect 15712 19952 15714 19961
rect 15488 19718 15516 19926
rect 15568 19916 15620 19922
rect 15658 19887 15714 19896
rect 15568 19858 15620 19864
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15488 18426 15516 18702
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15476 17604 15528 17610
rect 15476 17546 15528 17552
rect 15346 17190 15424 17218
rect 15290 17167 15346 17176
rect 14924 17128 14976 17134
rect 14924 17070 14976 17076
rect 15108 17128 15160 17134
rect 15108 17070 15160 17076
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 15292 16992 15344 16998
rect 15292 16934 15344 16940
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 14844 16794 14872 16934
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 15028 16250 15056 16934
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15016 16244 15068 16250
rect 15068 16204 15148 16232
rect 15016 16186 15068 16192
rect 15016 15904 15068 15910
rect 15016 15846 15068 15852
rect 14832 15564 14884 15570
rect 14832 15506 14884 15512
rect 14844 14958 14872 15506
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14936 14804 14964 14894
rect 14700 14436 14780 14464
rect 14844 14776 14964 14804
rect 14648 14418 14700 14424
rect 14556 14408 14608 14414
rect 14608 14356 14780 14362
rect 14556 14350 14780 14356
rect 14568 14334 14780 14350
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 14200 13462 14228 13874
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14292 13734 14320 13806
rect 14280 13728 14332 13734
rect 14280 13670 14332 13676
rect 14306 13628 14614 13637
rect 14306 13626 14312 13628
rect 14368 13626 14392 13628
rect 14448 13626 14472 13628
rect 14528 13626 14552 13628
rect 14608 13626 14614 13628
rect 14368 13574 14370 13626
rect 14550 13574 14552 13626
rect 14306 13572 14312 13574
rect 14368 13572 14392 13574
rect 14448 13572 14472 13574
rect 14528 13572 14552 13574
rect 14608 13572 14614 13574
rect 14306 13563 14614 13572
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14096 13388 14148 13394
rect 14096 13330 14148 13336
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 13646 13084 13954 13093
rect 13646 13082 13652 13084
rect 13708 13082 13732 13084
rect 13788 13082 13812 13084
rect 13868 13082 13892 13084
rect 13948 13082 13954 13084
rect 13708 13030 13710 13082
rect 13890 13030 13892 13082
rect 13646 13028 13652 13030
rect 13708 13028 13732 13030
rect 13788 13028 13812 13030
rect 13868 13028 13892 13030
rect 13948 13028 13954 13030
rect 13646 13019 13954 13028
rect 13544 12912 13596 12918
rect 13464 12872 13544 12900
rect 13176 12708 13228 12714
rect 13176 12650 13228 12656
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 12900 11756 12952 11762
rect 12900 11698 12952 11704
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12440 11076 12492 11082
rect 12440 11018 12492 11024
rect 12452 10266 12480 11018
rect 13004 10810 13032 11494
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12544 6934 12572 10610
rect 13096 10606 13124 12174
rect 13188 10810 13216 12650
rect 13464 11234 13492 12872
rect 13544 12854 13596 12860
rect 14004 12708 14056 12714
rect 14004 12650 14056 12656
rect 13646 11996 13954 12005
rect 13646 11994 13652 11996
rect 13708 11994 13732 11996
rect 13788 11994 13812 11996
rect 13868 11994 13892 11996
rect 13948 11994 13954 11996
rect 13708 11942 13710 11994
rect 13890 11942 13892 11994
rect 13646 11940 13652 11942
rect 13708 11940 13732 11942
rect 13788 11940 13812 11942
rect 13868 11940 13892 11942
rect 13948 11940 13954 11942
rect 13646 11931 13954 11940
rect 14016 11694 14044 12650
rect 14108 12374 14136 13330
rect 14200 12850 14228 13398
rect 14556 13388 14608 13394
rect 14556 13330 14608 13336
rect 14568 12986 14596 13330
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14660 12714 14688 14010
rect 14752 13394 14780 14334
rect 14844 14278 14872 14776
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14844 14074 14872 14214
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14936 13870 14964 14214
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14936 13462 14964 13806
rect 15028 13802 15056 15846
rect 15120 14074 15148 16204
rect 15212 15502 15240 16594
rect 15304 16114 15332 16934
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15304 15706 15332 16050
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15396 15570 15424 16934
rect 15488 16250 15516 17546
rect 15580 16794 15608 19858
rect 15764 19242 15792 21966
rect 16132 21690 16160 21966
rect 16120 21684 16172 21690
rect 16120 21626 16172 21632
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 15844 21480 15896 21486
rect 15896 21440 15976 21468
rect 15844 21422 15896 21428
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 15752 19236 15804 19242
rect 15752 19178 15804 19184
rect 15856 19122 15884 21286
rect 15948 21078 15976 21440
rect 16028 21412 16080 21418
rect 16028 21354 16080 21360
rect 15936 21072 15988 21078
rect 15936 21014 15988 21020
rect 15948 20398 15976 21014
rect 16040 20777 16068 21354
rect 16026 20768 16082 20777
rect 16026 20703 16082 20712
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15934 19952 15990 19961
rect 15934 19887 15990 19896
rect 15672 19094 15884 19122
rect 15672 17678 15700 19094
rect 15752 18896 15804 18902
rect 15752 18838 15804 18844
rect 15764 18408 15792 18838
rect 15844 18420 15896 18426
rect 15764 18380 15844 18408
rect 15844 18362 15896 18368
rect 15842 18320 15898 18329
rect 15842 18255 15898 18264
rect 15750 18184 15806 18193
rect 15856 18154 15884 18255
rect 15750 18119 15806 18128
rect 15844 18148 15896 18154
rect 15764 18086 15792 18119
rect 15844 18090 15896 18096
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15764 17746 15792 18022
rect 15752 17740 15804 17746
rect 15752 17682 15804 17688
rect 15660 17672 15712 17678
rect 15660 17614 15712 17620
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15672 16697 15700 17614
rect 15764 17202 15792 17682
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15948 17082 15976 19887
rect 16224 19802 16252 21558
rect 16408 21418 16436 22199
rect 16488 22170 16540 22176
rect 16592 21434 16620 22392
rect 16592 21418 16712 21434
rect 16396 21412 16448 21418
rect 16592 21412 16724 21418
rect 16592 21406 16672 21412
rect 16396 21354 16448 21360
rect 16672 21354 16724 21360
rect 16580 21344 16632 21350
rect 16580 21286 16632 21292
rect 16592 20534 16620 21286
rect 16670 21176 16726 21185
rect 16670 21111 16726 21120
rect 16684 20806 16712 21111
rect 16868 21078 16896 26302
rect 16960 26234 16988 30246
rect 17052 30190 17080 30534
rect 17328 30394 17356 30602
rect 17316 30388 17368 30394
rect 17316 30330 17368 30336
rect 17512 30258 17540 31078
rect 17788 30666 17816 32234
rect 18708 32026 18736 33544
rect 17868 32020 17920 32026
rect 17868 31962 17920 31968
rect 18696 32020 18748 32026
rect 18696 31962 18748 31968
rect 18788 32020 18840 32026
rect 18788 31962 18840 31968
rect 18972 32020 19024 32026
rect 18972 31962 19024 31968
rect 17880 31793 17908 31962
rect 18800 31929 18828 31962
rect 18786 31920 18842 31929
rect 18786 31855 18842 31864
rect 17866 31784 17922 31793
rect 17866 31719 17922 31728
rect 18420 31680 18472 31686
rect 18420 31622 18472 31628
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17776 30660 17828 30666
rect 17776 30602 17828 30608
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17040 30184 17092 30190
rect 17040 30126 17092 30132
rect 17052 29102 17080 30126
rect 18064 29850 18092 31214
rect 18432 30734 18460 31622
rect 18604 31136 18656 31142
rect 18604 31078 18656 31084
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 18616 30598 18644 31078
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18604 30592 18656 30598
rect 18604 30534 18656 30540
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 18512 29708 18564 29714
rect 18512 29650 18564 29656
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 17040 29096 17092 29102
rect 17040 29038 17092 29044
rect 17052 28082 17080 29038
rect 17132 28552 17184 28558
rect 17132 28494 17184 28500
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 17052 26586 17080 28018
rect 17144 27470 17172 28494
rect 17788 28422 17816 29582
rect 18328 29504 18380 29510
rect 18328 29446 18380 29452
rect 18340 29306 18368 29446
rect 18328 29300 18380 29306
rect 18328 29242 18380 29248
rect 18524 29170 18552 29650
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 17776 28416 17828 28422
rect 17776 28358 17828 28364
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17144 26858 17172 27270
rect 17512 27130 17540 27474
rect 17500 27124 17552 27130
rect 17500 27066 17552 27072
rect 17316 26920 17368 26926
rect 17316 26862 17368 26868
rect 17132 26852 17184 26858
rect 17132 26794 17184 26800
rect 17040 26580 17092 26586
rect 17092 26540 17172 26568
rect 17040 26522 17092 26528
rect 16960 26206 17080 26234
rect 17052 25906 17080 26206
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17052 25498 17080 25842
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 17144 24818 17172 26540
rect 17328 26042 17356 26862
rect 17500 26784 17552 26790
rect 17500 26726 17552 26732
rect 17316 26036 17368 26042
rect 17316 25978 17368 25984
rect 17224 25832 17276 25838
rect 17224 25774 17276 25780
rect 17132 24812 17184 24818
rect 17132 24754 17184 24760
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 17144 24274 17172 24550
rect 17132 24268 17184 24274
rect 17132 24210 17184 24216
rect 16948 24064 17000 24070
rect 16948 24006 17000 24012
rect 16960 21486 16988 24006
rect 17040 23520 17092 23526
rect 17040 23462 17092 23468
rect 17052 22778 17080 23462
rect 17040 22772 17092 22778
rect 17040 22714 17092 22720
rect 17132 21616 17184 21622
rect 17132 21558 17184 21564
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 17144 21418 17172 21558
rect 17132 21412 17184 21418
rect 17132 21354 17184 21360
rect 17236 21350 17264 25774
rect 17512 25702 17540 26726
rect 17500 25696 17552 25702
rect 17500 25638 17552 25644
rect 17512 24614 17540 25638
rect 17604 25362 17632 27814
rect 17684 27532 17736 27538
rect 17684 27474 17736 27480
rect 17696 27334 17724 27474
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 17788 26994 17816 28358
rect 17960 27940 18012 27946
rect 17960 27882 18012 27888
rect 17972 27674 18000 27882
rect 17960 27668 18012 27674
rect 17960 27610 18012 27616
rect 17776 26988 17828 26994
rect 17776 26930 17828 26936
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18432 25906 18460 26318
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 18524 25702 18552 26182
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 17592 25356 17644 25362
rect 17592 25298 17644 25304
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18328 25152 18380 25158
rect 18328 25094 18380 25100
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 24206 17540 24550
rect 17500 24200 17552 24206
rect 17500 24142 17552 24148
rect 17972 24138 18000 24618
rect 18144 24336 18196 24342
rect 18144 24278 18196 24284
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17592 23656 17644 23662
rect 17592 23598 17644 23604
rect 17604 23322 17632 23598
rect 17592 23316 17644 23322
rect 17592 23258 17644 23264
rect 17880 23186 17908 23802
rect 17868 23180 17920 23186
rect 17868 23122 17920 23128
rect 18052 23112 18104 23118
rect 18156 23089 18184 24278
rect 18340 23866 18368 25094
rect 18432 23866 18460 25230
rect 18524 24954 18552 25638
rect 18512 24948 18564 24954
rect 18512 24890 18564 24896
rect 18328 23860 18380 23866
rect 18328 23802 18380 23808
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18328 23520 18380 23526
rect 18328 23462 18380 23468
rect 18052 23054 18104 23060
rect 18142 23080 18198 23089
rect 17960 22500 18012 22506
rect 17960 22442 18012 22448
rect 17972 22234 18000 22442
rect 17960 22228 18012 22234
rect 17960 22170 18012 22176
rect 18064 21962 18092 23054
rect 18142 23015 18198 23024
rect 18052 21956 18104 21962
rect 18052 21898 18104 21904
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 16856 21072 16908 21078
rect 16856 21014 16908 21020
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 16580 20528 16632 20534
rect 16580 20470 16632 20476
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16132 19774 16252 19802
rect 16132 19258 16160 19774
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16040 19230 16160 19258
rect 16040 19174 16068 19230
rect 16028 19168 16080 19174
rect 16028 19110 16080 19116
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16132 18630 16160 19110
rect 16120 18624 16172 18630
rect 16120 18566 16172 18572
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16040 17338 16068 18158
rect 16132 17746 16160 18566
rect 16224 18222 16252 19654
rect 16500 18698 16528 19994
rect 16764 19984 16816 19990
rect 16764 19926 16816 19932
rect 16776 19786 16804 19926
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16764 19780 16816 19786
rect 16764 19722 16816 19728
rect 16488 18692 16540 18698
rect 16488 18634 16540 18640
rect 16500 18358 16528 18634
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16212 18216 16264 18222
rect 16212 18158 16264 18164
rect 16488 18216 16540 18222
rect 16540 18176 16620 18204
rect 16488 18158 16540 18164
rect 16120 17740 16172 17746
rect 16120 17682 16172 17688
rect 16224 17338 16252 18158
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 16212 17332 16264 17338
rect 16316 17320 16344 17818
rect 16408 17814 16436 18022
rect 16486 17912 16542 17921
rect 16486 17847 16542 17856
rect 16396 17808 16448 17814
rect 16396 17750 16448 17756
rect 16500 17610 16528 17847
rect 16488 17604 16540 17610
rect 16488 17546 16540 17552
rect 16396 17332 16448 17338
rect 16316 17292 16396 17320
rect 16212 17274 16264 17280
rect 16396 17274 16448 17280
rect 16120 17264 16172 17270
rect 16120 17206 16172 17212
rect 15856 17054 15976 17082
rect 15658 16688 15714 16697
rect 15714 16646 15792 16674
rect 15658 16623 15714 16632
rect 15764 16590 15792 16646
rect 15752 16584 15804 16590
rect 15752 16526 15804 16532
rect 15568 16448 15620 16454
rect 15568 16390 15620 16396
rect 15660 16448 15712 16454
rect 15660 16390 15712 16396
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15488 16153 15516 16186
rect 15474 16144 15530 16153
rect 15474 16079 15530 16088
rect 15476 16040 15528 16046
rect 15476 15982 15528 15988
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15488 15366 15516 15982
rect 15580 15570 15608 16390
rect 15672 16046 15700 16390
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15660 15632 15712 15638
rect 15856 15586 15884 17054
rect 15936 16992 15988 16998
rect 15936 16934 15988 16940
rect 15948 16454 15976 16934
rect 16132 16454 16160 17206
rect 16224 16658 16252 17274
rect 16304 17196 16356 17202
rect 16500 17184 16528 17546
rect 16592 17490 16620 18176
rect 16684 17814 16712 19722
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16776 18630 16804 19246
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 16592 17462 16712 17490
rect 16304 17138 16356 17144
rect 16408 17156 16528 17184
rect 16212 16652 16264 16658
rect 16212 16594 16264 16600
rect 15936 16448 15988 16454
rect 15936 16390 15988 16396
rect 16120 16448 16172 16454
rect 16120 16390 16172 16396
rect 15660 15574 15712 15580
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15568 15428 15620 15434
rect 15568 15370 15620 15376
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15382 15192 15438 15201
rect 15382 15127 15384 15136
rect 15436 15127 15438 15136
rect 15384 15098 15436 15104
rect 15396 15042 15424 15098
rect 15304 15014 15424 15042
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 15120 13530 15148 14010
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14648 12708 14700 12714
rect 14648 12650 14700 12656
rect 14752 12594 14780 13194
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14660 12566 14780 12594
rect 14306 12540 14614 12549
rect 14306 12538 14312 12540
rect 14368 12538 14392 12540
rect 14448 12538 14472 12540
rect 14528 12538 14552 12540
rect 14608 12538 14614 12540
rect 14368 12486 14370 12538
rect 14550 12486 14552 12538
rect 14306 12484 14312 12486
rect 14368 12484 14392 12486
rect 14448 12484 14472 12486
rect 14528 12484 14552 12486
rect 14608 12484 14614 12486
rect 14306 12475 14614 12484
rect 14660 12374 14688 12566
rect 14096 12368 14148 12374
rect 14096 12310 14148 12316
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14108 11898 14136 12310
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 14004 11688 14056 11694
rect 14004 11630 14056 11636
rect 13556 11354 13584 11630
rect 14306 11452 14614 11461
rect 14306 11450 14312 11452
rect 14368 11450 14392 11452
rect 14448 11450 14472 11452
rect 14528 11450 14552 11452
rect 14608 11450 14614 11452
rect 14368 11398 14370 11450
rect 14550 11398 14552 11450
rect 14306 11396 14312 11398
rect 14368 11396 14392 11398
rect 14448 11396 14472 11398
rect 14528 11396 14552 11398
rect 14608 11396 14614 11398
rect 14306 11387 14614 11396
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 14002 11248 14058 11257
rect 13464 11206 13584 11234
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13464 10674 13492 11018
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13084 10600 13136 10606
rect 13084 10542 13136 10548
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12728 10130 12756 10406
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 13556 9382 13584 11206
rect 14002 11183 14004 11192
rect 14056 11183 14058 11192
rect 14004 11154 14056 11160
rect 14936 11150 14964 11698
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 13646 10908 13954 10917
rect 13646 10906 13652 10908
rect 13708 10906 13732 10908
rect 13788 10906 13812 10908
rect 13868 10906 13892 10908
rect 13948 10906 13954 10908
rect 13708 10854 13710 10906
rect 13890 10854 13892 10906
rect 13646 10852 13652 10854
rect 13708 10852 13732 10854
rect 13788 10852 13812 10854
rect 13868 10852 13892 10854
rect 13948 10852 13954 10854
rect 13646 10843 13954 10852
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13646 9820 13954 9829
rect 13646 9818 13652 9820
rect 13708 9818 13732 9820
rect 13788 9818 13812 9820
rect 13868 9818 13892 9820
rect 13948 9818 13954 9820
rect 13708 9766 13710 9818
rect 13890 9766 13892 9818
rect 13646 9764 13652 9766
rect 13708 9764 13732 9766
rect 13788 9764 13812 9766
rect 13868 9764 13892 9766
rect 13948 9764 13954 9766
rect 13646 9755 13954 9764
rect 14016 9636 14044 10746
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 14108 10266 14136 10474
rect 14306 10364 14614 10373
rect 14306 10362 14312 10364
rect 14368 10362 14392 10364
rect 14448 10362 14472 10364
rect 14528 10362 14552 10364
rect 14608 10362 14614 10364
rect 14368 10310 14370 10362
rect 14550 10310 14552 10362
rect 14306 10308 14312 10310
rect 14368 10308 14392 10310
rect 14448 10308 14472 10310
rect 14528 10308 14552 10310
rect 14608 10308 14614 10310
rect 14306 10299 14614 10308
rect 14096 10260 14148 10266
rect 14096 10202 14148 10208
rect 14660 10062 14688 10542
rect 14936 10266 14964 11086
rect 15028 10674 15056 12786
rect 15304 12238 15332 15014
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14550 15516 14894
rect 15476 14544 15528 14550
rect 15476 14486 15528 14492
rect 15580 14482 15608 15370
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15672 13870 15700 15574
rect 15764 15558 15884 15586
rect 16132 15570 16160 16390
rect 16316 15978 16344 17138
rect 16304 15972 16356 15978
rect 16304 15914 16356 15920
rect 16120 15564 16172 15570
rect 15764 14822 15792 15558
rect 16120 15506 16172 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 15026 15884 15438
rect 15844 15020 15896 15026
rect 15844 14962 15896 14968
rect 16132 14958 16160 15506
rect 16120 14952 16172 14958
rect 16040 14912 16120 14940
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15764 12374 15792 13126
rect 15384 12368 15436 12374
rect 15384 12310 15436 12316
rect 15752 12368 15804 12374
rect 15752 12310 15804 12316
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15396 11830 15424 12310
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15856 11694 15884 14486
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15948 13530 15976 14350
rect 15936 13524 15988 13530
rect 15936 13466 15988 13472
rect 16040 13394 16068 14912
rect 16120 14894 16172 14900
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16132 13394 16160 14758
rect 16028 13388 16080 13394
rect 16028 13330 16080 13336
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16224 12434 16252 14758
rect 16408 13818 16436 17156
rect 16580 17128 16632 17134
rect 16486 17096 16542 17105
rect 16580 17070 16632 17076
rect 16486 17031 16542 17040
rect 16500 16794 16528 17031
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16592 16658 16620 17070
rect 16684 16998 16712 17462
rect 16776 17134 16804 18566
rect 16868 18222 16896 19246
rect 16948 19168 17000 19174
rect 16948 19110 17000 19116
rect 16960 18902 16988 19110
rect 16948 18896 17000 18902
rect 16948 18838 17000 18844
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16856 18216 16908 18222
rect 16856 18158 16908 18164
rect 16856 18080 16908 18086
rect 16854 18048 16856 18057
rect 16908 18048 16910 18057
rect 16854 17983 16910 17992
rect 16960 17746 16988 18702
rect 17052 18170 17080 20742
rect 17408 19236 17460 19242
rect 17408 19178 17460 19184
rect 17420 18970 17448 19178
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17052 18142 17264 18170
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16856 17604 16908 17610
rect 16856 17546 16908 17552
rect 16764 17128 16816 17134
rect 16764 17070 16816 17076
rect 16672 16992 16724 16998
rect 16868 16946 16896 17546
rect 16672 16934 16724 16940
rect 16776 16918 16896 16946
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16684 16250 16712 16594
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16580 16040 16632 16046
rect 16580 15982 16632 15988
rect 16672 16040 16724 16046
rect 16672 15982 16724 15988
rect 16592 15502 16620 15982
rect 16684 15570 16712 15982
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16592 14890 16620 15438
rect 16776 14906 16804 16918
rect 16960 16522 16988 17682
rect 17052 17202 17080 18022
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 17144 17202 17172 17614
rect 17236 17610 17264 18142
rect 17316 18080 17368 18086
rect 17316 18022 17368 18028
rect 17406 18048 17462 18057
rect 17224 17604 17276 17610
rect 17224 17546 17276 17552
rect 17328 17542 17356 18022
rect 17406 17983 17462 17992
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17132 17196 17184 17202
rect 17132 17138 17184 17144
rect 17038 17096 17094 17105
rect 17038 17031 17040 17040
rect 17092 17031 17094 17040
rect 17040 17002 17092 17008
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 17144 16182 17172 17138
rect 17328 17134 17356 17478
rect 17316 17128 17368 17134
rect 17236 17088 17316 17116
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16868 15162 16896 16050
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17052 15638 17080 15846
rect 17040 15632 17092 15638
rect 17040 15574 17092 15580
rect 17236 15570 17264 17088
rect 17316 17070 17368 17076
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16590 17356 16934
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17420 16454 17448 17983
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17420 16250 17448 16390
rect 17408 16244 17460 16250
rect 17408 16186 17460 16192
rect 17512 15706 17540 21422
rect 17590 19816 17646 19825
rect 17590 19751 17646 19760
rect 17604 18970 17632 19751
rect 17684 19712 17736 19718
rect 17684 19654 17736 19660
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17592 17740 17644 17746
rect 17592 17682 17644 17688
rect 17604 17338 17632 17682
rect 17696 17610 17724 19654
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17788 18426 17816 18702
rect 17776 18420 17828 18426
rect 17776 18362 17828 18368
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17604 16726 17632 17070
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 17696 16250 17724 17546
rect 17880 17542 17908 18702
rect 17972 17678 18000 21830
rect 18064 21486 18092 21898
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 18064 19174 18092 21422
rect 18156 19854 18184 23015
rect 18236 22160 18288 22166
rect 18236 22102 18288 22108
rect 18248 21690 18276 22102
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18340 20942 18368 23462
rect 18420 21684 18472 21690
rect 18420 21626 18472 21632
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18432 19922 18460 21626
rect 18616 19961 18644 30534
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18708 29238 18736 29582
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18708 23322 18736 23598
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18800 23202 18828 30602
rect 18984 30326 19012 31962
rect 20640 31958 20668 33544
rect 21456 32360 21508 32366
rect 21456 32302 21508 32308
rect 21928 32314 21956 33544
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 19524 31748 19576 31754
rect 19524 31690 19576 31696
rect 19536 30802 19564 31690
rect 21006 31580 21314 31589
rect 21006 31578 21012 31580
rect 21068 31578 21092 31580
rect 21148 31578 21172 31580
rect 21228 31578 21252 31580
rect 21308 31578 21314 31580
rect 21068 31526 21070 31578
rect 21250 31526 21252 31578
rect 21006 31524 21012 31526
rect 21068 31524 21092 31526
rect 21148 31524 21172 31526
rect 21228 31524 21252 31526
rect 21308 31524 21314 31526
rect 21006 31515 21314 31524
rect 21364 31136 21416 31142
rect 21364 31078 21416 31084
rect 21376 30870 21404 31078
rect 21364 30864 21416 30870
rect 21364 30806 21416 30812
rect 19524 30796 19576 30802
rect 19524 30738 19576 30744
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20260 30592 20312 30598
rect 20260 30534 20312 30540
rect 18972 30320 19024 30326
rect 20272 30274 20300 30534
rect 18972 30262 19024 30268
rect 18984 29850 19012 30262
rect 19340 30252 19392 30258
rect 19340 30194 19392 30200
rect 20180 30246 20300 30274
rect 18972 29844 19024 29850
rect 18972 29786 19024 29792
rect 19352 29782 19380 30194
rect 19708 30048 19760 30054
rect 19708 29990 19760 29996
rect 19892 30048 19944 30054
rect 19892 29990 19944 29996
rect 19720 29782 19748 29990
rect 19340 29776 19392 29782
rect 19340 29718 19392 29724
rect 19708 29776 19760 29782
rect 19708 29718 19760 29724
rect 19156 29504 19208 29510
rect 19156 29446 19208 29452
rect 19168 29102 19196 29446
rect 19156 29096 19208 29102
rect 19156 29038 19208 29044
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19812 28218 19840 28494
rect 19800 28212 19852 28218
rect 19800 28154 19852 28160
rect 19708 28008 19760 28014
rect 19708 27950 19760 27956
rect 19720 27538 19748 27950
rect 18972 27532 19024 27538
rect 18972 27474 19024 27480
rect 19708 27532 19760 27538
rect 19708 27474 19760 27480
rect 18984 26466 19012 27474
rect 19248 27464 19300 27470
rect 19248 27406 19300 27412
rect 19800 27464 19852 27470
rect 19800 27406 19852 27412
rect 19064 27328 19116 27334
rect 19064 27270 19116 27276
rect 19156 27328 19208 27334
rect 19156 27270 19208 27276
rect 19076 26858 19104 27270
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 19168 26518 19196 27270
rect 19260 26586 19288 27406
rect 19524 26852 19576 26858
rect 19524 26794 19576 26800
rect 19536 26586 19564 26794
rect 19812 26586 19840 27406
rect 19248 26580 19300 26586
rect 19248 26522 19300 26528
rect 19524 26580 19576 26586
rect 19524 26522 19576 26528
rect 19800 26580 19852 26586
rect 19800 26522 19852 26528
rect 18892 26450 19012 26466
rect 19156 26512 19208 26518
rect 19156 26454 19208 26460
rect 18880 26444 19012 26450
rect 18932 26438 19012 26444
rect 18880 26386 18932 26392
rect 18984 26234 19012 26438
rect 19432 26376 19484 26382
rect 19154 26344 19210 26353
rect 19210 26302 19288 26330
rect 19432 26318 19484 26324
rect 19154 26279 19210 26288
rect 18984 26206 19196 26234
rect 19064 25152 19116 25158
rect 19064 25094 19116 25100
rect 19076 24886 19104 25094
rect 18972 24880 19024 24886
rect 18972 24822 19024 24828
rect 19064 24880 19116 24886
rect 19064 24822 19116 24828
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18892 24070 18920 24210
rect 18984 24154 19012 24822
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19076 24342 19104 24686
rect 19064 24336 19116 24342
rect 19064 24278 19116 24284
rect 19168 24274 19196 26206
rect 19156 24268 19208 24274
rect 19156 24210 19208 24216
rect 18984 24126 19196 24154
rect 18880 24064 18932 24070
rect 18880 24006 18932 24012
rect 18892 23526 18920 24006
rect 18880 23520 18932 23526
rect 18880 23462 18932 23468
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 18708 23174 18828 23202
rect 18708 22794 18736 23174
rect 18892 22982 18920 23462
rect 18972 23112 19024 23118
rect 18972 23054 19024 23060
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18708 22766 18920 22794
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18800 21894 18828 21966
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18800 21554 18828 21830
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18708 20602 18736 20742
rect 18696 20596 18748 20602
rect 18696 20538 18748 20544
rect 18708 20466 18736 20538
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18602 19952 18658 19961
rect 18420 19916 18472 19922
rect 18602 19887 18658 19896
rect 18420 19858 18472 19864
rect 18144 19848 18196 19854
rect 18892 19825 18920 22766
rect 18984 22030 19012 23054
rect 19076 22574 19104 23462
rect 19168 22710 19196 24126
rect 19156 22704 19208 22710
rect 19156 22646 19208 22652
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18972 21888 19024 21894
rect 19168 21842 19196 22646
rect 19024 21836 19196 21842
rect 18972 21830 19196 21836
rect 18984 21814 19196 21830
rect 18144 19790 18196 19796
rect 18878 19816 18934 19825
rect 18878 19751 18934 19760
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18432 19310 18460 19654
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 18052 19168 18104 19174
rect 18052 19110 18104 19116
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17960 17536 18012 17542
rect 17960 17478 18012 17484
rect 17972 17270 18000 17478
rect 17960 17264 18012 17270
rect 17774 17232 17830 17241
rect 17960 17206 18012 17212
rect 18064 17202 18092 17750
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 18156 17270 18184 17546
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 17774 17167 17830 17176
rect 18052 17196 18104 17202
rect 17788 17082 17816 17167
rect 18052 17138 18104 17144
rect 17788 17066 18092 17082
rect 17788 17060 18104 17066
rect 17788 17054 18052 17060
rect 18052 17002 18104 17008
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17960 16992 18012 16998
rect 17960 16934 18012 16940
rect 17776 16720 17828 16726
rect 17776 16662 17828 16668
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17788 15978 17816 16662
rect 17880 16590 17908 16934
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17776 15972 17828 15978
rect 17776 15914 17828 15920
rect 17500 15700 17552 15706
rect 17328 15660 17500 15688
rect 17224 15564 17276 15570
rect 17224 15506 17276 15512
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 17040 15156 17092 15162
rect 17040 15098 17092 15104
rect 16580 14884 16632 14890
rect 16580 14826 16632 14832
rect 16684 14878 16804 14906
rect 16684 14482 16712 14878
rect 16672 14476 16724 14482
rect 16672 14418 16724 14424
rect 16684 14385 16712 14418
rect 16670 14376 16726 14385
rect 16670 14311 16726 14320
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16592 13938 16620 14214
rect 16580 13932 16632 13938
rect 16580 13874 16632 13880
rect 16408 13790 16620 13818
rect 16592 13530 16620 13790
rect 16684 13734 16712 14311
rect 16672 13728 16724 13734
rect 16672 13670 16724 13676
rect 16868 13530 16896 15098
rect 17052 14618 17080 15098
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16592 13258 16620 13466
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16868 12986 16896 13330
rect 16856 12980 16908 12986
rect 16856 12922 16908 12928
rect 16868 12832 16896 12922
rect 16960 12850 16988 14418
rect 17130 13696 17186 13705
rect 17130 13631 17186 13640
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 16776 12804 16896 12832
rect 16948 12844 17000 12850
rect 16672 12776 16724 12782
rect 16672 12718 16724 12724
rect 15948 12406 16252 12434
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15108 11212 15160 11218
rect 15108 11154 15160 11160
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 13924 9608 14044 9636
rect 13544 9376 13596 9382
rect 13544 9318 13596 9324
rect 13556 8974 13584 9318
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13924 8922 13952 9608
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 14016 9042 14044 9454
rect 14096 9376 14148 9382
rect 14096 9318 14148 9324
rect 14108 9178 14136 9318
rect 14306 9276 14614 9285
rect 14306 9274 14312 9276
rect 14368 9274 14392 9276
rect 14448 9274 14472 9276
rect 14528 9274 14552 9276
rect 14608 9274 14614 9276
rect 14368 9222 14370 9274
rect 14550 9222 14552 9274
rect 14306 9220 14312 9222
rect 14368 9220 14392 9222
rect 14448 9220 14472 9222
rect 14528 9220 14552 9222
rect 14608 9220 14614 9222
rect 14306 9211 14614 9220
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14096 8968 14148 8974
rect 13556 8430 13584 8910
rect 13924 8894 14044 8922
rect 14096 8910 14148 8916
rect 14016 8838 14044 8894
rect 14004 8832 14056 8838
rect 14004 8774 14056 8780
rect 13646 8732 13954 8741
rect 13646 8730 13652 8732
rect 13708 8730 13732 8732
rect 13788 8730 13812 8732
rect 13868 8730 13892 8732
rect 13948 8730 13954 8732
rect 13708 8678 13710 8730
rect 13890 8678 13892 8730
rect 13646 8676 13652 8678
rect 13708 8676 13732 8678
rect 13788 8676 13812 8678
rect 13868 8676 13892 8678
rect 13948 8676 13954 8678
rect 13646 8667 13954 8676
rect 14016 8566 14044 8774
rect 14004 8560 14056 8566
rect 14004 8502 14056 8508
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13820 8424 13872 8430
rect 13820 8366 13872 8372
rect 13556 8294 13584 8366
rect 13544 8288 13596 8294
rect 13266 8256 13322 8265
rect 13544 8230 13596 8236
rect 13266 8191 13322 8200
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 13188 7206 13216 7822
rect 13280 7546 13308 8191
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 12532 6928 12584 6934
rect 12532 6870 12584 6876
rect 12990 6896 13046 6905
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 12544 5234 12572 6870
rect 12990 6831 13046 6840
rect 13268 6860 13320 6866
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12900 6112 12952 6118
rect 12900 6054 12952 6060
rect 12820 5778 12848 6054
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 12912 5234 12940 6054
rect 13004 5914 13032 6831
rect 13268 6802 13320 6808
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13188 6458 13216 6598
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13280 6390 13308 6802
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 12992 5908 13044 5914
rect 12992 5850 13044 5856
rect 13004 5710 13032 5850
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12990 5536 13046 5545
rect 12990 5471 13046 5480
rect 13004 5370 13032 5471
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 12256 5228 12308 5234
rect 12256 5170 12308 5176
rect 12532 5228 12584 5234
rect 12900 5228 12952 5234
rect 12584 5188 12664 5216
rect 12532 5170 12584 5176
rect 12268 4826 12296 5170
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12636 4146 12664 5188
rect 12900 5170 12952 5176
rect 13004 4826 13032 5306
rect 12992 4820 13044 4826
rect 12992 4762 13044 4768
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 12636 3602 12664 4082
rect 13372 3738 13400 7822
rect 13728 7744 13780 7750
rect 13832 7732 13860 8366
rect 13912 7880 13964 7886
rect 13964 7840 14044 7868
rect 13912 7822 13964 7828
rect 13780 7704 13860 7732
rect 13728 7686 13780 7692
rect 13646 7644 13954 7653
rect 13646 7642 13652 7644
rect 13708 7642 13732 7644
rect 13788 7642 13812 7644
rect 13868 7642 13892 7644
rect 13948 7642 13954 7644
rect 13708 7590 13710 7642
rect 13890 7590 13892 7642
rect 13646 7588 13652 7590
rect 13708 7588 13732 7590
rect 13788 7588 13812 7590
rect 13868 7588 13892 7590
rect 13948 7588 13954 7590
rect 13646 7579 13954 7588
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13556 6866 13584 6938
rect 13648 6866 13676 7482
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13464 6100 13492 6802
rect 13646 6556 13954 6565
rect 13646 6554 13652 6556
rect 13708 6554 13732 6556
rect 13788 6554 13812 6556
rect 13868 6554 13892 6556
rect 13948 6554 13954 6556
rect 13708 6502 13710 6554
rect 13890 6502 13892 6554
rect 13646 6500 13652 6502
rect 13708 6500 13732 6502
rect 13788 6500 13812 6502
rect 13868 6500 13892 6502
rect 13948 6500 13954 6502
rect 13646 6491 13954 6500
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13544 6112 13596 6118
rect 13464 6072 13544 6100
rect 13544 6054 13596 6060
rect 13556 5352 13584 6054
rect 13924 5710 13952 6122
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13646 5468 13954 5477
rect 13646 5466 13652 5468
rect 13708 5466 13732 5468
rect 13788 5466 13812 5468
rect 13868 5466 13892 5468
rect 13948 5466 13954 5468
rect 13708 5414 13710 5466
rect 13890 5414 13892 5466
rect 13646 5412 13652 5414
rect 13708 5412 13732 5414
rect 13788 5412 13812 5414
rect 13868 5412 13892 5414
rect 13948 5412 13954 5414
rect 13646 5403 13954 5412
rect 13556 5324 13676 5352
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13464 4282 13492 4966
rect 13556 4826 13584 5034
rect 13648 4826 13676 5324
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 14016 4622 14044 7840
rect 14108 7274 14136 8910
rect 14384 8634 14412 9046
rect 14660 8974 14688 9998
rect 14936 9722 14964 9998
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 14648 8968 14700 8974
rect 14648 8910 14700 8916
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14306 8188 14614 8197
rect 14306 8186 14312 8188
rect 14368 8186 14392 8188
rect 14448 8186 14472 8188
rect 14528 8186 14552 8188
rect 14608 8186 14614 8188
rect 14368 8134 14370 8186
rect 14550 8134 14552 8186
rect 14306 8132 14312 8134
rect 14368 8132 14392 8134
rect 14448 8132 14472 8134
rect 14528 8132 14552 8134
rect 14608 8132 14614 8134
rect 14306 8123 14614 8132
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14200 7954 14228 8026
rect 14188 7948 14240 7954
rect 14188 7890 14240 7896
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14096 7268 14148 7274
rect 14096 7210 14148 7216
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 13452 4276 13504 4282
rect 13556 4264 13584 4558
rect 14004 4480 14056 4486
rect 14004 4422 14056 4428
rect 13646 4380 13954 4389
rect 13646 4378 13652 4380
rect 13708 4378 13732 4380
rect 13788 4378 13812 4380
rect 13868 4378 13892 4380
rect 13948 4378 13954 4380
rect 13708 4326 13710 4378
rect 13890 4326 13892 4378
rect 13646 4324 13652 4326
rect 13708 4324 13732 4326
rect 13788 4324 13812 4326
rect 13868 4324 13892 4326
rect 13948 4324 13954 4326
rect 13646 4315 13954 4324
rect 13556 4236 13676 4264
rect 13452 4218 13504 4224
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13556 3738 13584 3946
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13648 3602 13676 4236
rect 14016 3738 14044 4422
rect 14108 4146 14136 7210
rect 14200 6914 14228 7686
rect 14306 7100 14614 7109
rect 14306 7098 14312 7100
rect 14368 7098 14392 7100
rect 14448 7098 14472 7100
rect 14528 7098 14552 7100
rect 14608 7098 14614 7100
rect 14368 7046 14370 7098
rect 14550 7046 14552 7098
rect 14306 7044 14312 7046
rect 14368 7044 14392 7046
rect 14448 7044 14472 7046
rect 14528 7044 14552 7046
rect 14608 7044 14614 7046
rect 14306 7035 14614 7044
rect 14200 6886 14320 6914
rect 14188 6248 14240 6254
rect 14188 6190 14240 6196
rect 14200 5370 14228 6190
rect 14292 6186 14320 6886
rect 14660 6866 14688 8774
rect 14936 8634 14964 8910
rect 15028 8838 15056 9522
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14752 7750 14780 8570
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14844 7750 14872 8230
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14844 6662 14872 7686
rect 14936 6866 14964 8366
rect 15120 7478 15148 11154
rect 15200 10600 15252 10606
rect 15200 10542 15252 10548
rect 15212 9722 15240 10542
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15200 9716 15252 9722
rect 15200 9658 15252 9664
rect 15304 9586 15332 10406
rect 15396 10062 15424 10406
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15396 9722 15424 9998
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15488 9602 15516 11494
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15580 10538 15608 11086
rect 15660 10736 15712 10742
rect 15660 10678 15712 10684
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10266 15608 10474
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15396 9574 15516 9602
rect 15396 8838 15424 9574
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15028 6730 15056 6802
rect 15016 6724 15068 6730
rect 15016 6666 15068 6672
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14306 6012 14614 6021
rect 14306 6010 14312 6012
rect 14368 6010 14392 6012
rect 14448 6010 14472 6012
rect 14528 6010 14552 6012
rect 14608 6010 14614 6012
rect 14368 5958 14370 6010
rect 14550 5958 14552 6010
rect 14306 5956 14312 5958
rect 14368 5956 14392 5958
rect 14448 5956 14472 5958
rect 14528 5956 14552 5958
rect 14608 5956 14614 5958
rect 14306 5947 14614 5956
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14306 4924 14614 4933
rect 14306 4922 14312 4924
rect 14368 4922 14392 4924
rect 14448 4922 14472 4924
rect 14528 4922 14552 4924
rect 14608 4922 14614 4924
rect 14368 4870 14370 4922
rect 14550 4870 14552 4922
rect 14306 4868 14312 4870
rect 14368 4868 14392 4870
rect 14448 4868 14472 4870
rect 14528 4868 14552 4870
rect 14608 4868 14614 4870
rect 14306 4859 14614 4868
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14096 4140 14148 4146
rect 14096 4082 14148 4088
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13646 3292 13954 3301
rect 13646 3290 13652 3292
rect 13708 3290 13732 3292
rect 13788 3290 13812 3292
rect 13868 3290 13892 3292
rect 13948 3290 13954 3292
rect 13708 3238 13710 3290
rect 13890 3238 13892 3290
rect 13646 3236 13652 3238
rect 13708 3236 13732 3238
rect 13788 3236 13812 3238
rect 13868 3236 13892 3238
rect 13948 3236 13954 3238
rect 13646 3227 13954 3236
rect 14200 3194 14228 4558
rect 14660 4282 14688 6054
rect 14844 5914 14872 6598
rect 15028 6458 15056 6666
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14844 5778 14872 5850
rect 14832 5772 14884 5778
rect 14884 5732 14964 5760
rect 14832 5714 14884 5720
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14306 3836 14614 3845
rect 14306 3834 14312 3836
rect 14368 3834 14392 3836
rect 14448 3834 14472 3836
rect 14528 3834 14552 3836
rect 14608 3834 14614 3836
rect 14368 3782 14370 3834
rect 14550 3782 14552 3834
rect 14306 3780 14312 3782
rect 14368 3780 14392 3782
rect 14448 3780 14472 3782
rect 14528 3780 14552 3782
rect 14608 3780 14614 3782
rect 14306 3771 14614 3780
rect 14844 3194 14872 5510
rect 14936 5166 14964 5732
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15028 3194 15056 5646
rect 15120 4622 15148 7414
rect 15212 7342 15240 7822
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7546 15332 7686
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15396 7426 15424 8774
rect 15568 7812 15620 7818
rect 15568 7754 15620 7760
rect 15304 7398 15424 7426
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15200 6928 15252 6934
rect 15200 6870 15252 6876
rect 15212 5710 15240 6870
rect 15304 6662 15332 7398
rect 15580 7002 15608 7754
rect 15672 7274 15700 10678
rect 15948 10470 15976 12406
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15844 9648 15896 9654
rect 15844 9590 15896 9596
rect 15856 9178 15884 9590
rect 15948 9382 15976 10406
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15856 8634 15884 9114
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15948 8412 15976 9318
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8430 16160 8774
rect 16028 8424 16080 8430
rect 15948 8384 16028 8412
rect 15752 8288 15804 8294
rect 15752 8230 15804 8236
rect 15764 7954 15792 8230
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15660 7268 15712 7274
rect 15660 7210 15712 7216
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15304 6361 15332 6598
rect 15290 6352 15346 6361
rect 15290 6287 15346 6296
rect 15292 6248 15344 6254
rect 15292 6190 15344 6196
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15212 4622 15240 5170
rect 15304 4826 15332 6190
rect 15396 5914 15424 6870
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15488 5642 15516 6938
rect 15948 6730 15976 8384
rect 16028 8366 16080 8372
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15936 6724 15988 6730
rect 15936 6666 15988 6672
rect 15948 6458 15976 6666
rect 16224 6662 16252 11494
rect 16316 10674 16344 12174
rect 16684 12102 16712 12718
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16776 11558 16804 12804
rect 16948 12786 17000 12792
rect 17052 12782 17080 12922
rect 17144 12918 17172 13631
rect 17236 13326 17264 14758
rect 17328 14482 17356 15660
rect 17500 15642 17552 15648
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17500 15360 17552 15366
rect 17500 15302 17552 15308
rect 17512 14958 17540 15302
rect 17604 15026 17632 15370
rect 17972 15162 18000 16934
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 18156 15026 18184 15982
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17684 14884 17736 14890
rect 17684 14826 17736 14832
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16856 12640 16908 12646
rect 16856 12582 16908 12588
rect 16868 12306 16896 12582
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16948 12232 17000 12238
rect 16948 12174 17000 12180
rect 16856 12096 16908 12102
rect 16856 12038 16908 12044
rect 16764 11552 16816 11558
rect 16764 11494 16816 11500
rect 16776 11218 16804 11494
rect 16764 11212 16816 11218
rect 16764 11154 16816 11160
rect 16868 11082 16896 12038
rect 16960 11830 16988 12174
rect 17236 11830 17264 13262
rect 17328 12986 17356 14418
rect 17420 14278 17448 14758
rect 17696 14618 17724 14826
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 17684 14612 17736 14618
rect 17684 14554 17736 14560
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 13394 17448 14214
rect 17512 14074 17540 14350
rect 17500 14068 17552 14074
rect 17500 14010 17552 14016
rect 17972 13802 18000 14758
rect 18064 13938 18092 14758
rect 18156 14074 18184 14962
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17408 13388 17460 13394
rect 17408 13330 17460 13336
rect 17696 12986 17724 13670
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17684 12980 17736 12986
rect 17684 12922 17736 12928
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11830 17448 12038
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 16856 11076 16908 11082
rect 16856 11018 16908 11024
rect 16672 11008 16724 11014
rect 16672 10950 16724 10956
rect 16684 10674 16712 10950
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16672 10668 16724 10674
rect 16672 10610 16724 10616
rect 16764 10124 16816 10130
rect 16764 10066 16816 10072
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16592 9586 16620 9998
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16684 9178 16712 9454
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 16672 9036 16724 9042
rect 16672 8978 16724 8984
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 7002 16344 8910
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16500 8634 16528 8774
rect 16488 8628 16540 8634
rect 16488 8570 16540 8576
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 8022 16620 8298
rect 16580 8016 16632 8022
rect 16580 7958 16632 7964
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16304 6996 16356 7002
rect 16304 6938 16356 6944
rect 16408 6866 16436 7822
rect 16684 7546 16712 8978
rect 16776 8022 16804 10066
rect 16764 8016 16816 8022
rect 16764 7958 16816 7964
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16776 7342 16804 7958
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16764 7200 16816 7206
rect 16764 7142 16816 7148
rect 16776 6934 16804 7142
rect 16764 6928 16816 6934
rect 16764 6870 16816 6876
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 15936 6452 15988 6458
rect 15936 6394 15988 6400
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5914 15792 6054
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15476 5636 15528 5642
rect 15476 5578 15528 5584
rect 15750 5264 15806 5273
rect 15948 5234 15976 6394
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16028 5568 16080 5574
rect 16028 5510 16080 5516
rect 15750 5199 15752 5208
rect 15804 5199 15806 5208
rect 15936 5228 15988 5234
rect 15752 5170 15804 5176
rect 15936 5170 15988 5176
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15568 4684 15620 4690
rect 15568 4626 15620 4632
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 11520 2984 11572 2990
rect 11520 2926 11572 2932
rect 12268 800 12296 2994
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13648 1578 13676 2926
rect 14306 2748 14614 2757
rect 14306 2746 14312 2748
rect 14368 2746 14392 2748
rect 14448 2746 14472 2748
rect 14528 2746 14552 2748
rect 14608 2746 14614 2748
rect 14368 2694 14370 2746
rect 14550 2694 14552 2746
rect 14306 2692 14312 2694
rect 14368 2692 14392 2694
rect 14448 2692 14472 2694
rect 14528 2692 14552 2694
rect 14608 2692 14614 2694
rect 14306 2683 14614 2692
rect 13556 1550 13676 1578
rect 13556 800 13584 1550
rect 14844 800 14872 2994
rect 15396 2990 15424 3878
rect 15488 3602 15516 4014
rect 15580 3942 15608 4626
rect 15568 3936 15620 3942
rect 15568 3878 15620 3884
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15580 3126 15608 3878
rect 15856 3670 15884 3878
rect 16040 3738 16068 5510
rect 16408 5370 16436 6190
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16120 4616 16172 4622
rect 16120 4558 16172 4564
rect 16028 3732 16080 3738
rect 16028 3674 16080 3680
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 16132 3602 16160 4558
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16224 4282 16252 4422
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 16120 3596 16172 3602
rect 16120 3538 16172 3544
rect 15568 3120 15620 3126
rect 15568 3062 15620 3068
rect 16316 2990 16344 5102
rect 16396 4684 16448 4690
rect 16396 4626 16448 4632
rect 16408 3058 16436 4626
rect 16592 3738 16620 6054
rect 16684 5166 16712 6734
rect 16868 6390 16896 11018
rect 17328 10266 17356 11086
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16960 8634 16988 8774
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16868 5166 16896 6122
rect 17052 5166 17080 7278
rect 17328 6458 17356 7278
rect 17316 6452 17368 6458
rect 17316 6394 17368 6400
rect 17316 6248 17368 6254
rect 17316 6190 17368 6196
rect 17328 5914 17356 6190
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17144 5370 17172 5782
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 17040 5160 17092 5166
rect 17040 5102 17092 5108
rect 16948 3936 17000 3942
rect 17052 3924 17080 5102
rect 17512 4826 17540 12854
rect 17972 12782 18000 13466
rect 18156 12986 18184 14010
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 18248 12714 18276 17478
rect 18340 17105 18368 18362
rect 18524 17134 18552 18634
rect 18892 17785 18920 19751
rect 18984 17921 19012 21814
rect 19064 21072 19116 21078
rect 19064 21014 19116 21020
rect 19076 20602 19104 21014
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 19076 20058 19104 20334
rect 19260 20058 19288 26302
rect 19444 25702 19472 26318
rect 19536 26234 19564 26522
rect 19904 26466 19932 29990
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19996 27130 20024 27270
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 20076 26784 20128 26790
rect 20076 26726 20128 26732
rect 20180 26738 20208 30246
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20272 29306 20300 30126
rect 20364 29850 20392 30670
rect 20732 30394 20760 30670
rect 21006 30492 21314 30501
rect 21006 30490 21012 30492
rect 21068 30490 21092 30492
rect 21148 30490 21172 30492
rect 21228 30490 21252 30492
rect 21308 30490 21314 30492
rect 21068 30438 21070 30490
rect 21250 30438 21252 30490
rect 21006 30436 21012 30438
rect 21068 30436 21092 30438
rect 21148 30436 21172 30438
rect 21228 30436 21252 30438
rect 21308 30436 21314 30438
rect 21006 30427 21314 30436
rect 20720 30388 20772 30394
rect 20720 30330 20772 30336
rect 20444 30048 20496 30054
rect 20444 29990 20496 29996
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20260 29300 20312 29306
rect 20260 29242 20312 29248
rect 20364 28694 20392 29786
rect 20456 29782 20484 29990
rect 21468 29850 21496 32302
rect 21928 32286 22048 32314
rect 21666 32124 21974 32133
rect 21666 32122 21672 32124
rect 21728 32122 21752 32124
rect 21808 32122 21832 32124
rect 21888 32122 21912 32124
rect 21968 32122 21974 32124
rect 21728 32070 21730 32122
rect 21910 32070 21912 32122
rect 21666 32068 21672 32070
rect 21728 32068 21752 32070
rect 21808 32068 21832 32070
rect 21888 32068 21912 32070
rect 21968 32068 21974 32070
rect 21666 32059 21974 32068
rect 22020 32026 22048 32286
rect 22008 32020 22060 32026
rect 22008 31962 22060 31968
rect 23860 31958 23888 33544
rect 25148 31958 25176 33544
rect 25964 32292 26016 32298
rect 25964 32234 26016 32240
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 25792 32026 25820 32166
rect 25780 32020 25832 32026
rect 25780 31962 25832 31968
rect 23848 31952 23900 31958
rect 23848 31894 23900 31900
rect 25136 31952 25188 31958
rect 25136 31894 25188 31900
rect 24032 31884 24084 31890
rect 24032 31826 24084 31832
rect 25504 31884 25556 31890
rect 25504 31826 25556 31832
rect 24044 31754 24072 31826
rect 24044 31726 24164 31754
rect 22376 31680 22428 31686
rect 22376 31622 22428 31628
rect 22100 31272 22152 31278
rect 22100 31214 22152 31220
rect 21666 31036 21974 31045
rect 21666 31034 21672 31036
rect 21728 31034 21752 31036
rect 21808 31034 21832 31036
rect 21888 31034 21912 31036
rect 21968 31034 21974 31036
rect 21728 30982 21730 31034
rect 21910 30982 21912 31034
rect 21666 30980 21672 30982
rect 21728 30980 21752 30982
rect 21808 30980 21832 30982
rect 21888 30980 21912 30982
rect 21968 30980 21974 30982
rect 21666 30971 21974 30980
rect 22112 30394 22140 31214
rect 22388 30938 22416 31622
rect 23664 31408 23716 31414
rect 23664 31350 23716 31356
rect 23112 31272 23164 31278
rect 23112 31214 23164 31220
rect 22376 30932 22428 30938
rect 22376 30874 22428 30880
rect 22928 30728 22980 30734
rect 22928 30670 22980 30676
rect 22284 30592 22336 30598
rect 22284 30534 22336 30540
rect 22100 30388 22152 30394
rect 22100 30330 22152 30336
rect 22100 30252 22152 30258
rect 22100 30194 22152 30200
rect 21548 30184 21600 30190
rect 21548 30126 21600 30132
rect 20720 29844 20772 29850
rect 20720 29786 20772 29792
rect 21456 29844 21508 29850
rect 21456 29786 21508 29792
rect 20444 29776 20496 29782
rect 20444 29718 20496 29724
rect 20732 29034 20760 29786
rect 21560 29510 21588 30126
rect 22008 30116 22060 30122
rect 22008 30058 22060 30064
rect 21666 29948 21974 29957
rect 21666 29946 21672 29948
rect 21728 29946 21752 29948
rect 21808 29946 21832 29948
rect 21888 29946 21912 29948
rect 21968 29946 21974 29948
rect 21728 29894 21730 29946
rect 21910 29894 21912 29946
rect 21666 29892 21672 29894
rect 21728 29892 21752 29894
rect 21808 29892 21832 29894
rect 21888 29892 21912 29894
rect 21968 29892 21974 29894
rect 21666 29883 21974 29892
rect 22020 29850 22048 30058
rect 22008 29844 22060 29850
rect 22008 29786 22060 29792
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21006 29404 21314 29413
rect 21006 29402 21012 29404
rect 21068 29402 21092 29404
rect 21148 29402 21172 29404
rect 21228 29402 21252 29404
rect 21308 29402 21314 29404
rect 21068 29350 21070 29402
rect 21250 29350 21252 29402
rect 21006 29348 21012 29350
rect 21068 29348 21092 29350
rect 21148 29348 21172 29350
rect 21228 29348 21252 29350
rect 21308 29348 21314 29350
rect 21006 29339 21314 29348
rect 21560 29238 21588 29446
rect 21548 29232 21600 29238
rect 21548 29174 21600 29180
rect 22112 29170 22140 30194
rect 22296 30054 22324 30534
rect 22560 30388 22612 30394
rect 22560 30330 22612 30336
rect 22284 30048 22336 30054
rect 22284 29990 22336 29996
rect 22572 29714 22600 30330
rect 22744 30116 22796 30122
rect 22744 30058 22796 30064
rect 22756 29850 22784 30058
rect 22940 30054 22968 30670
rect 22928 30048 22980 30054
rect 22928 29990 22980 29996
rect 22744 29844 22796 29850
rect 22744 29786 22796 29792
rect 23124 29714 23152 31214
rect 23676 31142 23704 31350
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 24032 31272 24084 31278
rect 24032 31214 24084 31220
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23480 30252 23532 30258
rect 23480 30194 23532 30200
rect 22560 29708 22612 29714
rect 22560 29650 22612 29656
rect 23112 29708 23164 29714
rect 23112 29650 23164 29656
rect 22100 29164 22152 29170
rect 22100 29106 22152 29112
rect 20720 29028 20772 29034
rect 20720 28970 20772 28976
rect 20444 28960 20496 28966
rect 20444 28902 20496 28908
rect 20352 28688 20404 28694
rect 20352 28630 20404 28636
rect 20456 28422 20484 28902
rect 21666 28860 21974 28869
rect 21666 28858 21672 28860
rect 21728 28858 21752 28860
rect 21808 28858 21832 28860
rect 21888 28858 21912 28860
rect 21968 28858 21974 28860
rect 21728 28806 21730 28858
rect 21910 28806 21912 28858
rect 21666 28804 21672 28806
rect 21728 28804 21752 28806
rect 21808 28804 21832 28806
rect 21888 28804 21912 28806
rect 21968 28804 21974 28806
rect 21666 28795 21974 28804
rect 21364 28688 21416 28694
rect 21364 28630 21416 28636
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 20456 27606 20484 28358
rect 21006 28316 21314 28325
rect 21006 28314 21012 28316
rect 21068 28314 21092 28316
rect 21148 28314 21172 28316
rect 21228 28314 21252 28316
rect 21308 28314 21314 28316
rect 21068 28262 21070 28314
rect 21250 28262 21252 28314
rect 21006 28260 21012 28262
rect 21068 28260 21092 28262
rect 21148 28260 21172 28262
rect 21228 28260 21252 28262
rect 21308 28260 21314 28262
rect 21006 28251 21314 28260
rect 20444 27600 20496 27606
rect 20444 27542 20496 27548
rect 21006 27228 21314 27237
rect 21006 27226 21012 27228
rect 21068 27226 21092 27228
rect 21148 27226 21172 27228
rect 21228 27226 21252 27228
rect 21308 27226 21314 27228
rect 21068 27174 21070 27226
rect 21250 27174 21252 27226
rect 21006 27172 21012 27174
rect 21068 27172 21092 27174
rect 21148 27172 21172 27174
rect 21228 27172 21252 27174
rect 21308 27172 21314 27174
rect 21006 27163 21314 27172
rect 21376 26994 21404 28630
rect 22572 28626 22600 29650
rect 22652 29028 22704 29034
rect 22652 28970 22704 28976
rect 22664 28762 22692 28970
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 23492 28694 23520 30194
rect 23676 29646 23704 31078
rect 23768 30938 23796 31214
rect 23940 31136 23992 31142
rect 23940 31078 23992 31084
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23768 29850 23796 30874
rect 23848 30796 23900 30802
rect 23848 30738 23900 30744
rect 23860 30394 23888 30738
rect 23952 30394 23980 31078
rect 24044 30802 24072 31214
rect 24032 30796 24084 30802
rect 24032 30738 24084 30744
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 23940 30388 23992 30394
rect 23940 30330 23992 30336
rect 23756 29844 23808 29850
rect 23756 29786 23808 29792
rect 23664 29640 23716 29646
rect 23664 29582 23716 29588
rect 23768 29510 23796 29786
rect 23756 29504 23808 29510
rect 23756 29446 23808 29452
rect 23768 29322 23796 29446
rect 23768 29294 23888 29322
rect 23756 29164 23808 29170
rect 23756 29106 23808 29112
rect 23572 28960 23624 28966
rect 23572 28902 23624 28908
rect 23584 28762 23612 28902
rect 23572 28756 23624 28762
rect 23572 28698 23624 28704
rect 23480 28688 23532 28694
rect 23480 28630 23532 28636
rect 22100 28620 22152 28626
rect 22100 28562 22152 28568
rect 22560 28620 22612 28626
rect 22560 28562 22612 28568
rect 22112 28014 22140 28562
rect 22100 28008 22152 28014
rect 22100 27950 22152 27956
rect 23112 28008 23164 28014
rect 23112 27950 23164 27956
rect 21666 27772 21974 27781
rect 21666 27770 21672 27772
rect 21728 27770 21752 27772
rect 21808 27770 21832 27772
rect 21888 27770 21912 27772
rect 21968 27770 21974 27772
rect 21728 27718 21730 27770
rect 21910 27718 21912 27770
rect 21666 27716 21672 27718
rect 21728 27716 21752 27718
rect 21808 27716 21832 27718
rect 21888 27716 21912 27718
rect 21968 27716 21974 27718
rect 21666 27707 21974 27716
rect 22008 27532 22060 27538
rect 22112 27520 22140 27950
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22060 27492 22140 27520
rect 22008 27474 22060 27480
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 21364 26988 21416 26994
rect 21416 26948 21496 26976
rect 21364 26930 21416 26936
rect 20088 26586 20116 26726
rect 20180 26710 20484 26738
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19904 26438 20208 26466
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 19536 26206 19748 26234
rect 19720 26042 19748 26206
rect 19708 26036 19760 26042
rect 19708 25978 19760 25984
rect 19616 25900 19668 25906
rect 19616 25842 19668 25848
rect 19892 25900 19944 25906
rect 19892 25842 19944 25848
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 19352 23254 19380 24550
rect 19444 24206 19472 25638
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19536 24954 19564 25230
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19628 24818 19656 25842
rect 19904 25702 19932 25842
rect 19892 25696 19944 25702
rect 19892 25638 19944 25644
rect 20088 24818 20116 26250
rect 20180 26234 20208 26438
rect 20180 26206 20300 26234
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24342 20116 24754
rect 20076 24336 20128 24342
rect 20076 24278 20128 24284
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 19708 23656 19760 23662
rect 19708 23598 19760 23604
rect 19340 23248 19392 23254
rect 19340 23190 19392 23196
rect 19352 22506 19380 23190
rect 19340 22500 19392 22506
rect 19340 22442 19392 22448
rect 19720 22438 19748 23598
rect 19708 22432 19760 22438
rect 19708 22374 19760 22380
rect 19800 22432 19852 22438
rect 19800 22374 19852 22380
rect 20076 22432 20128 22438
rect 20076 22374 20128 22380
rect 19720 22030 19748 22374
rect 19812 22166 19840 22374
rect 20088 22234 20116 22374
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19800 22160 19852 22166
rect 19800 22102 19852 22108
rect 20272 22094 20300 26206
rect 20352 23520 20404 23526
rect 20352 23462 20404 23468
rect 20364 23254 20392 23462
rect 20352 23248 20404 23254
rect 20352 23190 20404 23196
rect 20180 22066 20300 22094
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 20088 21486 20116 21830
rect 20076 21480 20128 21486
rect 19996 21428 20076 21434
rect 19996 21422 20128 21428
rect 19800 21412 19852 21418
rect 19800 21354 19852 21360
rect 19996 21406 20116 21422
rect 19812 20466 19840 21354
rect 19800 20460 19852 20466
rect 19800 20402 19852 20408
rect 19064 20052 19116 20058
rect 19064 19994 19116 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19260 19334 19288 19994
rect 19812 19514 19840 20402
rect 19996 20330 20024 21406
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19800 19508 19852 19514
rect 19800 19450 19852 19456
rect 19168 19306 19288 19334
rect 19168 19242 19196 19306
rect 19156 19236 19208 19242
rect 19156 19178 19208 19184
rect 19168 18766 19196 19178
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19260 18902 19288 19110
rect 19248 18896 19300 18902
rect 19248 18838 19300 18844
rect 19156 18760 19208 18766
rect 19156 18702 19208 18708
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19168 18358 19196 18702
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19076 18057 19104 18294
rect 19248 18080 19300 18086
rect 19062 18048 19118 18057
rect 19248 18022 19300 18028
rect 19062 17983 19118 17992
rect 18970 17912 19026 17921
rect 18970 17847 19026 17856
rect 19076 17814 19104 17983
rect 19064 17808 19116 17814
rect 18878 17776 18934 17785
rect 19064 17750 19116 17756
rect 18878 17711 18934 17720
rect 19260 17134 19288 18022
rect 19352 17202 19380 18702
rect 19614 18456 19670 18465
rect 19614 18391 19670 18400
rect 19432 18352 19484 18358
rect 19522 18320 19578 18329
rect 19484 18300 19522 18306
rect 19432 18294 19522 18300
rect 19444 18278 19522 18294
rect 19628 18290 19656 18391
rect 19522 18255 19578 18264
rect 19616 18284 19668 18290
rect 19668 18244 19748 18272
rect 19616 18226 19668 18232
rect 19524 18216 19576 18222
rect 19524 18158 19576 18164
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19444 17746 19472 18090
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19340 17196 19392 17202
rect 19340 17138 19392 17144
rect 18512 17128 18564 17134
rect 18326 17096 18382 17105
rect 18512 17070 18564 17076
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 18326 17031 18382 17040
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 16114 18460 16390
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18328 14884 18380 14890
rect 18328 14826 18380 14832
rect 18340 14482 18368 14826
rect 18328 14476 18380 14482
rect 18328 14418 18380 14424
rect 18524 13530 18552 17070
rect 19444 16658 19472 17682
rect 19536 16658 19564 18158
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19432 16652 19484 16658
rect 19432 16594 19484 16600
rect 19524 16652 19576 16658
rect 19524 16594 19576 16600
rect 19156 15972 19208 15978
rect 19156 15914 19208 15920
rect 19168 15706 19196 15914
rect 19156 15700 19208 15706
rect 19156 15642 19208 15648
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18708 14618 18736 14894
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 19168 14482 19196 15370
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18616 14074 18644 14214
rect 18604 14068 18656 14074
rect 18604 14010 18656 14016
rect 18708 13802 18736 14214
rect 18696 13796 18748 13802
rect 18696 13738 18748 13744
rect 18892 13530 18920 14282
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18880 13524 18932 13530
rect 18880 13466 18932 13472
rect 18972 13388 19024 13394
rect 18972 13330 19024 13336
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18604 13184 18656 13190
rect 18524 13144 18604 13172
rect 18524 12730 18552 13144
rect 18604 13126 18656 13132
rect 18604 12844 18656 12850
rect 18708 12832 18736 13262
rect 18656 12804 18736 12832
rect 18604 12786 18656 12792
rect 18052 12708 18104 12714
rect 18052 12650 18104 12656
rect 18236 12708 18288 12714
rect 18236 12650 18288 12656
rect 18420 12708 18472 12714
rect 18524 12702 18644 12730
rect 18420 12650 18472 12656
rect 18064 12434 18092 12650
rect 18432 12442 18460 12650
rect 18420 12436 18472 12442
rect 18064 12406 18184 12434
rect 18156 12102 18184 12406
rect 18420 12378 18472 12384
rect 18616 12306 18644 12702
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18708 11694 18736 12804
rect 18984 12442 19012 13330
rect 18972 12436 19024 12442
rect 19260 12434 19288 15098
rect 19536 14890 19564 15302
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 19444 14074 19472 14350
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13530 19564 13670
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19524 13184 19576 13190
rect 19628 13172 19656 17614
rect 19576 13144 19656 13172
rect 19524 13126 19576 13132
rect 18972 12378 19024 12384
rect 19168 12406 19288 12434
rect 18984 11762 19012 12378
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19076 11762 19104 12038
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18696 11688 18748 11694
rect 18696 11630 18748 11636
rect 17960 11620 18012 11626
rect 17960 11562 18012 11568
rect 18420 11620 18472 11626
rect 18420 11562 18472 11568
rect 17972 11354 18000 11562
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 18432 11082 18460 11562
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18800 11014 18828 11494
rect 18984 11354 19012 11698
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18880 11280 18932 11286
rect 18880 11222 18932 11228
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18420 10532 18472 10538
rect 18420 10474 18472 10480
rect 18432 10266 18460 10474
rect 18800 10266 18828 10950
rect 18892 10810 18920 11222
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18420 10260 18472 10266
rect 18420 10202 18472 10208
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18800 10130 18828 10202
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 18512 9920 18564 9926
rect 18512 9862 18564 9868
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17696 8974 17724 9318
rect 17972 9110 18000 9862
rect 18052 9512 18104 9518
rect 18052 9454 18104 9460
rect 17960 9104 18012 9110
rect 17960 9046 18012 9052
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17696 6662 17724 8910
rect 17960 8900 18012 8906
rect 17960 8842 18012 8848
rect 17972 7546 18000 8842
rect 18064 8090 18092 9454
rect 18524 9042 18552 9862
rect 19168 9654 19196 12406
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19260 11150 19288 12242
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11830 19472 12174
rect 19720 11898 19748 18244
rect 19996 18222 20024 20266
rect 20180 19786 20208 22066
rect 20456 20448 20484 26710
rect 20548 25838 20576 26930
rect 21468 26450 21496 26948
rect 21666 26684 21974 26693
rect 21666 26682 21672 26684
rect 21728 26682 21752 26684
rect 21808 26682 21832 26684
rect 21888 26682 21912 26684
rect 21968 26682 21974 26684
rect 21728 26630 21730 26682
rect 21910 26630 21912 26682
rect 21666 26628 21672 26630
rect 21728 26628 21752 26630
rect 21808 26628 21832 26630
rect 21888 26628 21912 26630
rect 21968 26628 21974 26630
rect 21666 26619 21974 26628
rect 21456 26444 21508 26450
rect 21456 26386 21508 26392
rect 20628 26240 20680 26246
rect 20628 26182 20680 26188
rect 20536 25832 20588 25838
rect 20536 25774 20588 25780
rect 20548 25498 20576 25774
rect 20640 25770 20668 26182
rect 21006 26140 21314 26149
rect 21006 26138 21012 26140
rect 21068 26138 21092 26140
rect 21148 26138 21172 26140
rect 21228 26138 21252 26140
rect 21308 26138 21314 26140
rect 21068 26086 21070 26138
rect 21250 26086 21252 26138
rect 21006 26084 21012 26086
rect 21068 26084 21092 26086
rect 21148 26084 21172 26086
rect 21228 26084 21252 26086
rect 21308 26084 21314 26086
rect 21006 26075 21314 26084
rect 21468 26042 21496 26386
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21456 25832 21508 25838
rect 21456 25774 21508 25780
rect 20628 25764 20680 25770
rect 20628 25706 20680 25712
rect 20536 25492 20588 25498
rect 20536 25434 20588 25440
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 24750 20668 25094
rect 21006 25052 21314 25061
rect 21006 25050 21012 25052
rect 21068 25050 21092 25052
rect 21148 25050 21172 25052
rect 21228 25050 21252 25052
rect 21308 25050 21314 25052
rect 21068 24998 21070 25050
rect 21250 24998 21252 25050
rect 21006 24996 21012 24998
rect 21068 24996 21092 24998
rect 21148 24996 21172 24998
rect 21228 24996 21252 24998
rect 21308 24996 21314 24998
rect 21006 24987 21314 24996
rect 21468 24750 21496 25774
rect 22020 25770 22048 27474
rect 22756 27470 22784 27814
rect 23124 27470 23152 27950
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 22100 27328 22152 27334
rect 22100 27270 22152 27276
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 23112 27328 23164 27334
rect 23112 27270 23164 27276
rect 22112 26858 22140 27270
rect 22100 26852 22152 26858
rect 22100 26794 22152 26800
rect 22204 26586 22232 27270
rect 23124 27130 23152 27270
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23400 26586 23428 27474
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 22468 26512 22520 26518
rect 22468 26454 22520 26460
rect 22008 25764 22060 25770
rect 22008 25706 22060 25712
rect 22284 25764 22336 25770
rect 22284 25706 22336 25712
rect 22376 25764 22428 25770
rect 22376 25706 22428 25712
rect 21666 25596 21974 25605
rect 21666 25594 21672 25596
rect 21728 25594 21752 25596
rect 21808 25594 21832 25596
rect 21888 25594 21912 25596
rect 21968 25594 21974 25596
rect 21728 25542 21730 25594
rect 21910 25542 21912 25594
rect 21666 25540 21672 25542
rect 21728 25540 21752 25542
rect 21808 25540 21832 25542
rect 21888 25540 21912 25542
rect 21968 25540 21974 25542
rect 21666 25531 21974 25540
rect 22020 25362 22048 25706
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 20628 24744 20680 24750
rect 20628 24686 20680 24692
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21666 24508 21974 24517
rect 21666 24506 21672 24508
rect 21728 24506 21752 24508
rect 21808 24506 21832 24508
rect 21888 24506 21912 24508
rect 21968 24506 21974 24508
rect 21728 24454 21730 24506
rect 21910 24454 21912 24506
rect 21666 24452 21672 24454
rect 21728 24452 21752 24454
rect 21808 24452 21832 24454
rect 21888 24452 21912 24454
rect 21968 24452 21974 24454
rect 21666 24443 21974 24452
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21456 24064 21508 24070
rect 21456 24006 21508 24012
rect 21006 23964 21314 23973
rect 21006 23962 21012 23964
rect 21068 23962 21092 23964
rect 21148 23962 21172 23964
rect 21228 23962 21252 23964
rect 21308 23962 21314 23964
rect 21068 23910 21070 23962
rect 21250 23910 21252 23962
rect 21006 23908 21012 23910
rect 21068 23908 21092 23910
rect 21148 23908 21172 23910
rect 21228 23908 21252 23910
rect 21308 23908 21314 23910
rect 21006 23899 21314 23908
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20536 23588 20588 23594
rect 20536 23530 20588 23536
rect 20548 22574 20576 23530
rect 20916 22778 20944 23598
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21008 23254 21036 23462
rect 21468 23254 21496 24006
rect 21744 23662 21772 24346
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22100 24064 22152 24070
rect 22100 24006 22152 24012
rect 22112 23662 22140 24006
rect 21732 23656 21784 23662
rect 21560 23616 21732 23644
rect 20996 23248 21048 23254
rect 20996 23190 21048 23196
rect 21456 23248 21508 23254
rect 21456 23190 21508 23196
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21006 22876 21314 22885
rect 21006 22874 21012 22876
rect 21068 22874 21092 22876
rect 21148 22874 21172 22876
rect 21228 22874 21252 22876
rect 21308 22874 21314 22876
rect 21068 22822 21070 22874
rect 21250 22822 21252 22874
rect 21006 22820 21012 22822
rect 21068 22820 21092 22822
rect 21148 22820 21172 22822
rect 21228 22820 21252 22822
rect 21308 22820 21314 22822
rect 21006 22811 21314 22820
rect 21376 22778 21404 22918
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21560 22681 21588 23616
rect 21732 23598 21784 23604
rect 22100 23656 22152 23662
rect 22100 23598 22152 23604
rect 21666 23420 21974 23429
rect 21666 23418 21672 23420
rect 21728 23418 21752 23420
rect 21808 23418 21832 23420
rect 21888 23418 21912 23420
rect 21968 23418 21974 23420
rect 21728 23366 21730 23418
rect 21910 23366 21912 23418
rect 21666 23364 21672 23366
rect 21728 23364 21752 23366
rect 21808 23364 21832 23366
rect 21888 23364 21912 23366
rect 21968 23364 21974 23366
rect 21666 23355 21974 23364
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 21640 22704 21692 22710
rect 21546 22672 21602 22681
rect 21456 22636 21508 22642
rect 21640 22646 21692 22652
rect 21546 22607 21602 22616
rect 21456 22578 21508 22584
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20720 22568 20772 22574
rect 20720 22510 20772 22516
rect 20548 21486 20576 22510
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20640 21554 20668 21830
rect 20732 21690 20760 22510
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21376 22234 21404 22374
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20916 21690 20944 21966
rect 21006 21788 21314 21797
rect 21006 21786 21012 21788
rect 21068 21786 21092 21788
rect 21148 21786 21172 21788
rect 21228 21786 21252 21788
rect 21308 21786 21314 21788
rect 21068 21734 21070 21786
rect 21250 21734 21252 21786
rect 21006 21732 21012 21734
rect 21068 21732 21092 21734
rect 21148 21732 21172 21734
rect 21228 21732 21252 21734
rect 21308 21732 21314 21734
rect 21006 21723 21314 21732
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20536 21480 20588 21486
rect 20536 21422 20588 21428
rect 20640 21146 20668 21490
rect 21468 21350 21496 22578
rect 21560 22166 21588 22607
rect 21652 22545 21680 22646
rect 22112 22574 22140 23054
rect 22204 22778 22232 24142
rect 22296 23730 22324 25706
rect 22388 25498 22416 25706
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22480 25430 22508 26454
rect 23492 26450 23520 28630
rect 23768 28626 23796 29106
rect 23756 28620 23808 28626
rect 23756 28562 23808 28568
rect 23860 28218 23888 29294
rect 23940 28960 23992 28966
rect 23940 28902 23992 28908
rect 23952 28762 23980 28902
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 24032 28688 24084 28694
rect 24032 28630 24084 28636
rect 24044 28218 24072 28630
rect 23848 28212 23900 28218
rect 23848 28154 23900 28160
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 23584 27606 23612 27950
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23676 27470 23704 27950
rect 23940 27668 23992 27674
rect 23940 27610 23992 27616
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23572 27328 23624 27334
rect 23572 27270 23624 27276
rect 23584 27033 23612 27270
rect 23676 27130 23704 27406
rect 23664 27124 23716 27130
rect 23664 27066 23716 27072
rect 23570 27024 23626 27033
rect 23570 26959 23626 26968
rect 23584 26858 23612 26959
rect 23572 26852 23624 26858
rect 23572 26794 23624 26800
rect 23480 26444 23532 26450
rect 23480 26386 23532 26392
rect 23480 25832 23532 25838
rect 23480 25774 23532 25780
rect 22468 25424 22520 25430
rect 22468 25366 22520 25372
rect 22744 25288 22796 25294
rect 22744 25230 22796 25236
rect 22756 24750 22784 25230
rect 23492 24886 23520 25774
rect 23848 25696 23900 25702
rect 23848 25638 23900 25644
rect 23860 25498 23888 25638
rect 23848 25492 23900 25498
rect 23848 25434 23900 25440
rect 23952 25362 23980 27610
rect 24032 27600 24084 27606
rect 24032 27542 24084 27548
rect 24044 27402 24072 27542
rect 24032 27396 24084 27402
rect 24032 27338 24084 27344
rect 24136 26926 24164 31726
rect 24504 31470 24992 31498
rect 24504 31346 24532 31470
rect 24964 31414 24992 31470
rect 24584 31408 24636 31414
rect 24952 31408 25004 31414
rect 24636 31368 24716 31396
rect 24584 31350 24636 31356
rect 24492 31340 24544 31346
rect 24492 31282 24544 31288
rect 24688 31278 24716 31368
rect 24952 31350 25004 31356
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 25136 31272 25188 31278
rect 25136 31214 25188 31220
rect 24308 31204 24360 31210
rect 24308 31146 24360 31152
rect 24400 31204 24452 31210
rect 24400 31146 24452 31152
rect 24492 31204 24544 31210
rect 24492 31146 24544 31152
rect 24320 30870 24348 31146
rect 24308 30864 24360 30870
rect 24308 30806 24360 30812
rect 24412 30546 24440 31146
rect 24504 31113 24532 31146
rect 24490 31104 24546 31113
rect 24490 31039 24546 31048
rect 24596 30938 24624 31214
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24584 30932 24636 30938
rect 24584 30874 24636 30880
rect 24676 30864 24728 30870
rect 24676 30806 24728 30812
rect 24584 30592 24636 30598
rect 24412 30518 24532 30546
rect 24584 30534 24636 30540
rect 24400 30388 24452 30394
rect 24400 30330 24452 30336
rect 24412 29714 24440 30330
rect 24504 29850 24532 30518
rect 24596 30258 24624 30534
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 24492 29844 24544 29850
rect 24492 29786 24544 29792
rect 24688 29714 24716 30806
rect 24780 30802 24808 31078
rect 25148 30938 25176 31214
rect 25228 31136 25280 31142
rect 25226 31104 25228 31113
rect 25320 31136 25372 31142
rect 25280 31104 25282 31113
rect 25320 31078 25372 31084
rect 25226 31039 25282 31048
rect 25332 30954 25360 31078
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 25240 30926 25360 30954
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 24964 30394 24992 30874
rect 25044 30864 25096 30870
rect 25240 30818 25268 30926
rect 25096 30812 25268 30818
rect 25044 30806 25268 30812
rect 25056 30790 25268 30806
rect 25320 30796 25372 30802
rect 25320 30738 25372 30744
rect 25228 30728 25280 30734
rect 25228 30670 25280 30676
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 25240 30258 25268 30670
rect 25332 30394 25360 30738
rect 25320 30388 25372 30394
rect 25320 30330 25372 30336
rect 25228 30252 25280 30258
rect 25228 30194 25280 30200
rect 24768 29844 24820 29850
rect 25240 29832 25268 30194
rect 25516 30190 25544 31826
rect 25976 31822 26004 32234
rect 26436 31958 26464 33544
rect 28264 32224 28316 32230
rect 28264 32166 28316 32172
rect 26424 31952 26476 31958
rect 26424 31894 26476 31900
rect 28080 31952 28132 31958
rect 28080 31894 28132 31900
rect 25964 31816 26016 31822
rect 25964 31758 26016 31764
rect 25964 31680 26016 31686
rect 25964 31622 26016 31628
rect 25872 31408 25924 31414
rect 25872 31350 25924 31356
rect 25688 31272 25740 31278
rect 25688 31214 25740 31220
rect 25596 31204 25648 31210
rect 25596 31146 25648 31152
rect 25608 31113 25636 31146
rect 25594 31104 25650 31113
rect 25594 31039 25650 31048
rect 25700 30938 25728 31214
rect 25780 31136 25832 31142
rect 25780 31078 25832 31084
rect 25688 30932 25740 30938
rect 25688 30874 25740 30880
rect 25504 30184 25556 30190
rect 25792 30161 25820 31078
rect 25884 30802 25912 31350
rect 25872 30796 25924 30802
rect 25872 30738 25924 30744
rect 25884 30190 25912 30738
rect 25872 30184 25924 30190
rect 25504 30126 25556 30132
rect 25778 30152 25834 30161
rect 25872 30126 25924 30132
rect 25778 30087 25834 30096
rect 24768 29786 24820 29792
rect 25148 29804 25268 29832
rect 25688 29844 25740 29850
rect 24400 29708 24452 29714
rect 24400 29650 24452 29656
rect 24676 29708 24728 29714
rect 24676 29650 24728 29656
rect 24492 28144 24544 28150
rect 24492 28086 24544 28092
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 24308 27872 24360 27878
rect 24308 27814 24360 27820
rect 24320 27606 24348 27814
rect 24412 27674 24440 27950
rect 24400 27668 24452 27674
rect 24400 27610 24452 27616
rect 24308 27600 24360 27606
rect 24308 27542 24360 27548
rect 24216 27328 24268 27334
rect 24216 27270 24268 27276
rect 24228 27130 24256 27270
rect 24216 27124 24268 27130
rect 24216 27066 24268 27072
rect 24412 27033 24440 27610
rect 24504 27334 24532 28086
rect 24584 28008 24636 28014
rect 24584 27950 24636 27956
rect 24596 27470 24624 27950
rect 24584 27464 24636 27470
rect 24584 27406 24636 27412
rect 24492 27328 24544 27334
rect 24492 27270 24544 27276
rect 24584 27328 24636 27334
rect 24688 27282 24716 29650
rect 24780 29578 24808 29786
rect 24768 29572 24820 29578
rect 24768 29514 24820 29520
rect 24780 27674 24808 29514
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24964 29238 24992 29446
rect 24952 29232 25004 29238
rect 24952 29174 25004 29180
rect 25148 29170 25176 29804
rect 25884 29832 25912 30126
rect 25976 30122 26004 31622
rect 26332 31408 26384 31414
rect 26252 31368 26332 31396
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 26068 30852 26096 31282
rect 26252 30870 26280 31368
rect 26332 31350 26384 31356
rect 26332 31272 26384 31278
rect 26332 31214 26384 31220
rect 26424 31272 26476 31278
rect 26424 31214 26476 31220
rect 26884 31272 26936 31278
rect 26884 31214 26936 31220
rect 26240 30864 26292 30870
rect 26068 30824 26240 30852
rect 25964 30116 26016 30122
rect 25964 30058 26016 30064
rect 25740 29804 25912 29832
rect 25688 29786 25740 29792
rect 26068 29782 26096 30824
rect 26240 30806 26292 30812
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 26252 30274 26280 30534
rect 26160 30246 26280 30274
rect 26056 29776 26108 29782
rect 26056 29718 26108 29724
rect 25228 29708 25280 29714
rect 25228 29650 25280 29656
rect 25240 29170 25268 29650
rect 26068 29170 26096 29718
rect 26160 29510 26188 30246
rect 26344 29850 26372 31214
rect 26436 30938 26464 31214
rect 26516 31136 26568 31142
rect 26608 31136 26660 31142
rect 26516 31078 26568 31084
rect 26606 31104 26608 31113
rect 26660 31104 26662 31113
rect 26424 30932 26476 30938
rect 26424 30874 26476 30880
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26332 29844 26384 29850
rect 26332 29786 26384 29792
rect 26148 29504 26200 29510
rect 26148 29446 26200 29452
rect 26240 29504 26292 29510
rect 26240 29446 26292 29452
rect 25136 29164 25188 29170
rect 25136 29106 25188 29112
rect 25228 29164 25280 29170
rect 25228 29106 25280 29112
rect 26056 29164 26108 29170
rect 26056 29106 26108 29112
rect 25148 29034 25176 29106
rect 25136 29028 25188 29034
rect 25136 28970 25188 28976
rect 26056 28960 26108 28966
rect 26056 28902 26108 28908
rect 25136 28620 25188 28626
rect 25136 28562 25188 28568
rect 25148 28014 25176 28562
rect 26068 28082 26096 28902
rect 26160 28665 26188 29446
rect 26252 29306 26280 29446
rect 26240 29300 26292 29306
rect 26240 29242 26292 29248
rect 26436 28966 26464 30602
rect 26528 29170 26556 31078
rect 26606 31039 26662 31048
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26424 28960 26476 28966
rect 26424 28902 26476 28908
rect 26146 28656 26202 28665
rect 26146 28591 26202 28600
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 24768 27668 24820 27674
rect 24768 27610 24820 27616
rect 24952 27396 25004 27402
rect 24952 27338 25004 27344
rect 24636 27276 24716 27282
rect 24584 27270 24716 27276
rect 24398 27024 24454 27033
rect 24398 26959 24454 26968
rect 24504 26926 24532 27270
rect 24596 27254 24716 27270
rect 24124 26920 24176 26926
rect 24124 26862 24176 26868
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24492 26784 24544 26790
rect 24596 26738 24624 27254
rect 24860 26852 24912 26858
rect 24860 26794 24912 26800
rect 24544 26732 24624 26738
rect 24492 26726 24624 26732
rect 24504 26710 24624 26726
rect 24872 26246 24900 26794
rect 24964 26790 24992 27338
rect 25044 26852 25096 26858
rect 25044 26794 25096 26800
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24964 26314 24992 26726
rect 25056 26586 25084 26794
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24860 26240 24912 26246
rect 24860 26182 24912 26188
rect 24872 25362 24900 26182
rect 23940 25356 23992 25362
rect 23940 25298 23992 25304
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24964 25294 24992 26250
rect 25148 25922 25176 27950
rect 25596 27872 25648 27878
rect 25596 27814 25648 27820
rect 25872 27872 25924 27878
rect 25872 27814 25924 27820
rect 25608 27334 25636 27814
rect 25688 27668 25740 27674
rect 25688 27610 25740 27616
rect 25504 27328 25556 27334
rect 25504 27270 25556 27276
rect 25596 27328 25648 27334
rect 25596 27270 25648 27276
rect 25412 26920 25464 26926
rect 25412 26862 25464 26868
rect 25424 26586 25452 26862
rect 25412 26580 25464 26586
rect 25412 26522 25464 26528
rect 25228 26376 25280 26382
rect 25228 26318 25280 26324
rect 25240 26042 25268 26318
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 25148 25894 25268 25922
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 23480 24880 23532 24886
rect 23480 24822 23532 24828
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22744 24744 22796 24750
rect 22744 24686 22796 24692
rect 22664 24410 22692 24686
rect 22836 24608 22888 24614
rect 22836 24550 22888 24556
rect 24676 24608 24728 24614
rect 24676 24550 24728 24556
rect 22652 24404 22704 24410
rect 22652 24346 22704 24352
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22848 23118 22876 24550
rect 24124 24268 24176 24274
rect 24124 24210 24176 24216
rect 23940 24064 23992 24070
rect 23940 24006 23992 24012
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 23124 23118 23152 23666
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23204 22976 23256 22982
rect 23204 22918 23256 22924
rect 23216 22778 23244 22918
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 23204 22772 23256 22778
rect 23204 22714 23256 22720
rect 22100 22568 22152 22574
rect 21638 22536 21694 22545
rect 22100 22510 22152 22516
rect 21638 22471 21694 22480
rect 21666 22332 21974 22341
rect 21666 22330 21672 22332
rect 21728 22330 21752 22332
rect 21808 22330 21832 22332
rect 21888 22330 21912 22332
rect 21968 22330 21974 22332
rect 21728 22278 21730 22330
rect 21910 22278 21912 22330
rect 21666 22276 21672 22278
rect 21728 22276 21752 22278
rect 21808 22276 21832 22278
rect 21888 22276 21912 22278
rect 21968 22276 21974 22278
rect 21666 22267 21974 22276
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 21456 21344 21508 21350
rect 21456 21286 21508 21292
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 21560 21078 21588 22102
rect 22112 22030 22140 22510
rect 22204 22506 22232 22714
rect 22192 22500 22244 22506
rect 22192 22442 22244 22448
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22112 21350 22140 21966
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 22836 21412 22888 21418
rect 22836 21354 22888 21360
rect 22100 21344 22152 21350
rect 22100 21286 22152 21292
rect 21666 21244 21974 21253
rect 21666 21242 21672 21244
rect 21728 21242 21752 21244
rect 21808 21242 21832 21244
rect 21888 21242 21912 21244
rect 21968 21242 21974 21244
rect 21728 21190 21730 21242
rect 21910 21190 21912 21242
rect 21666 21188 21672 21190
rect 21728 21188 21752 21190
rect 21808 21188 21832 21190
rect 21888 21188 21912 21190
rect 21968 21188 21974 21190
rect 21666 21179 21974 21188
rect 20904 21072 20956 21078
rect 20904 21014 20956 21020
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 20812 21004 20864 21010
rect 20812 20946 20864 20952
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 20602 20760 20878
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20456 20420 20576 20448
rect 20442 20360 20498 20369
rect 20442 20295 20498 20304
rect 20456 20262 20484 20295
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 20456 20058 20484 20198
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 20260 19712 20312 19718
rect 20260 19654 20312 19660
rect 20076 18624 20128 18630
rect 20076 18566 20128 18572
rect 20088 18222 20116 18566
rect 20272 18222 20300 19654
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18766 20392 19110
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20442 18320 20498 18329
rect 20442 18255 20498 18264
rect 19800 18216 19852 18222
rect 19798 18184 19800 18193
rect 19984 18216 20036 18222
rect 19852 18184 19854 18193
rect 19984 18158 20036 18164
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 20260 18216 20312 18222
rect 20260 18158 20312 18164
rect 19798 18119 19854 18128
rect 20352 18148 20404 18154
rect 20352 18090 20404 18096
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 20088 16794 20116 17478
rect 20364 17066 20392 18090
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19996 16250 20024 16526
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 19800 16176 19852 16182
rect 19800 16118 19852 16124
rect 19812 15366 19840 16118
rect 19800 15360 19852 15366
rect 19800 15302 19852 15308
rect 19892 15360 19944 15366
rect 19892 15302 19944 15308
rect 19904 15026 19932 15302
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20364 14618 20392 14894
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20076 14272 20128 14278
rect 20074 14240 20076 14249
rect 20128 14240 20130 14249
rect 20074 14175 20130 14184
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 20088 12646 20116 13806
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20180 12442 20208 12650
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20456 12322 20484 18255
rect 20548 15502 20576 20420
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20640 18290 20668 19314
rect 20824 18465 20852 20946
rect 20916 20505 20944 21014
rect 22112 20874 22140 21286
rect 22100 20868 22152 20874
rect 22100 20810 22152 20816
rect 21006 20700 21314 20709
rect 21006 20698 21012 20700
rect 21068 20698 21092 20700
rect 21148 20698 21172 20700
rect 21228 20698 21252 20700
rect 21308 20698 21314 20700
rect 21068 20646 21070 20698
rect 21250 20646 21252 20698
rect 21006 20644 21012 20646
rect 21068 20644 21092 20646
rect 21148 20644 21172 20646
rect 21228 20644 21252 20646
rect 21308 20644 21314 20646
rect 21006 20635 21314 20644
rect 20902 20496 20958 20505
rect 22112 20466 22140 20810
rect 20902 20431 20958 20440
rect 21364 20460 21416 20466
rect 20916 19242 20944 20431
rect 21364 20402 21416 20408
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 20058 21128 20198
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 21006 19612 21314 19621
rect 21006 19610 21012 19612
rect 21068 19610 21092 19612
rect 21148 19610 21172 19612
rect 21228 19610 21252 19612
rect 21308 19610 21314 19612
rect 21068 19558 21070 19610
rect 21250 19558 21252 19610
rect 21006 19556 21012 19558
rect 21068 19556 21092 19558
rect 21148 19556 21172 19558
rect 21228 19556 21252 19558
rect 21308 19556 21314 19558
rect 21006 19547 21314 19556
rect 20904 19236 20956 19242
rect 20904 19178 20956 19184
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21088 18896 21140 18902
rect 21088 18838 21140 18844
rect 21100 18630 21128 18838
rect 21284 18714 21312 19110
rect 21376 18873 21404 20402
rect 22008 20324 22060 20330
rect 22008 20266 22060 20272
rect 21666 20156 21974 20165
rect 21666 20154 21672 20156
rect 21728 20154 21752 20156
rect 21808 20154 21832 20156
rect 21888 20154 21912 20156
rect 21968 20154 21974 20156
rect 21728 20102 21730 20154
rect 21910 20102 21912 20154
rect 21666 20100 21672 20102
rect 21728 20100 21752 20102
rect 21808 20100 21832 20102
rect 21888 20100 21912 20102
rect 21968 20100 21974 20102
rect 21666 20091 21974 20100
rect 22020 20058 22048 20266
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 21732 19848 21784 19854
rect 21732 19790 21784 19796
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21560 19174 21588 19654
rect 21744 19514 21772 19790
rect 21732 19508 21784 19514
rect 21732 19450 21784 19456
rect 21548 19168 21600 19174
rect 21548 19110 21600 19116
rect 21666 19068 21974 19077
rect 21666 19066 21672 19068
rect 21728 19066 21752 19068
rect 21808 19066 21832 19068
rect 21888 19066 21912 19068
rect 21968 19066 21974 19068
rect 21728 19014 21730 19066
rect 21910 19014 21912 19066
rect 21666 19012 21672 19014
rect 21728 19012 21752 19014
rect 21808 19012 21832 19014
rect 21888 19012 21912 19014
rect 21968 19012 21974 19014
rect 21666 19003 21974 19012
rect 21362 18864 21418 18873
rect 21362 18799 21418 18808
rect 21456 18760 21508 18766
rect 21362 18728 21418 18737
rect 21284 18686 21362 18714
rect 21456 18702 21508 18708
rect 21362 18663 21418 18672
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 21006 18524 21314 18533
rect 21006 18522 21012 18524
rect 21068 18522 21092 18524
rect 21148 18522 21172 18524
rect 21228 18522 21252 18524
rect 21308 18522 21314 18524
rect 21068 18470 21070 18522
rect 21250 18470 21252 18522
rect 21006 18468 21012 18470
rect 21068 18468 21092 18470
rect 21148 18468 21172 18470
rect 21228 18468 21252 18470
rect 21308 18468 21314 18470
rect 20810 18456 20866 18465
rect 21006 18459 21314 18468
rect 20810 18391 20866 18400
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20640 18193 20668 18226
rect 20626 18184 20682 18193
rect 20626 18119 20682 18128
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20640 17338 20668 17682
rect 21284 17678 21312 18022
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21006 17436 21314 17445
rect 21006 17434 21012 17436
rect 21068 17434 21092 17436
rect 21148 17434 21172 17436
rect 21228 17434 21252 17436
rect 21308 17434 21314 17436
rect 21068 17382 21070 17434
rect 21250 17382 21252 17434
rect 21006 17380 21012 17382
rect 21068 17380 21092 17382
rect 21148 17380 21172 17382
rect 21228 17380 21252 17382
rect 21308 17380 21314 17382
rect 21006 17371 21314 17380
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 21468 17134 21496 18702
rect 22008 18080 22060 18086
rect 22008 18022 22060 18028
rect 21666 17980 21974 17989
rect 21666 17978 21672 17980
rect 21728 17978 21752 17980
rect 21808 17978 21832 17980
rect 21888 17978 21912 17980
rect 21968 17978 21974 17980
rect 21728 17926 21730 17978
rect 21910 17926 21912 17978
rect 21666 17924 21672 17926
rect 21728 17924 21752 17926
rect 21808 17924 21832 17926
rect 21888 17924 21912 17926
rect 21968 17924 21974 17926
rect 21666 17915 21974 17924
rect 22020 17814 22048 18022
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 22112 17678 22140 20402
rect 22848 19922 22876 21354
rect 23308 21146 23336 21422
rect 23400 21418 23428 23530
rect 23480 23520 23532 23526
rect 23480 23462 23532 23468
rect 23492 22506 23520 23462
rect 23480 22500 23532 22506
rect 23480 22442 23532 22448
rect 23572 22160 23624 22166
rect 23572 22102 23624 22108
rect 23388 21412 23440 21418
rect 23388 21354 23440 21360
rect 23296 21140 23348 21146
rect 23296 21082 23348 21088
rect 23584 21010 23612 22102
rect 23952 22098 23980 24006
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24044 22234 24072 23054
rect 24032 22228 24084 22234
rect 24032 22170 24084 22176
rect 23940 22092 23992 22098
rect 23940 22034 23992 22040
rect 24136 21622 24164 24210
rect 24308 24200 24360 24206
rect 24308 24142 24360 24148
rect 24216 24132 24268 24138
rect 24216 24074 24268 24080
rect 24228 22234 24256 24074
rect 24320 22778 24348 24142
rect 24400 23520 24452 23526
rect 24400 23462 24452 23468
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 24412 22574 24440 23462
rect 24582 23352 24638 23361
rect 24582 23287 24638 23296
rect 24400 22568 24452 22574
rect 24400 22510 24452 22516
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 24596 22166 24624 23287
rect 24688 23186 24716 24550
rect 25148 24274 25176 25774
rect 25240 25362 25268 25894
rect 25320 25832 25372 25838
rect 25516 25786 25544 27270
rect 25700 26994 25728 27610
rect 25884 27062 25912 27814
rect 26068 27538 26096 28018
rect 26056 27532 26108 27538
rect 26056 27474 26108 27480
rect 26056 27328 26108 27334
rect 26056 27270 26108 27276
rect 25780 27056 25832 27062
rect 25778 27024 25780 27033
rect 25872 27056 25924 27062
rect 25832 27024 25834 27033
rect 25688 26988 25740 26994
rect 25872 26998 25924 27004
rect 25778 26959 25834 26968
rect 25688 26930 25740 26936
rect 25596 26784 25648 26790
rect 25596 26726 25648 26732
rect 25320 25774 25372 25780
rect 25332 25498 25360 25774
rect 25424 25758 25544 25786
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 25228 25356 25280 25362
rect 25228 25298 25280 25304
rect 25424 25226 25452 25758
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 25516 25362 25544 25638
rect 25608 25498 25636 26726
rect 25700 26602 25728 26930
rect 25700 26574 25820 26602
rect 25688 26512 25740 26518
rect 25688 26454 25740 26460
rect 25700 25498 25728 26454
rect 25596 25492 25648 25498
rect 25596 25434 25648 25440
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25504 25356 25556 25362
rect 25504 25298 25556 25304
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25516 24886 25544 25298
rect 25504 24880 25556 24886
rect 25504 24822 25556 24828
rect 25792 24614 25820 26574
rect 25884 25838 25912 26998
rect 25872 25832 25924 25838
rect 25872 25774 25924 25780
rect 25964 25492 26016 25498
rect 25964 25434 26016 25440
rect 25780 24608 25832 24614
rect 25832 24556 25912 24562
rect 25780 24550 25912 24556
rect 25792 24534 25912 24550
rect 25884 24274 25912 24534
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25412 24268 25464 24274
rect 25412 24210 25464 24216
rect 25596 24268 25648 24274
rect 25596 24210 25648 24216
rect 25872 24268 25924 24274
rect 25872 24210 25924 24216
rect 24860 24064 24912 24070
rect 24860 24006 24912 24012
rect 24952 24064 25004 24070
rect 24952 24006 25004 24012
rect 25136 24064 25188 24070
rect 25136 24006 25188 24012
rect 24872 23526 24900 24006
rect 24964 23594 24992 24006
rect 25148 23594 25176 24006
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 24952 23588 25004 23594
rect 24952 23530 25004 23536
rect 25136 23588 25188 23594
rect 25136 23530 25188 23536
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 25228 23316 25280 23322
rect 25228 23258 25280 23264
rect 24676 23180 24728 23186
rect 24676 23122 24728 23128
rect 24688 22778 24716 23122
rect 24952 23112 25004 23118
rect 25240 23066 25268 23258
rect 24952 23054 25004 23060
rect 24768 23044 24820 23050
rect 24768 22986 24820 22992
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24584 22160 24636 22166
rect 24676 22160 24728 22166
rect 24584 22102 24636 22108
rect 24674 22128 24676 22137
rect 24728 22128 24730 22137
rect 24674 22063 24730 22072
rect 24780 22030 24808 22986
rect 24860 22976 24912 22982
rect 24860 22918 24912 22924
rect 24492 22024 24544 22030
rect 24492 21966 24544 21972
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24504 21690 24532 21966
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24492 21684 24544 21690
rect 24492 21626 24544 21632
rect 24688 21622 24716 21830
rect 23756 21616 23808 21622
rect 23756 21558 23808 21564
rect 24124 21616 24176 21622
rect 24124 21558 24176 21564
rect 24676 21616 24728 21622
rect 24676 21558 24728 21564
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23020 20868 23072 20874
rect 23020 20810 23072 20816
rect 22928 20392 22980 20398
rect 22928 20334 22980 20340
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22744 19712 22796 19718
rect 22744 19654 22796 19660
rect 22756 19514 22784 19654
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22848 19334 22876 19858
rect 22940 19786 22968 20334
rect 23032 19922 23060 20810
rect 23388 20392 23440 20398
rect 23388 20334 23440 20340
rect 23020 19916 23072 19922
rect 23020 19858 23072 19864
rect 23204 19916 23256 19922
rect 23204 19858 23256 19864
rect 22928 19780 22980 19786
rect 22928 19722 22980 19728
rect 23216 19718 23244 19858
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 22756 19306 22876 19334
rect 22652 19236 22704 19242
rect 22652 19178 22704 19184
rect 22664 18970 22692 19178
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 22756 18834 22784 19306
rect 23400 18970 23428 20334
rect 23584 19922 23612 20946
rect 23768 20398 23796 21558
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24216 21344 24268 21350
rect 24216 21286 24268 21292
rect 24044 21010 24072 21286
rect 24228 21010 24256 21286
rect 24688 21146 24716 21558
rect 24676 21140 24728 21146
rect 24676 21082 24728 21088
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24216 21004 24268 21010
rect 24216 20946 24268 20952
rect 24400 21004 24452 21010
rect 24400 20946 24452 20952
rect 24584 21004 24636 21010
rect 24584 20946 24636 20952
rect 23940 20800 23992 20806
rect 23940 20742 23992 20748
rect 23952 20602 23980 20742
rect 23940 20596 23992 20602
rect 23940 20538 23992 20544
rect 24044 20466 24072 20946
rect 24124 20868 24176 20874
rect 24124 20810 24176 20816
rect 24136 20602 24164 20810
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 24032 20460 24084 20466
rect 24032 20402 24084 20408
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23848 20392 23900 20398
rect 23848 20334 23900 20340
rect 24124 20392 24176 20398
rect 24124 20334 24176 20340
rect 23664 20052 23716 20058
rect 23664 19994 23716 20000
rect 23572 19916 23624 19922
rect 23572 19858 23624 19864
rect 23676 19514 23704 19994
rect 23768 19689 23796 20334
rect 23860 20058 23888 20334
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 23848 20052 23900 20058
rect 23848 19994 23900 20000
rect 23952 19990 23980 20198
rect 23940 19984 23992 19990
rect 23940 19926 23992 19932
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23754 19680 23810 19689
rect 23754 19615 23810 19624
rect 23664 19508 23716 19514
rect 23664 19450 23716 19456
rect 23768 19394 23796 19615
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23676 19366 23796 19394
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 23492 18426 23520 19314
rect 23572 18624 23624 18630
rect 23572 18566 23624 18572
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22572 17882 22600 18158
rect 22836 18148 22888 18154
rect 22836 18090 22888 18096
rect 22848 17882 22876 18090
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 22560 17876 22612 17882
rect 22560 17818 22612 17824
rect 22836 17876 22888 17882
rect 22836 17818 22888 17824
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22112 17202 22140 17614
rect 22100 17196 22152 17202
rect 22100 17138 22152 17144
rect 21456 17128 21508 17134
rect 21456 17070 21508 17076
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21284 16794 21312 16934
rect 21666 16892 21974 16901
rect 21666 16890 21672 16892
rect 21728 16890 21752 16892
rect 21808 16890 21832 16892
rect 21888 16890 21912 16892
rect 21968 16890 21974 16892
rect 21728 16838 21730 16890
rect 21910 16838 21912 16890
rect 21666 16836 21672 16838
rect 21728 16836 21752 16838
rect 21808 16836 21832 16838
rect 21888 16836 21912 16838
rect 21968 16836 21974 16838
rect 21666 16827 21974 16836
rect 22848 16794 22876 17818
rect 23124 17134 23152 18022
rect 23584 17678 23612 18566
rect 23676 18426 23704 19366
rect 23756 19304 23808 19310
rect 23756 19246 23808 19252
rect 23768 18902 23796 19246
rect 23860 18970 23888 19790
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 23756 18896 23808 18902
rect 23756 18838 23808 18844
rect 23664 18420 23716 18426
rect 23664 18362 23716 18368
rect 23768 17678 23796 18838
rect 23952 18426 23980 19926
rect 24032 19508 24084 19514
rect 24032 19450 24084 19456
rect 24044 18834 24072 19450
rect 24136 18970 24164 20334
rect 24228 19786 24256 20946
rect 24412 20369 24440 20946
rect 24398 20360 24454 20369
rect 24398 20295 24454 20304
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24216 19780 24268 19786
rect 24216 19722 24268 19728
rect 24124 18964 24176 18970
rect 24124 18906 24176 18912
rect 24032 18828 24084 18834
rect 24032 18770 24084 18776
rect 23848 18420 23900 18426
rect 23848 18362 23900 18368
rect 23940 18420 23992 18426
rect 23940 18362 23992 18368
rect 23860 18222 23888 18362
rect 23848 18216 23900 18222
rect 23848 18158 23900 18164
rect 23860 17882 23888 18158
rect 23848 17876 23900 17882
rect 23848 17818 23900 17824
rect 24320 17814 24348 20198
rect 24596 20058 24624 20946
rect 24688 20466 24716 21082
rect 24780 21010 24808 21966
rect 24872 21010 24900 22918
rect 24964 21570 24992 23054
rect 25148 23038 25268 23066
rect 24964 21542 25084 21570
rect 25056 21486 25084 21542
rect 24952 21480 25004 21486
rect 24952 21422 25004 21428
rect 25044 21480 25096 21486
rect 25044 21422 25096 21428
rect 24964 21350 24992 21422
rect 24952 21344 25004 21350
rect 24952 21286 25004 21292
rect 24768 21004 24820 21010
rect 24768 20946 24820 20952
rect 24860 21004 24912 21010
rect 24860 20946 24912 20952
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 24584 20052 24636 20058
rect 24584 19994 24636 20000
rect 24596 19514 24624 19994
rect 24688 19514 24716 20198
rect 24780 19854 24808 20946
rect 24872 20398 24900 20946
rect 24964 20806 24992 21286
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 25056 20602 25084 21422
rect 25044 20596 25096 20602
rect 25044 20538 25096 20544
rect 25148 20466 25176 23038
rect 25228 22432 25280 22438
rect 25332 22409 25360 23802
rect 25424 22574 25452 24210
rect 25504 23724 25556 23730
rect 25504 23666 25556 23672
rect 25516 23633 25544 23666
rect 25502 23624 25558 23633
rect 25502 23559 25558 23568
rect 25608 23322 25636 24210
rect 25688 23724 25740 23730
rect 25688 23666 25740 23672
rect 25596 23316 25648 23322
rect 25596 23258 25648 23264
rect 25504 23248 25556 23254
rect 25504 23190 25556 23196
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25228 22374 25280 22380
rect 25318 22400 25374 22409
rect 25240 22030 25268 22374
rect 25318 22335 25374 22344
rect 25332 22080 25360 22335
rect 25424 22234 25452 22510
rect 25412 22228 25464 22234
rect 25412 22170 25464 22176
rect 25412 22092 25464 22098
rect 25332 22052 25412 22080
rect 25516 22094 25544 23190
rect 25700 22574 25728 23666
rect 25780 23520 25832 23526
rect 25832 23480 25912 23508
rect 25780 23462 25832 23468
rect 25884 23186 25912 23480
rect 25872 23180 25924 23186
rect 25872 23122 25924 23128
rect 25780 22976 25832 22982
rect 25884 22964 25912 23122
rect 25976 23050 26004 25434
rect 26068 25362 26096 27270
rect 26160 26790 26188 28591
rect 26436 28422 26464 28902
rect 26424 28416 26476 28422
rect 26424 28358 26476 28364
rect 26620 28218 26648 31039
rect 26792 30728 26844 30734
rect 26792 30670 26844 30676
rect 26804 29306 26832 30670
rect 26896 30394 26924 31214
rect 27160 31136 27212 31142
rect 27160 31078 27212 31084
rect 26884 30388 26936 30394
rect 26884 30330 26936 30336
rect 27172 30258 27200 31078
rect 27620 30932 27672 30938
rect 27620 30874 27672 30880
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27068 30252 27120 30258
rect 27068 30194 27120 30200
rect 27160 30252 27212 30258
rect 27160 30194 27212 30200
rect 26974 30152 27030 30161
rect 26974 30087 27030 30096
rect 27080 30138 27108 30194
rect 27080 30110 27292 30138
rect 26792 29300 26844 29306
rect 26792 29242 26844 29248
rect 26884 28960 26936 28966
rect 26884 28902 26936 28908
rect 26608 28212 26660 28218
rect 26528 28172 26608 28200
rect 26424 27940 26476 27946
rect 26424 27882 26476 27888
rect 26436 27606 26464 27882
rect 26424 27600 26476 27606
rect 26424 27542 26476 27548
rect 26332 27328 26384 27334
rect 26332 27270 26384 27276
rect 26344 27130 26372 27270
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26148 26784 26200 26790
rect 26148 26726 26200 26732
rect 26332 26784 26384 26790
rect 26332 26726 26384 26732
rect 26344 26518 26372 26726
rect 26332 26512 26384 26518
rect 26332 26454 26384 26460
rect 26436 26314 26464 27542
rect 26528 26518 26556 28172
rect 26608 28154 26660 28160
rect 26896 28014 26924 28902
rect 26988 28558 27016 30087
rect 27080 28762 27108 30110
rect 27264 30054 27292 30110
rect 27160 30048 27212 30054
rect 27160 29990 27212 29996
rect 27252 30048 27304 30054
rect 27252 29990 27304 29996
rect 27172 29578 27200 29990
rect 27160 29572 27212 29578
rect 27160 29514 27212 29520
rect 27540 29306 27568 30330
rect 27632 29306 27660 30874
rect 27896 30184 27948 30190
rect 27896 30126 27948 30132
rect 27908 29850 27936 30126
rect 27896 29844 27948 29850
rect 27896 29786 27948 29792
rect 28092 29730 28120 31894
rect 28172 30932 28224 30938
rect 28172 30874 28224 30880
rect 27908 29702 28120 29730
rect 27528 29300 27580 29306
rect 27528 29242 27580 29248
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 27540 28762 27568 29242
rect 27620 29096 27672 29102
rect 27620 29038 27672 29044
rect 27068 28756 27120 28762
rect 27068 28698 27120 28704
rect 27528 28756 27580 28762
rect 27528 28698 27580 28704
rect 27528 28620 27580 28626
rect 27632 28608 27660 29038
rect 27908 29034 27936 29702
rect 27988 29640 28040 29646
rect 27988 29582 28040 29588
rect 28000 29102 28028 29582
rect 28184 29170 28212 30874
rect 28276 30802 28304 32166
rect 28368 31822 28396 33544
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28644 31890 28672 32166
rect 29026 32124 29334 32133
rect 29026 32122 29032 32124
rect 29088 32122 29112 32124
rect 29168 32122 29192 32124
rect 29248 32122 29272 32124
rect 29328 32122 29334 32124
rect 29088 32070 29090 32122
rect 29270 32070 29272 32122
rect 29026 32068 29032 32070
rect 29088 32068 29112 32070
rect 29168 32068 29192 32070
rect 29248 32068 29272 32070
rect 29328 32068 29334 32070
rect 29026 32059 29334 32068
rect 28632 31884 28684 31890
rect 28632 31826 28684 31832
rect 28724 31884 28776 31890
rect 28724 31826 28776 31832
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 28366 31580 28674 31589
rect 28366 31578 28372 31580
rect 28428 31578 28452 31580
rect 28508 31578 28532 31580
rect 28588 31578 28612 31580
rect 28668 31578 28674 31580
rect 28428 31526 28430 31578
rect 28610 31526 28612 31578
rect 28366 31524 28372 31526
rect 28428 31524 28452 31526
rect 28508 31524 28532 31526
rect 28588 31524 28612 31526
rect 28668 31524 28674 31526
rect 28366 31515 28674 31524
rect 28736 30938 28764 31826
rect 29932 31754 29960 33646
rect 31574 33544 31630 34344
rect 32862 33674 32918 34344
rect 32600 33646 32918 33674
rect 31024 32020 31076 32026
rect 31024 31962 31076 31968
rect 29932 31726 30144 31754
rect 29642 31376 29698 31385
rect 30116 31346 30144 31726
rect 29642 31311 29698 31320
rect 30104 31340 30156 31346
rect 29656 31278 29684 31311
rect 30104 31282 30156 31288
rect 29644 31272 29696 31278
rect 29644 31214 29696 31220
rect 29026 31036 29334 31045
rect 29026 31034 29032 31036
rect 29088 31034 29112 31036
rect 29168 31034 29192 31036
rect 29248 31034 29272 31036
rect 29328 31034 29334 31036
rect 29088 30982 29090 31034
rect 29270 30982 29272 31034
rect 29026 30980 29032 30982
rect 29088 30980 29112 30982
rect 29168 30980 29192 30982
rect 29248 30980 29272 30982
rect 29328 30980 29334 30982
rect 29026 30971 29334 30980
rect 28724 30932 28776 30938
rect 28724 30874 28776 30880
rect 28264 30796 28316 30802
rect 28264 30738 28316 30744
rect 28816 30796 28868 30802
rect 28816 30738 28868 30744
rect 29828 30796 29880 30802
rect 29828 30738 29880 30744
rect 30380 30796 30432 30802
rect 30380 30738 30432 30744
rect 28724 30592 28776 30598
rect 28724 30534 28776 30540
rect 28366 30492 28674 30501
rect 28366 30490 28372 30492
rect 28428 30490 28452 30492
rect 28508 30490 28532 30492
rect 28588 30490 28612 30492
rect 28668 30490 28674 30492
rect 28428 30438 28430 30490
rect 28610 30438 28612 30490
rect 28366 30436 28372 30438
rect 28428 30436 28452 30438
rect 28508 30436 28532 30438
rect 28588 30436 28612 30438
rect 28668 30436 28674 30438
rect 28366 30427 28674 30436
rect 28264 30184 28316 30190
rect 28264 30126 28316 30132
rect 28276 29306 28304 30126
rect 28356 30116 28408 30122
rect 28356 30058 28408 30064
rect 28368 29646 28396 30058
rect 28736 29782 28764 30534
rect 28828 30394 28856 30738
rect 29736 30728 29788 30734
rect 29736 30670 29788 30676
rect 28816 30388 28868 30394
rect 28816 30330 28868 30336
rect 28724 29776 28776 29782
rect 28724 29718 28776 29724
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 28366 29404 28674 29413
rect 28366 29402 28372 29404
rect 28428 29402 28452 29404
rect 28508 29402 28532 29404
rect 28588 29402 28612 29404
rect 28668 29402 28674 29404
rect 28428 29350 28430 29402
rect 28610 29350 28612 29402
rect 28366 29348 28372 29350
rect 28428 29348 28452 29350
rect 28508 29348 28532 29350
rect 28588 29348 28612 29350
rect 28668 29348 28674 29350
rect 28366 29339 28674 29348
rect 28264 29300 28316 29306
rect 28264 29242 28316 29248
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 27988 29096 28040 29102
rect 27988 29038 28040 29044
rect 28632 29096 28684 29102
rect 28632 29038 28684 29044
rect 27896 29028 27948 29034
rect 27896 28970 27948 28976
rect 27908 28626 27936 28970
rect 27580 28580 27660 28608
rect 27528 28562 27580 28568
rect 26976 28552 27028 28558
rect 26976 28494 27028 28500
rect 27436 28484 27488 28490
rect 27436 28426 27488 28432
rect 26700 28008 26752 28014
rect 26700 27950 26752 27956
rect 26884 28008 26936 28014
rect 26884 27950 26936 27956
rect 26608 27328 26660 27334
rect 26608 27270 26660 27276
rect 26620 26518 26648 27270
rect 26516 26512 26568 26518
rect 26516 26454 26568 26460
rect 26608 26512 26660 26518
rect 26608 26454 26660 26460
rect 26424 26308 26476 26314
rect 26424 26250 26476 26256
rect 26332 25832 26384 25838
rect 26332 25774 26384 25780
rect 26056 25356 26108 25362
rect 26056 25298 26108 25304
rect 26344 25294 26372 25774
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26332 25288 26384 25294
rect 26332 25230 26384 25236
rect 26620 24274 26648 25638
rect 26712 25498 26740 27950
rect 26896 27674 26924 27950
rect 27252 27940 27304 27946
rect 27252 27882 27304 27888
rect 26976 27872 27028 27878
rect 26976 27814 27028 27820
rect 26884 27668 26936 27674
rect 26884 27610 26936 27616
rect 26884 27464 26936 27470
rect 26884 27406 26936 27412
rect 26792 27396 26844 27402
rect 26792 27338 26844 27344
rect 26804 26518 26832 27338
rect 26896 26586 26924 27406
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 26792 26512 26844 26518
rect 26792 26454 26844 26460
rect 26988 26382 27016 27814
rect 27264 27588 27292 27882
rect 27344 27600 27396 27606
rect 27264 27560 27344 27588
rect 27344 27542 27396 27548
rect 27356 26790 27384 27542
rect 27448 27402 27476 28426
rect 27632 28150 27660 28580
rect 27712 28620 27764 28626
rect 27896 28620 27948 28626
rect 27764 28580 27844 28608
rect 27712 28562 27764 28568
rect 27816 28506 27844 28580
rect 27896 28562 27948 28568
rect 28000 28506 28028 29038
rect 28644 28762 28672 29038
rect 28828 28994 28856 30330
rect 28908 30184 28960 30190
rect 28908 30126 28960 30132
rect 28920 29102 28948 30126
rect 29368 30048 29420 30054
rect 29368 29990 29420 29996
rect 29552 30048 29604 30054
rect 29552 29990 29604 29996
rect 29026 29948 29334 29957
rect 29026 29946 29032 29948
rect 29088 29946 29112 29948
rect 29168 29946 29192 29948
rect 29248 29946 29272 29948
rect 29328 29946 29334 29948
rect 29088 29894 29090 29946
rect 29270 29894 29272 29946
rect 29026 29892 29032 29894
rect 29088 29892 29112 29894
rect 29168 29892 29192 29894
rect 29248 29892 29272 29894
rect 29328 29892 29334 29894
rect 29026 29883 29334 29892
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 29276 29844 29328 29850
rect 29276 29786 29328 29792
rect 29012 29306 29040 29786
rect 29184 29708 29236 29714
rect 29184 29650 29236 29656
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 28908 29096 28960 29102
rect 28908 29038 28960 29044
rect 28736 28966 28856 28994
rect 28632 28756 28684 28762
rect 28632 28698 28684 28704
rect 27816 28478 28028 28506
rect 28172 28552 28224 28558
rect 28172 28494 28224 28500
rect 27620 28144 27672 28150
rect 27620 28086 27672 28092
rect 27620 28008 27672 28014
rect 27620 27950 27672 27956
rect 27528 27940 27580 27946
rect 27528 27882 27580 27888
rect 27436 27396 27488 27402
rect 27436 27338 27488 27344
rect 27540 27033 27568 27882
rect 27632 27538 27660 27950
rect 27816 27878 27844 28478
rect 27896 28076 27948 28082
rect 27896 28018 27948 28024
rect 27804 27872 27856 27878
rect 27804 27814 27856 27820
rect 27620 27532 27672 27538
rect 27620 27474 27672 27480
rect 27526 27024 27582 27033
rect 27526 26959 27582 26968
rect 27344 26784 27396 26790
rect 27344 26726 27396 26732
rect 27356 26586 27384 26726
rect 27540 26586 27568 26959
rect 27344 26580 27396 26586
rect 27344 26522 27396 26528
rect 27528 26580 27580 26586
rect 27528 26522 27580 26528
rect 27816 26450 27844 27814
rect 27908 26926 27936 28018
rect 28184 27946 28212 28494
rect 28366 28316 28674 28325
rect 28366 28314 28372 28316
rect 28428 28314 28452 28316
rect 28508 28314 28532 28316
rect 28588 28314 28612 28316
rect 28668 28314 28674 28316
rect 28428 28262 28430 28314
rect 28610 28262 28612 28314
rect 28366 28260 28372 28262
rect 28428 28260 28452 28262
rect 28508 28260 28532 28262
rect 28588 28260 28612 28262
rect 28668 28260 28674 28262
rect 28366 28251 28674 28260
rect 28736 28218 28764 28966
rect 28920 28665 28948 29038
rect 29196 28994 29224 29650
rect 29288 29510 29316 29786
rect 29276 29504 29328 29510
rect 29276 29446 29328 29452
rect 29380 29306 29408 29990
rect 29564 29510 29592 29990
rect 29748 29850 29776 30670
rect 29736 29844 29788 29850
rect 29736 29786 29788 29792
rect 29552 29504 29604 29510
rect 29552 29446 29604 29452
rect 29368 29300 29420 29306
rect 29368 29242 29420 29248
rect 29196 28966 29500 28994
rect 29026 28860 29334 28869
rect 29026 28858 29032 28860
rect 29088 28858 29112 28860
rect 29168 28858 29192 28860
rect 29248 28858 29272 28860
rect 29328 28858 29334 28860
rect 29088 28806 29090 28858
rect 29270 28806 29272 28858
rect 29026 28804 29032 28806
rect 29088 28804 29112 28806
rect 29168 28804 29192 28806
rect 29248 28804 29272 28806
rect 29328 28804 29334 28806
rect 29026 28795 29334 28804
rect 28906 28656 28962 28665
rect 28816 28620 28868 28626
rect 28906 28591 28962 28600
rect 28816 28562 28868 28568
rect 28828 28218 28856 28562
rect 28920 28558 28948 28591
rect 28908 28552 28960 28558
rect 28908 28494 28960 28500
rect 28540 28212 28592 28218
rect 28540 28154 28592 28160
rect 28724 28212 28776 28218
rect 28724 28154 28776 28160
rect 28816 28212 28868 28218
rect 28816 28154 28868 28160
rect 28264 28144 28316 28150
rect 28264 28086 28316 28092
rect 28172 27940 28224 27946
rect 28172 27882 28224 27888
rect 28184 27674 28212 27882
rect 28172 27668 28224 27674
rect 28172 27610 28224 27616
rect 28184 27538 28212 27610
rect 28172 27532 28224 27538
rect 28172 27474 28224 27480
rect 27988 27464 28040 27470
rect 27988 27406 28040 27412
rect 28000 27130 28028 27406
rect 27988 27124 28040 27130
rect 27988 27066 28040 27072
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27804 26444 27856 26450
rect 27804 26386 27856 26392
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 27712 26308 27764 26314
rect 27712 26250 27764 26256
rect 26700 25492 26752 25498
rect 26700 25434 26752 25440
rect 27724 24818 27752 26250
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 26700 24404 26752 24410
rect 26700 24346 26752 24352
rect 26240 24268 26292 24274
rect 26240 24210 26292 24216
rect 26608 24268 26660 24274
rect 26608 24210 26660 24216
rect 26056 23520 26108 23526
rect 26056 23462 26108 23468
rect 26068 23361 26096 23462
rect 26054 23352 26110 23361
rect 26252 23322 26280 24210
rect 26424 23792 26476 23798
rect 26476 23752 26556 23780
rect 26424 23734 26476 23740
rect 26332 23656 26384 23662
rect 26332 23598 26384 23604
rect 26424 23656 26476 23662
rect 26424 23598 26476 23604
rect 26054 23287 26110 23296
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 26056 23248 26108 23254
rect 26056 23190 26108 23196
rect 25964 23044 26016 23050
rect 25964 22986 26016 22992
rect 25832 22936 25912 22964
rect 25780 22918 25832 22924
rect 26068 22778 26096 23190
rect 26252 23050 26280 23258
rect 26344 23050 26372 23598
rect 26240 23044 26292 23050
rect 26240 22986 26292 22992
rect 26332 23044 26384 23050
rect 26332 22986 26384 22992
rect 26056 22772 26108 22778
rect 26056 22714 26108 22720
rect 26054 22672 26110 22681
rect 26054 22607 26110 22616
rect 26068 22574 26096 22607
rect 25688 22568 25740 22574
rect 25688 22510 25740 22516
rect 26056 22568 26108 22574
rect 26056 22510 26108 22516
rect 25516 22066 25636 22094
rect 25412 22034 25464 22040
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25240 21622 25268 21966
rect 25228 21616 25280 21622
rect 25228 21558 25280 21564
rect 25424 21350 25452 22034
rect 25504 21956 25556 21962
rect 25504 21898 25556 21904
rect 25412 21344 25464 21350
rect 25412 21286 25464 21292
rect 25516 21078 25544 21898
rect 25504 21072 25556 21078
rect 25504 21014 25556 21020
rect 25320 20936 25372 20942
rect 25320 20878 25372 20884
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24860 20392 24912 20398
rect 24860 20334 24912 20340
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 25136 19712 25188 19718
rect 25332 19689 25360 20878
rect 25516 20602 25544 20878
rect 25608 20602 25636 22066
rect 25872 22092 25924 22098
rect 25872 22034 25924 22040
rect 25780 21888 25832 21894
rect 25780 21830 25832 21836
rect 25688 21412 25740 21418
rect 25688 21354 25740 21360
rect 25700 21010 25728 21354
rect 25792 21162 25820 21830
rect 25884 21418 25912 22034
rect 26068 21894 26096 22510
rect 26344 22506 26372 22986
rect 26436 22658 26464 23598
rect 26528 22760 26556 23752
rect 26620 23186 26648 24210
rect 26712 23866 26740 24346
rect 26700 23860 26752 23866
rect 26700 23802 26752 23808
rect 26712 23662 26740 23802
rect 27816 23662 27844 26386
rect 27908 25770 27936 26726
rect 28276 26450 28304 28086
rect 28552 27538 28580 28154
rect 28724 28076 28776 28082
rect 28724 28018 28776 28024
rect 28632 28008 28684 28014
rect 28632 27950 28684 27956
rect 28540 27532 28592 27538
rect 28540 27474 28592 27480
rect 28644 27470 28672 27950
rect 28736 27860 28764 28018
rect 28816 27872 28868 27878
rect 28736 27832 28816 27860
rect 28816 27814 28868 27820
rect 28632 27464 28684 27470
rect 28920 27418 28948 28494
rect 29184 28484 29236 28490
rect 29184 28426 29236 28432
rect 29196 28150 29224 28426
rect 29472 28218 29500 28966
rect 29564 28694 29592 29446
rect 29552 28688 29604 28694
rect 29552 28630 29604 28636
rect 29460 28212 29512 28218
rect 29460 28154 29512 28160
rect 29184 28144 29236 28150
rect 29184 28086 29236 28092
rect 29458 28112 29514 28121
rect 29368 28076 29420 28082
rect 29458 28047 29514 28056
rect 29368 28018 29420 28024
rect 29380 27985 29408 28018
rect 29366 27976 29422 27985
rect 29472 27946 29500 28047
rect 29366 27911 29422 27920
rect 29460 27940 29512 27946
rect 29460 27882 29512 27888
rect 29026 27772 29334 27781
rect 29026 27770 29032 27772
rect 29088 27770 29112 27772
rect 29168 27770 29192 27772
rect 29248 27770 29272 27772
rect 29328 27770 29334 27772
rect 29088 27718 29090 27770
rect 29270 27718 29272 27770
rect 29026 27716 29032 27718
rect 29088 27716 29112 27718
rect 29168 27716 29192 27718
rect 29248 27716 29272 27718
rect 29328 27716 29334 27718
rect 29026 27707 29334 27716
rect 29564 27538 29592 28630
rect 29644 28144 29696 28150
rect 29644 28086 29696 28092
rect 29000 27532 29052 27538
rect 29000 27474 29052 27480
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 28632 27406 28684 27412
rect 28736 27390 28948 27418
rect 28366 27228 28674 27237
rect 28366 27226 28372 27228
rect 28428 27226 28452 27228
rect 28508 27226 28532 27228
rect 28588 27226 28612 27228
rect 28668 27226 28674 27228
rect 28428 27174 28430 27226
rect 28610 27174 28612 27226
rect 28366 27172 28372 27174
rect 28428 27172 28452 27174
rect 28508 27172 28532 27174
rect 28588 27172 28612 27174
rect 28668 27172 28674 27174
rect 28366 27163 28674 27172
rect 28736 27112 28764 27390
rect 28908 27328 28960 27334
rect 28908 27270 28960 27276
rect 28644 27084 28764 27112
rect 28448 26920 28500 26926
rect 28448 26862 28500 26868
rect 28460 26586 28488 26862
rect 28448 26580 28500 26586
rect 28448 26522 28500 26528
rect 28644 26450 28672 27084
rect 28920 27062 28948 27270
rect 28908 27056 28960 27062
rect 28908 26998 28960 27004
rect 29012 26874 29040 27474
rect 29550 27432 29606 27441
rect 29550 27367 29552 27376
rect 29604 27367 29606 27376
rect 29552 27338 29604 27344
rect 28828 26846 29040 26874
rect 28828 26450 28856 26846
rect 29368 26784 29420 26790
rect 29368 26726 29420 26732
rect 29460 26784 29512 26790
rect 29460 26726 29512 26732
rect 29026 26684 29334 26693
rect 29026 26682 29032 26684
rect 29088 26682 29112 26684
rect 29168 26682 29192 26684
rect 29248 26682 29272 26684
rect 29328 26682 29334 26684
rect 29088 26630 29090 26682
rect 29270 26630 29272 26682
rect 29026 26628 29032 26630
rect 29088 26628 29112 26630
rect 29168 26628 29192 26630
rect 29248 26628 29272 26630
rect 29328 26628 29334 26630
rect 29026 26619 29334 26628
rect 29092 26512 29144 26518
rect 29092 26454 29144 26460
rect 28264 26444 28316 26450
rect 28264 26386 28316 26392
rect 28632 26444 28684 26450
rect 28632 26386 28684 26392
rect 28816 26444 28868 26450
rect 28816 26386 28868 26392
rect 28172 26376 28224 26382
rect 28172 26318 28224 26324
rect 28184 25906 28212 26318
rect 28816 26240 28868 26246
rect 28816 26182 28868 26188
rect 28908 26240 28960 26246
rect 28908 26182 28960 26188
rect 28366 26140 28674 26149
rect 28366 26138 28372 26140
rect 28428 26138 28452 26140
rect 28508 26138 28532 26140
rect 28588 26138 28612 26140
rect 28668 26138 28674 26140
rect 28428 26086 28430 26138
rect 28610 26086 28612 26138
rect 28366 26084 28372 26086
rect 28428 26084 28452 26086
rect 28508 26084 28532 26086
rect 28588 26084 28612 26086
rect 28668 26084 28674 26086
rect 28366 26075 28674 26084
rect 28172 25900 28224 25906
rect 28224 25860 28304 25888
rect 28172 25842 28224 25848
rect 27896 25764 27948 25770
rect 27896 25706 27948 25712
rect 27896 25492 27948 25498
rect 27896 25434 27948 25440
rect 27908 24954 27936 25434
rect 28172 25220 28224 25226
rect 28172 25162 28224 25168
rect 27988 25152 28040 25158
rect 27988 25094 28040 25100
rect 28000 24954 28028 25094
rect 28184 24954 28212 25162
rect 27896 24948 27948 24954
rect 27896 24890 27948 24896
rect 27988 24948 28040 24954
rect 27988 24890 28040 24896
rect 28172 24948 28224 24954
rect 28172 24890 28224 24896
rect 28276 24818 28304 25860
rect 28828 25838 28856 26182
rect 28920 25974 28948 26182
rect 28908 25968 28960 25974
rect 28908 25910 28960 25916
rect 28816 25832 28868 25838
rect 28816 25774 28868 25780
rect 29104 25702 29132 26454
rect 29380 26042 29408 26726
rect 29472 26586 29500 26726
rect 29460 26580 29512 26586
rect 29460 26522 29512 26528
rect 29368 26036 29420 26042
rect 29368 25978 29420 25984
rect 29092 25696 29144 25702
rect 29092 25638 29144 25644
rect 29026 25596 29334 25605
rect 29026 25594 29032 25596
rect 29088 25594 29112 25596
rect 29168 25594 29192 25596
rect 29248 25594 29272 25596
rect 29328 25594 29334 25596
rect 29088 25542 29090 25594
rect 29270 25542 29272 25594
rect 29026 25540 29032 25542
rect 29088 25540 29112 25542
rect 29168 25540 29192 25542
rect 29248 25540 29272 25542
rect 29328 25540 29334 25542
rect 29026 25531 29334 25540
rect 29380 25362 29408 25978
rect 29368 25356 29420 25362
rect 29368 25298 29420 25304
rect 29184 25152 29236 25158
rect 29184 25094 29236 25100
rect 28366 25052 28674 25061
rect 28366 25050 28372 25052
rect 28428 25050 28452 25052
rect 28508 25050 28532 25052
rect 28588 25050 28612 25052
rect 28668 25050 28674 25052
rect 28428 24998 28430 25050
rect 28610 24998 28612 25050
rect 28366 24996 28372 24998
rect 28428 24996 28452 24998
rect 28508 24996 28532 24998
rect 28588 24996 28612 24998
rect 28668 24996 28674 24998
rect 28366 24987 28674 24996
rect 28264 24812 28316 24818
rect 28264 24754 28316 24760
rect 27896 24744 27948 24750
rect 27896 24686 27948 24692
rect 27988 24744 28040 24750
rect 27988 24686 28040 24692
rect 27908 24342 27936 24686
rect 27896 24336 27948 24342
rect 27896 24278 27948 24284
rect 26700 23656 26752 23662
rect 26884 23656 26936 23662
rect 26700 23598 26752 23604
rect 26790 23624 26846 23633
rect 26884 23598 26936 23604
rect 27804 23656 27856 23662
rect 27804 23598 27856 23604
rect 26790 23559 26846 23568
rect 26608 23180 26660 23186
rect 26608 23122 26660 23128
rect 26700 23180 26752 23186
rect 26700 23122 26752 23128
rect 26528 22732 26648 22760
rect 26436 22630 26556 22658
rect 26424 22568 26476 22574
rect 26424 22510 26476 22516
rect 26332 22500 26384 22506
rect 26332 22442 26384 22448
rect 26332 22024 26384 22030
rect 26332 21966 26384 21972
rect 26056 21888 26108 21894
rect 26056 21830 26108 21836
rect 26068 21690 26096 21830
rect 26056 21684 26108 21690
rect 26056 21626 26108 21632
rect 26148 21548 26200 21554
rect 26148 21490 26200 21496
rect 25872 21412 25924 21418
rect 25872 21354 25924 21360
rect 25792 21134 26004 21162
rect 25976 21026 26004 21134
rect 25688 21004 25740 21010
rect 25976 20998 26096 21026
rect 25688 20946 25740 20952
rect 25700 20890 25728 20946
rect 26068 20942 26096 20998
rect 26160 20942 26188 21490
rect 26344 21434 26372 21966
rect 26436 21554 26464 22510
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26344 21406 26464 21434
rect 26056 20936 26108 20942
rect 25700 20862 25820 20890
rect 26056 20878 26108 20884
rect 26148 20936 26200 20942
rect 26148 20878 26200 20884
rect 25688 20800 25740 20806
rect 25688 20742 25740 20748
rect 25700 20602 25728 20742
rect 25504 20596 25556 20602
rect 25504 20538 25556 20544
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25688 20596 25740 20602
rect 25688 20538 25740 20544
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 25136 19654 25188 19660
rect 25318 19680 25374 19689
rect 24780 19514 24808 19654
rect 24584 19508 24636 19514
rect 24504 19468 24584 19496
rect 24400 19168 24452 19174
rect 24400 19110 24452 19116
rect 24412 18426 24440 19110
rect 24400 18420 24452 18426
rect 24400 18362 24452 18368
rect 24504 18222 24532 19468
rect 24584 19450 24636 19456
rect 24676 19508 24728 19514
rect 24676 19450 24728 19456
rect 24768 19508 24820 19514
rect 24768 19450 24820 19456
rect 24584 19168 24636 19174
rect 24584 19110 24636 19116
rect 24596 18426 24624 19110
rect 24688 18834 24716 19450
rect 24780 18834 24808 19450
rect 25148 18902 25176 19654
rect 25318 19615 25374 19624
rect 25332 19394 25360 19615
rect 25516 19446 25544 20402
rect 25792 20398 25820 20862
rect 26436 20806 26464 21406
rect 26528 21350 26556 22630
rect 26620 22250 26648 22732
rect 26712 22545 26740 23122
rect 26804 23050 26832 23559
rect 26896 23186 26924 23598
rect 27344 23520 27396 23526
rect 27344 23462 27396 23468
rect 27250 23352 27306 23361
rect 27250 23287 27306 23296
rect 26884 23180 26936 23186
rect 26884 23122 26936 23128
rect 26792 23044 26844 23050
rect 26792 22986 26844 22992
rect 26804 22574 26832 22986
rect 26792 22568 26844 22574
rect 26698 22536 26754 22545
rect 26792 22510 26844 22516
rect 26698 22471 26754 22480
rect 27264 22438 27292 23287
rect 27160 22432 27212 22438
rect 26974 22400 27030 22409
rect 27030 22380 27160 22386
rect 27030 22374 27212 22380
rect 27252 22432 27304 22438
rect 27252 22374 27304 22380
rect 27030 22358 27200 22374
rect 26974 22335 27030 22344
rect 26620 22222 26924 22250
rect 26700 22160 26752 22166
rect 26700 22102 26752 22108
rect 26712 21894 26740 22102
rect 26700 21888 26752 21894
rect 26700 21830 26752 21836
rect 26792 21888 26844 21894
rect 26896 21876 26924 22222
rect 27356 22166 27384 23462
rect 27528 23112 27580 23118
rect 27580 23060 27752 23066
rect 27528 23054 27752 23060
rect 27540 23038 27752 23054
rect 27724 22574 27752 23038
rect 27908 22710 27936 24278
rect 28000 23866 28028 24686
rect 28080 24064 28132 24070
rect 28080 24006 28132 24012
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 27988 23588 28040 23594
rect 27988 23530 28040 23536
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27908 22574 27936 22646
rect 27528 22568 27580 22574
rect 27434 22536 27490 22545
rect 27490 22516 27528 22522
rect 27490 22510 27580 22516
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27896 22568 27948 22574
rect 27896 22510 27948 22516
rect 27490 22494 27568 22510
rect 27434 22471 27490 22480
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 27344 22160 27396 22166
rect 27342 22128 27344 22137
rect 27396 22128 27398 22137
rect 27540 22098 27568 22374
rect 27342 22063 27398 22072
rect 27528 22092 27580 22098
rect 27632 22094 27660 22510
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27816 22234 27844 22374
rect 27804 22228 27856 22234
rect 28000 22216 28028 23530
rect 27804 22170 27856 22176
rect 27908 22188 28028 22216
rect 27632 22066 27844 22094
rect 27528 22034 27580 22040
rect 27436 22024 27488 22030
rect 27436 21966 27488 21972
rect 26976 21888 27028 21894
rect 26896 21848 26976 21876
rect 26792 21830 26844 21836
rect 26976 21830 27028 21836
rect 26804 21554 26832 21830
rect 26792 21548 26844 21554
rect 26792 21490 26844 21496
rect 27068 21548 27120 21554
rect 27068 21490 27120 21496
rect 27080 21434 27108 21490
rect 26988 21418 27108 21434
rect 26976 21412 27108 21418
rect 27028 21406 27108 21412
rect 26976 21354 27028 21360
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26792 21344 26844 21350
rect 26792 21286 26844 21292
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 26148 20528 26200 20534
rect 26148 20470 26200 20476
rect 25688 20392 25740 20398
rect 25688 20334 25740 20340
rect 25780 20392 25832 20398
rect 25780 20334 25832 20340
rect 25700 19922 25728 20334
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25688 19780 25740 19786
rect 25688 19722 25740 19728
rect 25504 19440 25556 19446
rect 25332 19366 25452 19394
rect 25504 19382 25556 19388
rect 25424 19310 25452 19366
rect 25412 19304 25464 19310
rect 25412 19246 25464 19252
rect 25136 18896 25188 18902
rect 25136 18838 25188 18844
rect 25596 18896 25648 18902
rect 25596 18838 25648 18844
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24768 18828 24820 18834
rect 24768 18770 24820 18776
rect 25608 18426 25636 18838
rect 25700 18426 25728 19722
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25976 19378 26004 19654
rect 25964 19372 26016 19378
rect 25964 19314 26016 19320
rect 26160 19334 26188 20470
rect 26436 20466 26464 20742
rect 26804 20602 26832 21286
rect 26792 20596 26844 20602
rect 26792 20538 26844 20544
rect 26424 20460 26476 20466
rect 26424 20402 26476 20408
rect 26332 20392 26384 20398
rect 26332 20334 26384 20340
rect 26344 20058 26372 20334
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26332 19916 26384 19922
rect 26332 19858 26384 19864
rect 26344 19514 26372 19858
rect 26332 19508 26384 19514
rect 26332 19450 26384 19456
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25872 19168 25924 19174
rect 25872 19110 25924 19116
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 24492 18216 24544 18222
rect 24492 18158 24544 18164
rect 24952 18216 25004 18222
rect 24952 18158 25004 18164
rect 25320 18216 25372 18222
rect 25320 18158 25372 18164
rect 24308 17808 24360 17814
rect 24308 17750 24360 17756
rect 23572 17672 23624 17678
rect 23572 17614 23624 17620
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 24964 17134 24992 18158
rect 25332 17882 25360 18158
rect 25700 17882 25728 18362
rect 25792 18086 25820 19110
rect 25884 18766 25912 19110
rect 25872 18760 25924 18766
rect 25872 18702 25924 18708
rect 25976 18222 26004 19314
rect 26160 19306 26372 19334
rect 26240 18692 26292 18698
rect 26240 18634 26292 18640
rect 26252 18306 26280 18634
rect 26068 18290 26280 18306
rect 26056 18284 26280 18290
rect 26108 18278 26280 18284
rect 26056 18226 26108 18232
rect 25964 18216 26016 18222
rect 26344 18204 26372 19306
rect 26436 18970 26464 20402
rect 26700 20256 26752 20262
rect 26700 20198 26752 20204
rect 26712 19854 26740 20198
rect 27448 20058 27476 21966
rect 27712 21344 27764 21350
rect 27712 21286 27764 21292
rect 27724 21078 27752 21286
rect 27816 21146 27844 22066
rect 27804 21140 27856 21146
rect 27804 21082 27856 21088
rect 27712 21072 27764 21078
rect 27712 21014 27764 21020
rect 27620 20800 27672 20806
rect 27620 20742 27672 20748
rect 27712 20800 27764 20806
rect 27712 20742 27764 20748
rect 27436 20052 27488 20058
rect 27356 20012 27436 20040
rect 26700 19848 26752 19854
rect 26700 19790 26752 19796
rect 26608 19712 26660 19718
rect 26608 19654 26660 19660
rect 27252 19712 27304 19718
rect 27252 19654 27304 19660
rect 26620 19514 26648 19654
rect 26608 19508 26660 19514
rect 26608 19450 26660 19456
rect 27264 19378 27292 19654
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27356 19174 27384 20012
rect 27436 19994 27488 20000
rect 27528 20052 27580 20058
rect 27528 19994 27580 20000
rect 27436 19304 27488 19310
rect 27436 19246 27488 19252
rect 27344 19168 27396 19174
rect 27344 19110 27396 19116
rect 26424 18964 26476 18970
rect 26424 18906 26476 18912
rect 26516 18964 26568 18970
rect 26516 18906 26568 18912
rect 26528 18426 26556 18906
rect 26792 18896 26844 18902
rect 26792 18838 26844 18844
rect 26882 18864 26938 18873
rect 26516 18420 26568 18426
rect 26516 18362 26568 18368
rect 26804 18290 26832 18838
rect 26882 18799 26938 18808
rect 26896 18680 26924 18799
rect 26976 18692 27028 18698
rect 26896 18652 26976 18680
rect 26896 18290 26924 18652
rect 26976 18634 27028 18640
rect 27448 18426 27476 19246
rect 27540 18698 27568 19994
rect 27632 19922 27660 20742
rect 27724 19990 27752 20742
rect 27712 19984 27764 19990
rect 27712 19926 27764 19932
rect 27620 19916 27672 19922
rect 27620 19858 27672 19864
rect 27816 19718 27844 21082
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27908 19496 27936 22188
rect 28092 22098 28120 24006
rect 28276 23186 28304 24754
rect 29196 24614 29224 25094
rect 29184 24608 29236 24614
rect 29184 24550 29236 24556
rect 29026 24508 29334 24517
rect 29026 24506 29032 24508
rect 29088 24506 29112 24508
rect 29168 24506 29192 24508
rect 29248 24506 29272 24508
rect 29328 24506 29334 24508
rect 29088 24454 29090 24506
rect 29270 24454 29272 24506
rect 29026 24452 29032 24454
rect 29088 24452 29112 24454
rect 29168 24452 29192 24454
rect 29248 24452 29272 24454
rect 29328 24452 29334 24454
rect 29026 24443 29334 24452
rect 29460 24132 29512 24138
rect 29460 24074 29512 24080
rect 28366 23964 28674 23973
rect 28366 23962 28372 23964
rect 28428 23962 28452 23964
rect 28508 23962 28532 23964
rect 28588 23962 28612 23964
rect 28668 23962 28674 23964
rect 28428 23910 28430 23962
rect 28610 23910 28612 23962
rect 28366 23908 28372 23910
rect 28428 23908 28452 23910
rect 28508 23908 28532 23910
rect 28588 23908 28612 23910
rect 28668 23908 28674 23910
rect 28366 23899 28674 23908
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28264 23180 28316 23186
rect 28264 23122 28316 23128
rect 28724 22976 28776 22982
rect 28724 22918 28776 22924
rect 28366 22876 28674 22885
rect 28366 22874 28372 22876
rect 28428 22874 28452 22876
rect 28508 22874 28532 22876
rect 28588 22874 28612 22876
rect 28668 22874 28674 22876
rect 28428 22822 28430 22874
rect 28610 22822 28612 22874
rect 28366 22820 28372 22822
rect 28428 22820 28452 22822
rect 28508 22820 28532 22822
rect 28588 22820 28612 22822
rect 28668 22820 28674 22822
rect 28366 22811 28674 22820
rect 27988 22092 28040 22098
rect 27988 22034 28040 22040
rect 28080 22092 28132 22098
rect 28080 22034 28132 22040
rect 28000 21690 28028 22034
rect 28366 21788 28674 21797
rect 28366 21786 28372 21788
rect 28428 21786 28452 21788
rect 28508 21786 28532 21788
rect 28588 21786 28612 21788
rect 28668 21786 28674 21788
rect 28428 21734 28430 21786
rect 28610 21734 28612 21786
rect 28366 21732 28372 21734
rect 28428 21732 28452 21734
rect 28508 21732 28532 21734
rect 28588 21732 28612 21734
rect 28668 21732 28674 21734
rect 28366 21723 28674 21732
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 28736 21350 28764 22918
rect 28828 22710 28856 23598
rect 29368 23520 29420 23526
rect 29368 23462 29420 23468
rect 29026 23420 29334 23429
rect 29026 23418 29032 23420
rect 29088 23418 29112 23420
rect 29168 23418 29192 23420
rect 29248 23418 29272 23420
rect 29328 23418 29334 23420
rect 29088 23366 29090 23418
rect 29270 23366 29272 23418
rect 29026 23364 29032 23366
rect 29088 23364 29112 23366
rect 29168 23364 29192 23366
rect 29248 23364 29272 23366
rect 29328 23364 29334 23366
rect 29026 23355 29334 23364
rect 28908 23112 28960 23118
rect 28908 23054 28960 23060
rect 28920 22778 28948 23054
rect 29380 22778 29408 23462
rect 28908 22772 28960 22778
rect 28908 22714 28960 22720
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 28816 22704 28868 22710
rect 28816 22646 28868 22652
rect 29472 22574 29500 24074
rect 29656 23798 29684 28086
rect 29736 27532 29788 27538
rect 29736 27474 29788 27480
rect 29748 25362 29776 27474
rect 29840 27130 29868 30738
rect 30392 30394 30420 30738
rect 30380 30388 30432 30394
rect 30380 30330 30432 30336
rect 29920 30184 29972 30190
rect 29920 30126 29972 30132
rect 30012 30184 30064 30190
rect 30012 30126 30064 30132
rect 30656 30184 30708 30190
rect 30656 30126 30708 30132
rect 30932 30184 30984 30190
rect 30932 30126 30984 30132
rect 29932 29850 29960 30126
rect 29920 29844 29972 29850
rect 29920 29786 29972 29792
rect 30024 28966 30052 30126
rect 30196 29844 30248 29850
rect 30196 29786 30248 29792
rect 30012 28960 30064 28966
rect 30012 28902 30064 28908
rect 30208 28608 30236 29786
rect 30380 29708 30432 29714
rect 30380 29650 30432 29656
rect 30392 28665 30420 29650
rect 30668 29306 30696 30126
rect 30656 29300 30708 29306
rect 30656 29242 30708 29248
rect 30944 29102 30972 30126
rect 30932 29096 30984 29102
rect 30932 29038 30984 29044
rect 30840 28960 30892 28966
rect 30840 28902 30892 28908
rect 30852 28694 30880 28902
rect 30840 28688 30892 28694
rect 29932 28580 30236 28608
rect 30378 28656 30434 28665
rect 30840 28630 30892 28636
rect 30378 28591 30434 28600
rect 29932 28150 29960 28580
rect 30196 28416 30248 28422
rect 30196 28358 30248 28364
rect 30208 28218 30236 28358
rect 30196 28212 30248 28218
rect 30196 28154 30248 28160
rect 30380 28212 30432 28218
rect 30380 28154 30432 28160
rect 29920 28144 29972 28150
rect 29920 28086 29972 28092
rect 30194 28112 30250 28121
rect 29932 27878 29960 28086
rect 30194 28047 30196 28056
rect 30248 28047 30250 28056
rect 30196 28018 30248 28024
rect 30104 28008 30156 28014
rect 30104 27950 30156 27956
rect 29920 27872 29972 27878
rect 29920 27814 29972 27820
rect 30116 27441 30144 27950
rect 30392 27674 30420 28154
rect 30746 27976 30802 27985
rect 30802 27934 30880 27962
rect 30746 27911 30802 27920
rect 30852 27878 30880 27934
rect 30748 27872 30800 27878
rect 30748 27814 30800 27820
rect 30840 27872 30892 27878
rect 30840 27814 30892 27820
rect 30760 27674 30788 27814
rect 30380 27668 30432 27674
rect 30380 27610 30432 27616
rect 30748 27668 30800 27674
rect 30748 27610 30800 27616
rect 30392 27470 30420 27610
rect 30564 27600 30616 27606
rect 30564 27542 30616 27548
rect 30380 27464 30432 27470
rect 30102 27432 30158 27441
rect 30380 27406 30432 27412
rect 30102 27367 30158 27376
rect 30472 27328 30524 27334
rect 30472 27270 30524 27276
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 30484 27062 30512 27270
rect 30472 27056 30524 27062
rect 30472 26998 30524 27004
rect 30576 26926 30604 27542
rect 30852 27538 30880 27814
rect 30840 27532 30892 27538
rect 30840 27474 30892 27480
rect 30656 27464 30708 27470
rect 30656 27406 30708 27412
rect 30564 26920 30616 26926
rect 30564 26862 30616 26868
rect 30104 26852 30156 26858
rect 30104 26794 30156 26800
rect 30116 25770 30144 26794
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30288 26308 30340 26314
rect 30288 26250 30340 26256
rect 30104 25764 30156 25770
rect 30104 25706 30156 25712
rect 29736 25356 29788 25362
rect 29736 25298 29788 25304
rect 29748 24954 29776 25298
rect 29736 24948 29788 24954
rect 29736 24890 29788 24896
rect 30300 24750 30328 26250
rect 30392 25838 30420 26726
rect 30668 26586 30696 27406
rect 30852 27130 30880 27474
rect 30944 27470 30972 29038
rect 30932 27464 30984 27470
rect 30932 27406 30984 27412
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30656 26580 30708 26586
rect 30656 26522 30708 26528
rect 30944 26450 30972 27406
rect 30932 26444 30984 26450
rect 30932 26386 30984 26392
rect 30380 25832 30432 25838
rect 30380 25774 30432 25780
rect 30392 25158 30420 25774
rect 30748 25492 30800 25498
rect 30748 25434 30800 25440
rect 30380 25152 30432 25158
rect 30380 25094 30432 25100
rect 30288 24744 30340 24750
rect 30288 24686 30340 24692
rect 30380 24200 30432 24206
rect 30380 24142 30432 24148
rect 29644 23792 29696 23798
rect 29644 23734 29696 23740
rect 30392 23322 30420 24142
rect 30380 23316 30432 23322
rect 30380 23258 30432 23264
rect 29920 23248 29972 23254
rect 29920 23190 29972 23196
rect 29932 22778 29960 23190
rect 30288 23112 30340 23118
rect 30288 23054 30340 23060
rect 29920 22772 29972 22778
rect 29920 22714 29972 22720
rect 30300 22642 30328 23054
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 29460 22568 29512 22574
rect 29460 22510 29512 22516
rect 29736 22500 29788 22506
rect 29736 22442 29788 22448
rect 29026 22332 29334 22341
rect 29026 22330 29032 22332
rect 29088 22330 29112 22332
rect 29168 22330 29192 22332
rect 29248 22330 29272 22332
rect 29328 22330 29334 22332
rect 29088 22278 29090 22330
rect 29270 22278 29272 22330
rect 29026 22276 29032 22278
rect 29088 22276 29112 22278
rect 29168 22276 29192 22278
rect 29248 22276 29272 22278
rect 29328 22276 29334 22278
rect 29026 22267 29334 22276
rect 29748 22094 29776 22442
rect 30300 22094 30328 22578
rect 29748 22066 29960 22094
rect 28172 21344 28224 21350
rect 28172 21286 28224 21292
rect 28724 21344 28776 21350
rect 28724 21286 28776 21292
rect 28184 21146 28212 21286
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28366 20700 28674 20709
rect 28366 20698 28372 20700
rect 28428 20698 28452 20700
rect 28508 20698 28532 20700
rect 28588 20698 28612 20700
rect 28668 20698 28674 20700
rect 28428 20646 28430 20698
rect 28610 20646 28612 20698
rect 28366 20644 28372 20646
rect 28428 20644 28452 20646
rect 28508 20644 28532 20646
rect 28588 20644 28612 20646
rect 28668 20644 28674 20646
rect 28366 20635 28674 20644
rect 27988 20596 28040 20602
rect 27988 20538 28040 20544
rect 28000 19922 28028 20538
rect 28078 20496 28134 20505
rect 28134 20454 28212 20482
rect 28078 20431 28134 20440
rect 28184 20398 28212 20454
rect 28172 20392 28224 20398
rect 28224 20352 28304 20380
rect 28172 20334 28224 20340
rect 28080 20324 28132 20330
rect 28080 20266 28132 20272
rect 27988 19916 28040 19922
rect 27988 19858 28040 19864
rect 27724 19468 27936 19496
rect 27724 19242 27752 19468
rect 27908 19378 27936 19468
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 27896 19372 27948 19378
rect 27896 19314 27948 19320
rect 27712 19236 27764 19242
rect 27712 19178 27764 19184
rect 27816 18970 27844 19314
rect 28000 19174 28028 19858
rect 28092 19514 28120 20266
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28184 20058 28212 20198
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28276 19990 28304 20352
rect 28264 19984 28316 19990
rect 28264 19926 28316 19932
rect 28736 19786 28764 21286
rect 29026 21244 29334 21253
rect 29026 21242 29032 21244
rect 29088 21242 29112 21244
rect 29168 21242 29192 21244
rect 29248 21242 29272 21244
rect 29328 21242 29334 21244
rect 29088 21190 29090 21242
rect 29270 21190 29272 21242
rect 29026 21188 29032 21190
rect 29088 21188 29112 21190
rect 29168 21188 29192 21190
rect 29248 21188 29272 21190
rect 29328 21188 29334 21190
rect 29026 21179 29334 21188
rect 29734 21040 29790 21049
rect 29790 20998 29868 21026
rect 29734 20975 29790 20984
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 29026 20156 29334 20165
rect 29026 20154 29032 20156
rect 29088 20154 29112 20156
rect 29168 20154 29192 20156
rect 29248 20154 29272 20156
rect 29328 20154 29334 20156
rect 29088 20102 29090 20154
rect 29270 20102 29272 20154
rect 29026 20100 29032 20102
rect 29088 20100 29112 20102
rect 29168 20100 29192 20102
rect 29248 20100 29272 20102
rect 29328 20100 29334 20102
rect 29026 20091 29334 20100
rect 28908 19984 28960 19990
rect 28908 19926 28960 19932
rect 28724 19780 28776 19786
rect 28724 19722 28776 19728
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28276 19378 28304 19654
rect 28366 19612 28674 19621
rect 28366 19610 28372 19612
rect 28428 19610 28452 19612
rect 28508 19610 28532 19612
rect 28588 19610 28612 19612
rect 28668 19610 28674 19612
rect 28428 19558 28430 19610
rect 28610 19558 28612 19610
rect 28366 19556 28372 19558
rect 28428 19556 28452 19558
rect 28508 19556 28532 19558
rect 28588 19556 28612 19558
rect 28668 19556 28674 19558
rect 28366 19547 28674 19556
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28736 19310 28764 19722
rect 28920 19514 28948 19926
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 29012 19394 29040 19790
rect 28920 19366 29040 19394
rect 28724 19304 28776 19310
rect 28724 19246 28776 19252
rect 27988 19168 28040 19174
rect 27988 19110 28040 19116
rect 28356 19168 28408 19174
rect 28356 19110 28408 19116
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 28368 18834 28396 19110
rect 28920 18834 28948 19366
rect 29380 19174 29408 20402
rect 29460 20324 29512 20330
rect 29460 20266 29512 20272
rect 29472 19718 29500 20266
rect 29564 20058 29592 20878
rect 29656 20602 29684 20878
rect 29840 20602 29868 20998
rect 29644 20596 29696 20602
rect 29644 20538 29696 20544
rect 29828 20596 29880 20602
rect 29828 20538 29880 20544
rect 29840 20058 29868 20538
rect 29552 20052 29604 20058
rect 29552 19994 29604 20000
rect 29828 20052 29880 20058
rect 29828 19994 29880 20000
rect 29932 19990 29960 22066
rect 30208 22066 30328 22094
rect 30208 21554 30236 22066
rect 30196 21548 30248 21554
rect 30196 21490 30248 21496
rect 30012 20800 30064 20806
rect 30012 20742 30064 20748
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30024 20330 30052 20742
rect 30012 20324 30064 20330
rect 30012 20266 30064 20272
rect 30116 20262 30144 20742
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 29920 19984 29972 19990
rect 29920 19926 29972 19932
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 29552 19236 29604 19242
rect 29552 19178 29604 19184
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29026 19068 29334 19077
rect 29026 19066 29032 19068
rect 29088 19066 29112 19068
rect 29168 19066 29192 19068
rect 29248 19066 29272 19068
rect 29328 19066 29334 19068
rect 29088 19014 29090 19066
rect 29270 19014 29272 19066
rect 29026 19012 29032 19014
rect 29088 19012 29112 19014
rect 29168 19012 29192 19014
rect 29248 19012 29272 19014
rect 29328 19012 29334 19014
rect 29026 19003 29334 19012
rect 28356 18828 28408 18834
rect 28356 18770 28408 18776
rect 28908 18828 28960 18834
rect 28908 18770 28960 18776
rect 28814 18728 28870 18737
rect 27528 18692 27580 18698
rect 28814 18663 28870 18672
rect 28908 18692 28960 18698
rect 27528 18634 27580 18640
rect 27436 18420 27488 18426
rect 27436 18362 27488 18368
rect 26792 18284 26844 18290
rect 26792 18226 26844 18232
rect 26884 18284 26936 18290
rect 26884 18226 26936 18232
rect 26424 18216 26476 18222
rect 26344 18176 26424 18204
rect 25964 18158 26016 18164
rect 26424 18158 26476 18164
rect 25780 18080 25832 18086
rect 25780 18022 25832 18028
rect 25320 17876 25372 17882
rect 25320 17818 25372 17824
rect 25688 17876 25740 17882
rect 25688 17818 25740 17824
rect 25044 17808 25096 17814
rect 25044 17750 25096 17756
rect 25056 17338 25084 17750
rect 25688 17740 25740 17746
rect 25688 17682 25740 17688
rect 25412 17672 25464 17678
rect 25412 17614 25464 17620
rect 25044 17332 25096 17338
rect 25044 17274 25096 17280
rect 23112 17128 23164 17134
rect 23112 17070 23164 17076
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 23664 17060 23716 17066
rect 23664 17002 23716 17008
rect 21272 16788 21324 16794
rect 21272 16730 21324 16736
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 21006 16348 21314 16357
rect 21006 16346 21012 16348
rect 21068 16346 21092 16348
rect 21148 16346 21172 16348
rect 21228 16346 21252 16348
rect 21308 16346 21314 16348
rect 21068 16294 21070 16346
rect 21250 16294 21252 16346
rect 21006 16292 21012 16294
rect 21068 16292 21092 16294
rect 21148 16292 21172 16294
rect 21228 16292 21252 16294
rect 21308 16292 21314 16294
rect 21006 16283 21314 16292
rect 23112 16176 23164 16182
rect 23112 16118 23164 16124
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14482 20668 14894
rect 20916 14550 20944 16050
rect 21666 15804 21974 15813
rect 21666 15802 21672 15804
rect 21728 15802 21752 15804
rect 21808 15802 21832 15804
rect 21888 15802 21912 15804
rect 21968 15802 21974 15804
rect 21728 15750 21730 15802
rect 21910 15750 21912 15802
rect 21666 15748 21672 15750
rect 21728 15748 21752 15750
rect 21808 15748 21832 15750
rect 21888 15748 21912 15750
rect 21968 15748 21974 15750
rect 21666 15739 21974 15748
rect 23124 15706 23152 16118
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 21548 15632 21600 15638
rect 21548 15574 21600 15580
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21006 15260 21314 15269
rect 21006 15258 21012 15260
rect 21068 15258 21092 15260
rect 21148 15258 21172 15260
rect 21228 15258 21252 15260
rect 21308 15258 21314 15260
rect 21068 15206 21070 15258
rect 21250 15206 21252 15258
rect 21006 15204 21012 15206
rect 21068 15204 21092 15206
rect 21148 15204 21172 15206
rect 21228 15204 21252 15206
rect 21308 15204 21314 15206
rect 21006 15195 21314 15204
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14550 21036 14758
rect 20904 14544 20956 14550
rect 20904 14486 20956 14492
rect 20996 14544 21048 14550
rect 20996 14486 21048 14492
rect 20628 14476 20680 14482
rect 20628 14418 20680 14424
rect 20640 12442 20668 14418
rect 21376 14414 21404 15302
rect 21560 14822 21588 15574
rect 23124 15570 23152 15642
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 23112 15564 23164 15570
rect 23112 15506 23164 15512
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22192 15020 22244 15026
rect 22192 14962 22244 14968
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 20824 14074 20852 14350
rect 20904 14340 20956 14346
rect 20904 14282 20956 14288
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20916 13938 20944 14282
rect 21006 14172 21314 14181
rect 21006 14170 21012 14172
rect 21068 14170 21092 14172
rect 21148 14170 21172 14172
rect 21228 14170 21252 14172
rect 21308 14170 21314 14172
rect 21068 14118 21070 14170
rect 21250 14118 21252 14170
rect 21006 14116 21012 14118
rect 21068 14116 21092 14118
rect 21148 14116 21172 14118
rect 21228 14116 21252 14118
rect 21308 14116 21314 14118
rect 21006 14107 21314 14116
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20824 12986 20852 13806
rect 20904 13728 20956 13734
rect 20904 13670 20956 13676
rect 20916 13530 20944 13670
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21376 13326 21404 14350
rect 21468 13462 21496 14758
rect 21666 14716 21974 14725
rect 21666 14714 21672 14716
rect 21728 14714 21752 14716
rect 21808 14714 21832 14716
rect 21888 14714 21912 14716
rect 21968 14714 21974 14716
rect 21728 14662 21730 14714
rect 21910 14662 21912 14714
rect 21666 14660 21672 14662
rect 21728 14660 21752 14662
rect 21808 14660 21832 14662
rect 21888 14660 21912 14662
rect 21968 14660 21974 14662
rect 21666 14651 21974 14660
rect 21548 13728 21600 13734
rect 21548 13670 21600 13676
rect 21456 13456 21508 13462
rect 21456 13398 21508 13404
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21006 13084 21314 13093
rect 21006 13082 21012 13084
rect 21068 13082 21092 13084
rect 21148 13082 21172 13084
rect 21228 13082 21252 13084
rect 21308 13082 21314 13084
rect 21068 13030 21070 13082
rect 21250 13030 21252 13082
rect 21006 13028 21012 13030
rect 21068 13028 21092 13030
rect 21148 13028 21172 13030
rect 21228 13028 21252 13030
rect 21308 13028 21314 13030
rect 21006 13019 21314 13028
rect 20812 12980 20864 12986
rect 20812 12922 20864 12928
rect 21376 12918 21404 13262
rect 21560 12986 21588 13670
rect 21666 13628 21974 13637
rect 21666 13626 21672 13628
rect 21728 13626 21752 13628
rect 21808 13626 21832 13628
rect 21888 13626 21912 13628
rect 21968 13626 21974 13628
rect 21728 13574 21730 13626
rect 21910 13574 21912 13626
rect 21666 13572 21672 13574
rect 21728 13572 21752 13574
rect 21808 13572 21832 13574
rect 21888 13572 21912 13574
rect 21968 13572 21974 13574
rect 21666 13563 21974 13572
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 21836 12986 21864 13262
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21364 12912 21416 12918
rect 21364 12854 21416 12860
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20456 12294 20668 12322
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19708 11892 19760 11898
rect 19708 11834 19760 11840
rect 19432 11824 19484 11830
rect 19432 11766 19484 11772
rect 19996 11286 20024 12038
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 20536 11688 20588 11694
rect 20536 11630 20588 11636
rect 19984 11280 20036 11286
rect 19984 11222 20036 11228
rect 20180 11218 20208 11630
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10674 19288 11086
rect 20272 10810 20300 11154
rect 20260 10804 20312 10810
rect 20260 10746 20312 10752
rect 19340 10736 19392 10742
rect 19340 10678 19392 10684
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19248 10464 19300 10470
rect 19248 10406 19300 10412
rect 19260 10062 19288 10406
rect 19352 10266 19380 10678
rect 19340 10260 19392 10266
rect 19340 10202 19392 10208
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 20258 9616 20314 9625
rect 20258 9551 20260 9560
rect 20312 9551 20314 9560
rect 20260 9522 20312 9528
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18616 9178 18644 9386
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 18984 9110 19012 9318
rect 19628 9110 19656 9318
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 19616 9104 19668 9110
rect 19616 9046 19668 9052
rect 18512 9036 18564 9042
rect 18512 8978 18564 8984
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18236 8356 18288 8362
rect 18236 8298 18288 8304
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 18248 7546 18276 8298
rect 18340 7954 18368 8570
rect 18432 8022 18460 8774
rect 18420 8016 18472 8022
rect 18420 7958 18472 7964
rect 18328 7948 18380 7954
rect 18328 7890 18380 7896
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18524 7342 18552 8978
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18696 8832 18748 8838
rect 18696 8774 18748 8780
rect 18708 8634 18736 8774
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18800 8430 18828 8910
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18892 8498 18920 8842
rect 18984 8566 19012 9046
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19260 8634 19288 8910
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18236 7268 18288 7274
rect 18236 7210 18288 7216
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17684 6384 17736 6390
rect 17684 6326 17736 6332
rect 17696 5914 17724 6326
rect 17972 6254 18000 6666
rect 18248 6390 18276 7210
rect 18602 6896 18658 6905
rect 18420 6860 18472 6866
rect 18602 6831 18658 6840
rect 18420 6802 18472 6808
rect 18432 6458 18460 6802
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 17960 6248 18012 6254
rect 17960 6190 18012 6196
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17960 5364 18012 5370
rect 17960 5306 18012 5312
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17000 3896 17080 3924
rect 16948 3878 17000 3884
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 17052 3602 17080 3896
rect 17604 3738 17632 4150
rect 17972 4078 18000 5306
rect 18064 5273 18092 5306
rect 18050 5264 18106 5273
rect 18050 5199 18106 5208
rect 18064 5166 18092 5199
rect 18052 5160 18104 5166
rect 18052 5102 18104 5108
rect 18144 5160 18196 5166
rect 18144 5102 18196 5108
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18064 4282 18092 4626
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17880 3738 17908 3946
rect 18064 3890 18092 4218
rect 17972 3862 18092 3890
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17040 3596 17092 3602
rect 17040 3538 17092 3544
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 15384 2984 15436 2990
rect 15384 2926 15436 2932
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16960 2774 16988 3470
rect 17972 2990 18000 3862
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 16776 2746 16988 2774
rect 16776 800 16804 2746
rect 18064 800 18092 2994
rect 18156 2922 18184 5102
rect 18248 4690 18276 6326
rect 18616 5914 18644 6831
rect 18800 6254 18828 8366
rect 19708 8356 19760 8362
rect 19708 8298 19760 8304
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19260 8090 19288 8230
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19340 7880 19392 7886
rect 19340 7822 19392 7828
rect 19352 7002 19380 7822
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19076 6458 19104 6598
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18788 6248 18840 6254
rect 18788 6190 18840 6196
rect 18604 5908 18656 5914
rect 18604 5850 18656 5856
rect 18696 5840 18748 5846
rect 18696 5782 18748 5788
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18248 3058 18276 4014
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18340 2922 18368 5102
rect 18432 4758 18460 5510
rect 18512 5228 18564 5234
rect 18564 5188 18644 5216
rect 18512 5170 18564 5176
rect 18616 5137 18644 5188
rect 18602 5128 18658 5137
rect 18602 5063 18658 5072
rect 18420 4752 18472 4758
rect 18420 4694 18472 4700
rect 18432 4214 18460 4694
rect 18708 4690 18736 5782
rect 18800 5710 18828 6190
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18788 5704 18840 5710
rect 18788 5646 18840 5652
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18708 4078 18736 4626
rect 18800 4146 18828 5646
rect 19076 5234 19104 5850
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19536 5370 19564 5646
rect 19524 5364 19576 5370
rect 19524 5306 19576 5312
rect 19246 5264 19302 5273
rect 19064 5228 19116 5234
rect 19246 5199 19248 5208
rect 19064 5170 19116 5176
rect 19300 5199 19302 5208
rect 19248 5170 19300 5176
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 18892 4282 18920 5102
rect 18984 4950 19288 4978
rect 18984 4758 19012 4950
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18788 4140 18840 4146
rect 18788 4082 18840 4088
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 18328 2916 18380 2922
rect 18328 2858 18380 2864
rect 18708 2854 18736 4014
rect 19076 3058 19104 4762
rect 19260 4554 19288 4950
rect 19432 4616 19484 4622
rect 19432 4558 19484 4564
rect 19248 4548 19300 4554
rect 19248 4490 19300 4496
rect 19444 3738 19472 4558
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19536 4010 19564 4422
rect 19628 4282 19656 4422
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19524 4004 19576 4010
rect 19524 3946 19576 3952
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19432 3052 19484 3058
rect 19432 2994 19484 3000
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 19444 1442 19472 2994
rect 19720 2854 19748 8298
rect 20180 7954 20208 9318
rect 20364 8430 20392 9454
rect 20352 8424 20404 8430
rect 20352 8366 20404 8372
rect 20364 7954 20392 8366
rect 20444 8288 20496 8294
rect 20444 8230 20496 8236
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20352 7948 20404 7954
rect 20352 7890 20404 7896
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20088 6934 20116 7822
rect 20456 7206 20484 8230
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20456 6798 20484 7142
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20260 6724 20312 6730
rect 20260 6666 20312 6672
rect 20272 6118 20300 6666
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20076 5296 20128 5302
rect 20076 5238 20128 5244
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 19812 3670 19840 4694
rect 20088 4282 20116 5238
rect 20548 4978 20576 11630
rect 20640 8922 20668 12294
rect 21006 11996 21314 12005
rect 21006 11994 21012 11996
rect 21068 11994 21092 11996
rect 21148 11994 21172 11996
rect 21228 11994 21252 11996
rect 21308 11994 21314 11996
rect 21068 11942 21070 11994
rect 21250 11942 21252 11994
rect 21006 11940 21012 11942
rect 21068 11940 21092 11942
rect 21148 11940 21172 11942
rect 21228 11940 21252 11942
rect 21308 11940 21314 11942
rect 21006 11931 21314 11940
rect 21376 11762 21404 12854
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21468 12374 21496 12786
rect 21456 12368 21508 12374
rect 21456 12310 21508 12316
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 20720 11688 20772 11694
rect 20720 11630 20772 11636
rect 20732 10810 20760 11630
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20732 10538 20760 10746
rect 20720 10532 20772 10538
rect 20720 10474 20772 10480
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20732 9110 20760 9862
rect 20824 9518 20852 11086
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21006 10908 21314 10917
rect 21006 10906 21012 10908
rect 21068 10906 21092 10908
rect 21148 10906 21172 10908
rect 21228 10906 21252 10908
rect 21308 10906 21314 10908
rect 21068 10854 21070 10906
rect 21250 10854 21252 10906
rect 21006 10852 21012 10854
rect 21068 10852 21092 10854
rect 21148 10852 21172 10854
rect 21228 10852 21252 10854
rect 21308 10852 21314 10854
rect 21006 10843 21314 10852
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20916 9586 20944 10746
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21008 10198 21036 10406
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 21006 9820 21314 9829
rect 21006 9818 21012 9820
rect 21068 9818 21092 9820
rect 21148 9818 21172 9820
rect 21228 9818 21252 9820
rect 21308 9818 21314 9820
rect 21068 9766 21070 9818
rect 21250 9766 21252 9818
rect 21006 9764 21012 9766
rect 21068 9764 21092 9766
rect 21148 9764 21172 9766
rect 21228 9764 21252 9766
rect 21308 9764 21314 9766
rect 21006 9755 21314 9764
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20812 9512 20864 9518
rect 20812 9454 20864 9460
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 20640 8894 20852 8922
rect 20628 6860 20680 6866
rect 20628 6802 20680 6808
rect 20640 5914 20668 6802
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20732 6458 20760 6734
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20640 5166 20668 5850
rect 20628 5160 20680 5166
rect 20720 5160 20772 5166
rect 20628 5102 20680 5108
rect 20718 5128 20720 5137
rect 20772 5128 20774 5137
rect 20718 5063 20774 5072
rect 20548 4950 20668 4978
rect 20352 4616 20404 4622
rect 20352 4558 20404 4564
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 20272 4146 20300 4422
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 19800 3664 19852 3670
rect 19800 3606 19852 3612
rect 20272 3534 20300 4082
rect 20364 4010 20392 4558
rect 20444 4480 20496 4486
rect 20444 4422 20496 4428
rect 20352 4004 20404 4010
rect 20352 3946 20404 3952
rect 20456 3738 20484 4422
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20640 3398 20668 4950
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20732 3466 20760 4626
rect 20824 3482 20852 8894
rect 21192 8838 21220 9318
rect 21284 9110 21312 9454
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21006 8732 21314 8741
rect 21006 8730 21012 8732
rect 21068 8730 21092 8732
rect 21148 8730 21172 8732
rect 21228 8730 21252 8732
rect 21308 8730 21314 8732
rect 21068 8678 21070 8730
rect 21250 8678 21252 8730
rect 21006 8676 21012 8678
rect 21068 8676 21092 8678
rect 21148 8676 21172 8678
rect 21228 8676 21252 8678
rect 21308 8676 21314 8678
rect 21006 8667 21314 8676
rect 21376 8634 21404 11018
rect 21456 10532 21508 10538
rect 21456 10474 21508 10480
rect 21468 9926 21496 10474
rect 21456 9920 21508 9926
rect 21456 9862 21508 9868
rect 21468 9042 21496 9862
rect 21456 9036 21508 9042
rect 21456 8978 21508 8984
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 20904 8356 20956 8362
rect 20904 8298 20956 8304
rect 20916 7750 20944 8298
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 21006 7644 21314 7653
rect 21006 7642 21012 7644
rect 21068 7642 21092 7644
rect 21148 7642 21172 7644
rect 21228 7642 21252 7644
rect 21308 7642 21314 7644
rect 21068 7590 21070 7642
rect 21250 7590 21252 7642
rect 21006 7588 21012 7590
rect 21068 7588 21092 7590
rect 21148 7588 21172 7590
rect 21228 7588 21252 7590
rect 21308 7588 21314 7590
rect 21006 7579 21314 7588
rect 21468 7410 21496 8978
rect 21560 8362 21588 12922
rect 22020 12850 22048 14758
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 22112 13530 22140 13806
rect 22100 13524 22152 13530
rect 22100 13466 22152 13472
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21666 12540 21974 12549
rect 21666 12538 21672 12540
rect 21728 12538 21752 12540
rect 21808 12538 21832 12540
rect 21888 12538 21912 12540
rect 21968 12538 21974 12540
rect 21728 12486 21730 12538
rect 21910 12486 21912 12538
rect 21666 12484 21672 12486
rect 21728 12484 21752 12486
rect 21808 12484 21832 12486
rect 21888 12484 21912 12486
rect 21968 12484 21974 12486
rect 21666 12475 21974 12484
rect 22100 12368 22152 12374
rect 22204 12356 22232 14962
rect 22480 14958 22508 15302
rect 22560 15156 22612 15162
rect 22560 15098 22612 15104
rect 22572 14958 22600 15098
rect 22940 15026 23244 15042
rect 22928 15020 23244 15026
rect 22980 15014 23244 15020
rect 22928 14962 22980 14968
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22296 12374 22324 13874
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22388 12442 22416 12718
rect 22376 12436 22428 12442
rect 22376 12378 22428 12384
rect 22152 12328 22232 12356
rect 22284 12368 22336 12374
rect 22100 12310 22152 12316
rect 22284 12310 22336 12316
rect 21666 11452 21974 11461
rect 21666 11450 21672 11452
rect 21728 11450 21752 11452
rect 21808 11450 21832 11452
rect 21888 11450 21912 11452
rect 21968 11450 21974 11452
rect 21728 11398 21730 11450
rect 21910 11398 21912 11450
rect 21666 11396 21672 11398
rect 21728 11396 21752 11398
rect 21808 11396 21832 11398
rect 21888 11396 21912 11398
rect 21968 11396 21974 11398
rect 21666 11387 21974 11396
rect 22572 11354 22600 14894
rect 23216 14822 23244 15014
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23204 14816 23256 14822
rect 23204 14758 23256 14764
rect 22848 14464 22876 14758
rect 23032 14618 23060 14758
rect 23584 14618 23612 15574
rect 23020 14612 23072 14618
rect 23020 14554 23072 14560
rect 23572 14612 23624 14618
rect 23572 14554 23624 14560
rect 23676 14482 23704 17002
rect 25424 16998 25452 17614
rect 25412 16992 25464 16998
rect 25412 16934 25464 16940
rect 25504 16992 25556 16998
rect 25504 16934 25556 16940
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24136 15706 24164 15982
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24584 15904 24636 15910
rect 24584 15846 24636 15852
rect 24412 15706 24440 15846
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 24400 15700 24452 15706
rect 24400 15642 24452 15648
rect 24596 15570 24624 15846
rect 24584 15564 24636 15570
rect 24584 15506 24636 15512
rect 24596 15366 24624 15506
rect 24584 15360 24636 15366
rect 24584 15302 24636 15308
rect 24308 14952 24360 14958
rect 24308 14894 24360 14900
rect 22928 14476 22980 14482
rect 22756 14436 22928 14464
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22664 13938 22692 14214
rect 22652 13932 22704 13938
rect 22652 13874 22704 13880
rect 22652 13456 22704 13462
rect 22652 13398 22704 13404
rect 22664 12442 22692 13398
rect 22756 12442 22784 14436
rect 22928 14418 22980 14424
rect 23664 14476 23716 14482
rect 23664 14418 23716 14424
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 22836 12708 22888 12714
rect 22836 12650 22888 12656
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22744 12436 22796 12442
rect 22848 12434 22876 12650
rect 22928 12436 22980 12442
rect 22848 12406 22928 12434
rect 22744 12378 22796 12384
rect 22928 12378 22980 12384
rect 23400 12306 23428 13670
rect 23492 13394 23520 13806
rect 24044 13530 24072 14418
rect 24320 14346 24348 14894
rect 24768 14816 24820 14822
rect 24768 14758 24820 14764
rect 24308 14340 24360 14346
rect 24308 14282 24360 14288
rect 24780 14278 24808 14758
rect 25424 14414 25452 16934
rect 25516 16114 25544 16934
rect 25504 16108 25556 16114
rect 25504 16050 25556 16056
rect 25412 14408 25464 14414
rect 25412 14350 25464 14356
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24124 13796 24176 13802
rect 24124 13738 24176 13744
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24136 13462 24164 13738
rect 24780 13530 24808 14214
rect 24860 13796 24912 13802
rect 24860 13738 24912 13744
rect 24872 13530 24900 13738
rect 24768 13524 24820 13530
rect 24768 13466 24820 13472
rect 24860 13524 24912 13530
rect 24860 13466 24912 13472
rect 24124 13456 24176 13462
rect 24124 13398 24176 13404
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23492 12374 23520 13330
rect 23940 12776 23992 12782
rect 23940 12718 23992 12724
rect 23952 12442 23980 12718
rect 24136 12442 24164 13398
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 25608 12986 25636 13330
rect 25596 12980 25648 12986
rect 25596 12922 25648 12928
rect 25700 12442 25728 17682
rect 26804 17678 26832 18226
rect 26896 17746 26924 18226
rect 27540 18222 27568 18634
rect 27896 18624 27948 18630
rect 27896 18566 27948 18572
rect 28724 18624 28776 18630
rect 28724 18566 28776 18572
rect 27528 18216 27580 18222
rect 27528 18158 27580 18164
rect 27908 17814 27936 18566
rect 28366 18524 28674 18533
rect 28366 18522 28372 18524
rect 28428 18522 28452 18524
rect 28508 18522 28532 18524
rect 28588 18522 28612 18524
rect 28668 18522 28674 18524
rect 28428 18470 28430 18522
rect 28610 18470 28612 18522
rect 28366 18468 28372 18470
rect 28428 18468 28452 18470
rect 28508 18468 28532 18470
rect 28588 18468 28612 18470
rect 28668 18468 28674 18470
rect 28366 18459 28674 18468
rect 28080 18080 28132 18086
rect 28080 18022 28132 18028
rect 28092 17814 28120 18022
rect 28736 17882 28764 18566
rect 28828 17882 28856 18663
rect 28908 18634 28960 18640
rect 28724 17876 28776 17882
rect 28724 17818 28776 17824
rect 28816 17876 28868 17882
rect 28816 17818 28868 17824
rect 28920 17814 28948 18634
rect 29026 17980 29334 17989
rect 29026 17978 29032 17980
rect 29088 17978 29112 17980
rect 29168 17978 29192 17980
rect 29248 17978 29272 17980
rect 29328 17978 29334 17980
rect 29088 17926 29090 17978
rect 29270 17926 29272 17978
rect 29026 17924 29032 17926
rect 29088 17924 29112 17926
rect 29168 17924 29192 17926
rect 29248 17924 29272 17926
rect 29328 17924 29334 17926
rect 29026 17915 29334 17924
rect 27896 17808 27948 17814
rect 27896 17750 27948 17756
rect 28080 17808 28132 17814
rect 28080 17750 28132 17756
rect 28908 17808 28960 17814
rect 28908 17750 28960 17756
rect 26884 17740 26936 17746
rect 26884 17682 26936 17688
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 16794 26372 17478
rect 28366 17436 28674 17445
rect 28366 17434 28372 17436
rect 28428 17434 28452 17436
rect 28508 17434 28532 17436
rect 28588 17434 28612 17436
rect 28668 17434 28674 17436
rect 28428 17382 28430 17434
rect 28610 17382 28612 17434
rect 28366 17380 28372 17382
rect 28428 17380 28452 17382
rect 28508 17380 28532 17382
rect 28588 17380 28612 17382
rect 28668 17380 28674 17382
rect 28366 17371 28674 17380
rect 28920 17338 28948 17750
rect 29380 17678 29408 19110
rect 29564 18970 29592 19178
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29828 18760 29880 18766
rect 29828 18702 29880 18708
rect 29840 18630 29868 18702
rect 29828 18624 29880 18630
rect 29828 18566 29880 18572
rect 29460 18216 29512 18222
rect 29460 18158 29512 18164
rect 29000 17672 29052 17678
rect 29000 17614 29052 17620
rect 29368 17672 29420 17678
rect 29368 17614 29420 17620
rect 28908 17332 28960 17338
rect 28908 17274 28960 17280
rect 29012 17202 29040 17614
rect 29472 17338 29500 18158
rect 29920 17740 29972 17746
rect 29920 17682 29972 17688
rect 29552 17536 29604 17542
rect 29552 17478 29604 17484
rect 29460 17332 29512 17338
rect 29460 17274 29512 17280
rect 29000 17196 29052 17202
rect 29000 17138 29052 17144
rect 27344 17060 27396 17066
rect 27344 17002 27396 17008
rect 26516 16992 26568 16998
rect 26516 16934 26568 16940
rect 27068 16992 27120 16998
rect 27068 16934 27120 16940
rect 26332 16788 26384 16794
rect 26332 16730 26384 16736
rect 26528 16726 26556 16934
rect 27080 16794 27108 16934
rect 27356 16794 27384 17002
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 27068 16788 27120 16794
rect 27068 16730 27120 16736
rect 27344 16788 27396 16794
rect 27344 16730 27396 16736
rect 28920 16726 28948 16934
rect 29026 16892 29334 16901
rect 29026 16890 29032 16892
rect 29088 16890 29112 16892
rect 29168 16890 29192 16892
rect 29248 16890 29272 16892
rect 29328 16890 29334 16892
rect 29088 16838 29090 16890
rect 29270 16838 29272 16890
rect 29026 16836 29032 16838
rect 29088 16836 29112 16838
rect 29168 16836 29192 16838
rect 29248 16836 29272 16838
rect 29328 16836 29334 16838
rect 29026 16827 29334 16836
rect 29564 16726 29592 17478
rect 29932 17338 29960 17682
rect 29920 17332 29972 17338
rect 29920 17274 29972 17280
rect 26516 16720 26568 16726
rect 26516 16662 26568 16668
rect 28908 16720 28960 16726
rect 28908 16662 28960 16668
rect 29552 16720 29604 16726
rect 29552 16662 29604 16668
rect 29368 16584 29420 16590
rect 29368 16526 29420 16532
rect 28366 16348 28674 16357
rect 28366 16346 28372 16348
rect 28428 16346 28452 16348
rect 28508 16346 28532 16348
rect 28588 16346 28612 16348
rect 28668 16346 28674 16348
rect 28428 16294 28430 16346
rect 28610 16294 28612 16346
rect 28366 16292 28372 16294
rect 28428 16292 28452 16294
rect 28508 16292 28532 16294
rect 28588 16292 28612 16294
rect 28668 16292 28674 16294
rect 28366 16283 28674 16292
rect 29380 16114 29408 16526
rect 30024 16250 30052 19654
rect 30208 18834 30236 21490
rect 30656 20256 30708 20262
rect 30656 20198 30708 20204
rect 30668 19961 30696 20198
rect 30654 19952 30710 19961
rect 30654 19887 30656 19896
rect 30708 19887 30710 19896
rect 30656 19858 30708 19864
rect 30654 19816 30710 19825
rect 30654 19751 30710 19760
rect 30668 19718 30696 19751
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30288 19236 30340 19242
rect 30288 19178 30340 19184
rect 30300 18970 30328 19178
rect 30288 18964 30340 18970
rect 30288 18906 30340 18912
rect 30196 18828 30248 18834
rect 30196 18770 30248 18776
rect 30288 18284 30340 18290
rect 30288 18226 30340 18232
rect 30012 16244 30064 16250
rect 30012 16186 30064 16192
rect 29368 16108 29420 16114
rect 29368 16050 29420 16056
rect 29828 16108 29880 16114
rect 29828 16050 29880 16056
rect 26608 16040 26660 16046
rect 26608 15982 26660 15988
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26056 15632 26108 15638
rect 26056 15574 26108 15580
rect 26068 14958 26096 15574
rect 26344 15026 26372 15846
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 25872 14952 25924 14958
rect 25872 14894 25924 14900
rect 26056 14952 26108 14958
rect 26056 14894 26108 14900
rect 25884 14618 25912 14894
rect 25872 14612 25924 14618
rect 25872 14554 25924 14560
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25792 14074 25820 14350
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25884 13954 25912 14554
rect 26068 14550 26096 14894
rect 26056 14544 26108 14550
rect 26056 14486 26108 14492
rect 25792 13926 25912 13954
rect 25792 12782 25820 13926
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25884 13530 25912 13806
rect 25872 13524 25924 13530
rect 25872 13466 25924 13472
rect 26068 12850 26096 14486
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 13870 26188 14214
rect 26620 14074 26648 15982
rect 29026 15804 29334 15813
rect 29026 15802 29032 15804
rect 29088 15802 29112 15804
rect 29168 15802 29192 15804
rect 29248 15802 29272 15804
rect 29328 15802 29334 15804
rect 29088 15750 29090 15802
rect 29270 15750 29272 15802
rect 29026 15748 29032 15750
rect 29088 15748 29112 15750
rect 29168 15748 29192 15750
rect 29248 15748 29272 15750
rect 29328 15748 29334 15750
rect 29026 15739 29334 15748
rect 27804 15632 27856 15638
rect 27804 15574 27856 15580
rect 26884 15496 26936 15502
rect 26884 15438 26936 15444
rect 26896 15162 26924 15438
rect 26884 15156 26936 15162
rect 26884 15098 26936 15104
rect 27816 14618 27844 15574
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 28172 15360 28224 15366
rect 28172 15302 28224 15308
rect 27896 14816 27948 14822
rect 27896 14758 27948 14764
rect 27160 14612 27212 14618
rect 27160 14554 27212 14560
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27172 14074 27200 14554
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 27712 14476 27764 14482
rect 27712 14418 27764 14424
rect 27344 14272 27396 14278
rect 27344 14214 27396 14220
rect 26608 14068 26660 14074
rect 26608 14010 26660 14016
rect 27160 14068 27212 14074
rect 27160 14010 27212 14016
rect 27356 13870 27384 14214
rect 27540 14006 27568 14418
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27528 14000 27580 14006
rect 27528 13942 27580 13948
rect 26148 13864 26200 13870
rect 26148 13806 26200 13812
rect 27344 13864 27396 13870
rect 27344 13806 27396 13812
rect 26160 12889 26188 13806
rect 26976 13796 27028 13802
rect 26976 13738 27028 13744
rect 26988 13462 27016 13738
rect 26976 13456 27028 13462
rect 26976 13398 27028 13404
rect 26424 13320 26476 13326
rect 26424 13262 26476 13268
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26146 12880 26202 12889
rect 26056 12844 26108 12850
rect 26146 12815 26202 12824
rect 26332 12844 26384 12850
rect 26056 12786 26108 12792
rect 26332 12786 26384 12792
rect 25780 12776 25832 12782
rect 25780 12718 25832 12724
rect 23756 12436 23808 12442
rect 23756 12378 23808 12384
rect 23940 12436 23992 12442
rect 23940 12378 23992 12384
rect 24124 12436 24176 12442
rect 24124 12378 24176 12384
rect 24860 12436 24912 12442
rect 24860 12378 24912 12384
rect 25688 12436 25740 12442
rect 25688 12378 25740 12384
rect 23480 12368 23532 12374
rect 23480 12310 23532 12316
rect 22836 12300 22888 12306
rect 22836 12242 22888 12248
rect 23388 12300 23440 12306
rect 23388 12242 23440 12248
rect 22848 12102 22876 12242
rect 23768 12238 23796 12378
rect 23756 12232 23808 12238
rect 23756 12174 23808 12180
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 23480 12096 23532 12102
rect 23480 12038 23532 12044
rect 22848 11370 22876 12038
rect 23492 11898 23520 12038
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22756 11342 22876 11370
rect 22100 11212 22152 11218
rect 22100 11154 22152 11160
rect 22376 11212 22428 11218
rect 22376 11154 22428 11160
rect 22008 10532 22060 10538
rect 22008 10474 22060 10480
rect 21666 10364 21974 10373
rect 21666 10362 21672 10364
rect 21728 10362 21752 10364
rect 21808 10362 21832 10364
rect 21888 10362 21912 10364
rect 21968 10362 21974 10364
rect 21728 10310 21730 10362
rect 21910 10310 21912 10362
rect 21666 10308 21672 10310
rect 21728 10308 21752 10310
rect 21808 10308 21832 10310
rect 21888 10308 21912 10310
rect 21968 10308 21974 10310
rect 21666 10299 21974 10308
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 21836 9489 21864 9658
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21928 9518 21956 9590
rect 21916 9512 21968 9518
rect 21822 9480 21878 9489
rect 21916 9454 21968 9460
rect 21822 9415 21878 9424
rect 21666 9276 21974 9285
rect 21666 9274 21672 9276
rect 21728 9274 21752 9276
rect 21808 9274 21832 9276
rect 21888 9274 21912 9276
rect 21968 9274 21974 9276
rect 21728 9222 21730 9274
rect 21910 9222 21912 9274
rect 21666 9220 21672 9222
rect 21728 9220 21752 9222
rect 21808 9220 21832 9222
rect 21888 9220 21912 9222
rect 21968 9220 21974 9222
rect 21666 9211 21974 9220
rect 21732 8832 21784 8838
rect 21732 8774 21784 8780
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21744 8430 21772 8774
rect 21928 8634 21956 8774
rect 22020 8634 22048 10474
rect 22112 9518 22140 11154
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22100 9512 22152 9518
rect 22100 9454 22152 9460
rect 21916 8628 21968 8634
rect 21916 8570 21968 8576
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 22204 8498 22232 11086
rect 22284 10600 22336 10606
rect 22284 10542 22336 10548
rect 22296 10266 22324 10542
rect 22388 10470 22416 11154
rect 22376 10464 22428 10470
rect 22376 10406 22428 10412
rect 22284 10260 22336 10266
rect 22284 10202 22336 10208
rect 22388 10062 22416 10406
rect 22376 10056 22428 10062
rect 22376 9998 22428 10004
rect 22284 9512 22336 9518
rect 22388 9500 22416 9998
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 22336 9472 22416 9500
rect 22480 9489 22508 9590
rect 22466 9480 22522 9489
rect 22284 9454 22336 9460
rect 22192 8492 22244 8498
rect 22192 8434 22244 8440
rect 21732 8424 21784 8430
rect 21730 8392 21732 8401
rect 21784 8392 21786 8401
rect 22296 8378 22324 9454
rect 22466 9415 22522 9424
rect 21548 8356 21600 8362
rect 21730 8327 21786 8336
rect 22008 8356 22060 8362
rect 21548 8298 21600 8304
rect 22008 8298 22060 8304
rect 22112 8350 22324 8378
rect 21666 8188 21974 8197
rect 21666 8186 21672 8188
rect 21728 8186 21752 8188
rect 21808 8186 21832 8188
rect 21888 8186 21912 8188
rect 21968 8186 21974 8188
rect 21728 8134 21730 8186
rect 21910 8134 21912 8186
rect 21666 8132 21672 8134
rect 21728 8132 21752 8134
rect 21808 8132 21832 8134
rect 21888 8132 21912 8134
rect 21968 8132 21974 8134
rect 21666 8123 21974 8132
rect 21916 7880 21968 7886
rect 22020 7868 22048 8298
rect 22112 8022 22140 8350
rect 22192 8288 22244 8294
rect 22192 8230 22244 8236
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 21968 7840 22048 7868
rect 21916 7822 21968 7828
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21916 7404 21968 7410
rect 21968 7364 22048 7392
rect 21916 7346 21968 7352
rect 21666 7100 21974 7109
rect 21666 7098 21672 7100
rect 21728 7098 21752 7100
rect 21808 7098 21832 7100
rect 21888 7098 21912 7100
rect 21968 7098 21974 7100
rect 21728 7046 21730 7098
rect 21910 7046 21912 7098
rect 21666 7044 21672 7046
rect 21728 7044 21752 7046
rect 21808 7044 21832 7046
rect 21888 7044 21912 7046
rect 21968 7044 21974 7046
rect 21666 7035 21974 7044
rect 22020 6914 22048 7364
rect 22204 7274 22232 8230
rect 22480 7750 22508 9415
rect 22572 7954 22600 9658
rect 22756 9654 22784 11342
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22940 9450 22968 10678
rect 23204 10600 23256 10606
rect 23204 10542 23256 10548
rect 23020 10464 23072 10470
rect 23020 10406 23072 10412
rect 22928 9444 22980 9450
rect 22928 9386 22980 9392
rect 22560 7948 22612 7954
rect 22560 7890 22612 7896
rect 22940 7818 22968 9386
rect 23032 7954 23060 10406
rect 23216 9722 23244 10542
rect 23664 10532 23716 10538
rect 23664 10474 23716 10480
rect 23388 10124 23440 10130
rect 23388 10066 23440 10072
rect 23204 9716 23256 9722
rect 23204 9658 23256 9664
rect 23400 9450 23428 10066
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23492 9518 23520 9862
rect 23584 9654 23612 9998
rect 23572 9648 23624 9654
rect 23570 9616 23572 9625
rect 23624 9616 23626 9625
rect 23570 9551 23626 9560
rect 23676 9518 23704 10474
rect 23480 9512 23532 9518
rect 23664 9512 23716 9518
rect 23480 9454 23532 9460
rect 23662 9480 23664 9489
rect 23716 9480 23718 9489
rect 23388 9444 23440 9450
rect 23662 9415 23718 9424
rect 23388 9386 23440 9392
rect 23768 8838 23796 10746
rect 24136 10606 24164 12378
rect 24582 12200 24638 12209
rect 24582 12135 24638 12144
rect 24490 11928 24546 11937
rect 24490 11863 24546 11872
rect 24504 11830 24532 11863
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 24492 11824 24544 11830
rect 24492 11766 24544 11772
rect 24124 10600 24176 10606
rect 24124 10542 24176 10548
rect 24136 10198 24164 10542
rect 24124 10192 24176 10198
rect 24124 10134 24176 10140
rect 24136 9722 24164 10134
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23860 9042 23888 9454
rect 23940 9444 23992 9450
rect 23940 9386 23992 9392
rect 23952 9178 23980 9386
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 23848 9036 23900 9042
rect 23848 8978 23900 8984
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23296 8424 23348 8430
rect 23296 8366 23348 8372
rect 23386 8392 23442 8401
rect 23112 8288 23164 8294
rect 23112 8230 23164 8236
rect 23124 7954 23152 8230
rect 23308 8090 23336 8366
rect 23386 8327 23442 8336
rect 23400 8294 23428 8327
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23112 7948 23164 7954
rect 23112 7890 23164 7896
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22560 7540 22612 7546
rect 22560 7482 22612 7488
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22572 7206 22600 7482
rect 22652 7268 22704 7274
rect 22652 7210 22704 7216
rect 22560 7200 22612 7206
rect 22560 7142 22612 7148
rect 22664 7002 22692 7210
rect 22652 6996 22704 7002
rect 22652 6938 22704 6944
rect 22940 6934 22968 7754
rect 23400 7546 23428 8230
rect 23480 7880 23532 7886
rect 24228 7834 24256 11766
rect 24596 11694 24624 12135
rect 24872 11694 24900 12378
rect 24952 12300 25004 12306
rect 24952 12242 25004 12248
rect 25688 12300 25740 12306
rect 25688 12242 25740 12248
rect 24964 11830 24992 12242
rect 25136 12096 25188 12102
rect 25136 12038 25188 12044
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 24964 11694 24992 11766
rect 25148 11694 25176 12038
rect 24584 11688 24636 11694
rect 24584 11630 24636 11636
rect 24860 11688 24912 11694
rect 24860 11630 24912 11636
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 25136 11688 25188 11694
rect 25413 11688 25465 11694
rect 25136 11630 25188 11636
rect 25332 11648 25413 11676
rect 25136 11552 25188 11558
rect 25136 11494 25188 11500
rect 25228 11552 25280 11558
rect 25228 11494 25280 11500
rect 25148 11286 25176 11494
rect 25136 11280 25188 11286
rect 25136 11222 25188 11228
rect 25136 11144 25188 11150
rect 25136 11086 25188 11092
rect 24400 11008 24452 11014
rect 24400 10950 24452 10956
rect 24412 10470 24440 10950
rect 25148 10810 25176 11086
rect 25136 10804 25188 10810
rect 25136 10746 25188 10752
rect 25240 10674 25268 11494
rect 25332 11014 25360 11648
rect 25700 11642 25728 12242
rect 25413 11630 25465 11636
rect 25608 11626 25728 11642
rect 25504 11620 25556 11626
rect 25504 11562 25556 11568
rect 25596 11620 25728 11626
rect 25648 11614 25728 11620
rect 25596 11562 25648 11568
rect 25412 11280 25464 11286
rect 25516 11268 25544 11562
rect 25464 11240 25544 11268
rect 25412 11222 25464 11228
rect 25320 11008 25372 11014
rect 25320 10950 25372 10956
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 24860 10532 24912 10538
rect 24860 10474 24912 10480
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24400 10464 24452 10470
rect 24400 10406 24452 10412
rect 24320 9722 24348 10406
rect 24308 9716 24360 9722
rect 24308 9658 24360 9664
rect 24320 8974 24348 9658
rect 24412 9382 24440 10406
rect 24872 10130 24900 10474
rect 25504 10192 25556 10198
rect 25504 10134 25556 10140
rect 24860 10124 24912 10130
rect 24860 10066 24912 10072
rect 25412 10124 25464 10130
rect 25412 10066 25464 10072
rect 25424 9654 25452 10066
rect 25516 9674 25544 10134
rect 25792 10130 25820 12718
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26252 12170 26280 12650
rect 26344 12374 26372 12786
rect 26332 12368 26384 12374
rect 26332 12310 26384 12316
rect 26436 12186 26464 13262
rect 26712 12442 26740 13262
rect 26792 13184 26844 13190
rect 26792 13126 26844 13132
rect 26804 12986 26832 13126
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 26884 12980 26936 12986
rect 26884 12922 26936 12928
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26896 12374 26924 12922
rect 26988 12434 27016 13398
rect 27632 13326 27660 14350
rect 27724 14074 27752 14418
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27712 14068 27764 14074
rect 27712 14010 27764 14016
rect 27816 13938 27844 14282
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27620 13320 27672 13326
rect 27620 13262 27672 13268
rect 27632 12714 27660 13262
rect 27816 12850 27844 13874
rect 27908 13870 27936 14758
rect 28000 14414 28028 15302
rect 28080 15020 28132 15026
rect 28080 14962 28132 14968
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27896 13864 27948 13870
rect 27896 13806 27948 13812
rect 27804 12844 27856 12850
rect 27804 12786 27856 12792
rect 27908 12730 27936 13806
rect 27988 13728 28040 13734
rect 27988 13670 28040 13676
rect 28000 13258 28028 13670
rect 27988 13252 28040 13258
rect 27988 13194 28040 13200
rect 27620 12708 27672 12714
rect 27620 12650 27672 12656
rect 27724 12702 27936 12730
rect 26988 12406 27108 12434
rect 26608 12368 26660 12374
rect 26608 12310 26660 12316
rect 26884 12368 26936 12374
rect 26884 12310 26936 12316
rect 27080 12322 27108 12406
rect 26620 12209 26648 12310
rect 26976 12300 27028 12306
rect 27080 12294 27660 12322
rect 26976 12242 27028 12248
rect 26148 12164 26200 12170
rect 26148 12106 26200 12112
rect 26240 12164 26292 12170
rect 26240 12106 26292 12112
rect 26344 12158 26464 12186
rect 26606 12200 26662 12209
rect 25872 12096 25924 12102
rect 25872 12038 25924 12044
rect 26160 12050 26188 12106
rect 26344 12050 26372 12158
rect 26606 12135 26662 12144
rect 25884 11694 25912 12038
rect 26160 12022 26372 12050
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 25872 11688 25924 11694
rect 26252 11642 26280 12022
rect 26620 11898 26648 12038
rect 26608 11892 26660 11898
rect 26608 11834 26660 11840
rect 26988 11694 27016 12242
rect 27436 12232 27488 12238
rect 27436 12174 27488 12180
rect 27448 11898 27476 12174
rect 27436 11892 27488 11898
rect 27436 11834 27488 11840
rect 27252 11824 27304 11830
rect 27252 11766 27304 11772
rect 25872 11630 25924 11636
rect 26160 11626 26280 11642
rect 26976 11688 27028 11694
rect 26976 11630 27028 11636
rect 26148 11620 26280 11626
rect 26200 11614 26280 11620
rect 26424 11620 26476 11626
rect 26148 11562 26200 11568
rect 26424 11562 26476 11568
rect 26884 11620 26936 11626
rect 26884 11562 26936 11568
rect 26160 10146 26188 11562
rect 26332 11552 26384 11558
rect 26332 11494 26384 11500
rect 26240 11212 26292 11218
rect 26240 11154 26292 11160
rect 26252 10266 26280 11154
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 25780 10124 25832 10130
rect 26160 10118 26280 10146
rect 25780 10066 25832 10072
rect 25412 9648 25464 9654
rect 25516 9646 25728 9674
rect 25412 9590 25464 9596
rect 25700 9518 25728 9646
rect 24768 9512 24820 9518
rect 24768 9454 24820 9460
rect 25228 9512 25280 9518
rect 25228 9454 25280 9460
rect 25688 9512 25740 9518
rect 25740 9472 25820 9500
rect 26252 9489 26280 10118
rect 25688 9454 25740 9460
rect 24584 9444 24636 9450
rect 24584 9386 24636 9392
rect 24400 9376 24452 9382
rect 24400 9318 24452 9324
rect 24412 9110 24440 9318
rect 24400 9104 24452 9110
rect 24400 9046 24452 9052
rect 24308 8968 24360 8974
rect 24308 8910 24360 8916
rect 24320 8430 24348 8910
rect 24596 8430 24624 9386
rect 24780 9042 24808 9454
rect 25136 9444 25188 9450
rect 25136 9386 25188 9392
rect 24768 9036 24820 9042
rect 24768 8978 24820 8984
rect 24952 9036 25004 9042
rect 24952 8978 25004 8984
rect 24676 8968 24728 8974
rect 24964 8922 24992 8978
rect 24676 8910 24728 8916
rect 24688 8498 24716 8910
rect 24780 8894 24992 8922
rect 24676 8492 24728 8498
rect 24676 8434 24728 8440
rect 24308 8424 24360 8430
rect 24308 8366 24360 8372
rect 24584 8424 24636 8430
rect 24584 8366 24636 8372
rect 24780 7954 24808 8894
rect 25148 8634 25176 9386
rect 25240 8838 25268 9454
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25424 9178 25452 9318
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25688 9036 25740 9042
rect 25688 8978 25740 8984
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25700 8634 25728 8978
rect 25792 8838 25820 9472
rect 26238 9480 26294 9489
rect 26344 9450 26372 11494
rect 26436 11354 26464 11562
rect 26424 11348 26476 11354
rect 26424 11290 26476 11296
rect 26896 11286 26924 11562
rect 26884 11280 26936 11286
rect 26884 11222 26936 11228
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 26424 10600 26476 10606
rect 26424 10542 26476 10548
rect 26436 10266 26464 10542
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26896 10130 26924 11222
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27080 10810 27108 11086
rect 27068 10804 27120 10810
rect 27068 10746 27120 10752
rect 27172 10674 27200 11222
rect 27160 10668 27212 10674
rect 27160 10610 27212 10616
rect 27264 10130 27292 11766
rect 27448 11694 27476 11834
rect 27436 11688 27488 11694
rect 27436 11630 27488 11636
rect 27632 10198 27660 12294
rect 27724 11914 27752 12702
rect 27804 12640 27856 12646
rect 27804 12582 27856 12588
rect 27816 12306 27844 12582
rect 27804 12300 27856 12306
rect 27804 12242 27856 12248
rect 27724 11886 27844 11914
rect 27816 11694 27844 11886
rect 28000 11694 28028 13194
rect 28092 12714 28120 14962
rect 28184 12850 28212 15302
rect 28366 15260 28674 15269
rect 28366 15258 28372 15260
rect 28428 15258 28452 15260
rect 28508 15258 28532 15260
rect 28588 15258 28612 15260
rect 28668 15258 28674 15260
rect 28428 15206 28430 15258
rect 28610 15206 28612 15258
rect 28366 15204 28372 15206
rect 28428 15204 28452 15206
rect 28508 15204 28532 15206
rect 28588 15204 28612 15206
rect 28668 15204 28674 15206
rect 28366 15195 28674 15204
rect 28448 14952 28500 14958
rect 28448 14894 28500 14900
rect 28632 14952 28684 14958
rect 28632 14894 28684 14900
rect 28460 14618 28488 14894
rect 28540 14884 28592 14890
rect 28540 14826 28592 14832
rect 28552 14618 28580 14826
rect 28448 14612 28500 14618
rect 28448 14554 28500 14560
rect 28540 14612 28592 14618
rect 28540 14554 28592 14560
rect 28644 14482 28672 14894
rect 29026 14716 29334 14725
rect 29026 14714 29032 14716
rect 29088 14714 29112 14716
rect 29168 14714 29192 14716
rect 29248 14714 29272 14716
rect 29328 14714 29334 14716
rect 29088 14662 29090 14714
rect 29270 14662 29272 14714
rect 29026 14660 29032 14662
rect 29088 14660 29112 14662
rect 29168 14660 29192 14662
rect 29248 14660 29272 14662
rect 29328 14660 29334 14662
rect 29026 14651 29334 14660
rect 28816 14544 28868 14550
rect 28816 14486 28868 14492
rect 28632 14476 28684 14482
rect 28684 14436 28764 14464
rect 28632 14418 28684 14424
rect 28366 14172 28674 14181
rect 28366 14170 28372 14172
rect 28428 14170 28452 14172
rect 28508 14170 28532 14172
rect 28588 14170 28612 14172
rect 28668 14170 28674 14172
rect 28428 14118 28430 14170
rect 28610 14118 28612 14170
rect 28366 14116 28372 14118
rect 28428 14116 28452 14118
rect 28508 14116 28532 14118
rect 28588 14116 28612 14118
rect 28668 14116 28674 14118
rect 28366 14107 28674 14116
rect 28736 13954 28764 14436
rect 28828 14006 28856 14486
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 28908 14340 28960 14346
rect 28908 14282 28960 14288
rect 28644 13926 28764 13954
rect 28816 14000 28868 14006
rect 28816 13942 28868 13948
rect 28644 13870 28672 13926
rect 28632 13864 28684 13870
rect 28632 13806 28684 13812
rect 28724 13864 28776 13870
rect 28920 13852 28948 14282
rect 29288 14074 29316 14350
rect 29380 14074 29408 16050
rect 29736 14952 29788 14958
rect 29736 14894 29788 14900
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 29472 14090 29500 14758
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29472 14074 29592 14090
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 29368 14068 29420 14074
rect 29368 14010 29420 14016
rect 29472 14068 29604 14074
rect 29472 14062 29552 14068
rect 28776 13824 28948 13852
rect 29000 13864 29052 13870
rect 28998 13832 29000 13841
rect 29052 13832 29054 13841
rect 28724 13806 28776 13812
rect 28644 13462 28672 13806
rect 28632 13456 28684 13462
rect 28632 13398 28684 13404
rect 28736 13190 28764 13806
rect 28998 13767 29054 13776
rect 29026 13628 29334 13637
rect 29026 13626 29032 13628
rect 29088 13626 29112 13628
rect 29168 13626 29192 13628
rect 29248 13626 29272 13628
rect 29328 13626 29334 13628
rect 29088 13574 29090 13626
rect 29270 13574 29272 13626
rect 29026 13572 29032 13574
rect 29088 13572 29112 13574
rect 29168 13572 29192 13574
rect 29248 13572 29272 13574
rect 29328 13572 29334 13574
rect 29026 13563 29334 13572
rect 29380 13462 29408 14010
rect 29368 13456 29420 13462
rect 29012 13394 29132 13410
rect 29368 13398 29420 13404
rect 29000 13388 29132 13394
rect 29052 13382 29132 13388
rect 29000 13330 29052 13336
rect 28998 13288 29054 13297
rect 28998 13223 29000 13232
rect 29052 13223 29054 13232
rect 29000 13194 29052 13200
rect 28448 13184 28500 13190
rect 28276 13144 28448 13172
rect 28172 12844 28224 12850
rect 28172 12786 28224 12792
rect 28080 12708 28132 12714
rect 28080 12650 28132 12656
rect 28172 12640 28224 12646
rect 28172 12582 28224 12588
rect 28184 11694 28212 12582
rect 27712 11688 27764 11694
rect 27712 11630 27764 11636
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27988 11688 28040 11694
rect 27988 11630 28040 11636
rect 28172 11688 28224 11694
rect 28172 11630 28224 11636
rect 27724 11014 27752 11630
rect 27804 11552 27856 11558
rect 27804 11494 27856 11500
rect 28080 11552 28132 11558
rect 28080 11494 28132 11500
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27620 10192 27672 10198
rect 27620 10134 27672 10140
rect 26884 10124 26936 10130
rect 26884 10066 26936 10072
rect 27252 10124 27304 10130
rect 27252 10066 27304 10072
rect 27264 9722 27292 10066
rect 27724 10062 27752 10950
rect 27816 10198 27844 11494
rect 28092 10266 28120 11494
rect 28080 10260 28132 10266
rect 28080 10202 28132 10208
rect 27804 10192 27856 10198
rect 27804 10134 27856 10140
rect 28172 10192 28224 10198
rect 28172 10134 28224 10140
rect 27712 10056 27764 10062
rect 27712 9998 27764 10004
rect 27436 9920 27488 9926
rect 27436 9862 27488 9868
rect 26608 9716 26660 9722
rect 26608 9658 26660 9664
rect 27252 9716 27304 9722
rect 27252 9658 27304 9664
rect 26620 9518 26648 9658
rect 26608 9512 26660 9518
rect 26608 9454 26660 9460
rect 26238 9415 26240 9424
rect 26292 9415 26294 9424
rect 26332 9444 26384 9450
rect 26240 9386 26292 9392
rect 26332 9386 26384 9392
rect 26976 9444 27028 9450
rect 26976 9386 27028 9392
rect 25872 9376 25924 9382
rect 25872 9318 25924 9324
rect 25884 8974 25912 9318
rect 25872 8968 25924 8974
rect 25872 8910 25924 8916
rect 26344 8838 26372 9386
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26608 9172 26660 9178
rect 26608 9114 26660 9120
rect 26620 9042 26648 9114
rect 26424 9036 26476 9042
rect 26424 8978 26476 8984
rect 26608 9036 26660 9042
rect 26608 8978 26660 8984
rect 25780 8832 25832 8838
rect 25780 8774 25832 8780
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 25136 8628 25188 8634
rect 25136 8570 25188 8576
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25148 8537 25176 8570
rect 25134 8528 25190 8537
rect 26160 8498 26188 8774
rect 25134 8463 25190 8472
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 25320 8424 25372 8430
rect 25320 8366 25372 8372
rect 25872 8424 25924 8430
rect 25872 8366 25924 8372
rect 24768 7948 24820 7954
rect 24768 7890 24820 7896
rect 23480 7822 23532 7828
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 22928 6928 22980 6934
rect 22020 6886 22140 6914
rect 21548 6860 21600 6866
rect 21548 6802 21600 6808
rect 21006 6556 21314 6565
rect 21006 6554 21012 6556
rect 21068 6554 21092 6556
rect 21148 6554 21172 6556
rect 21228 6554 21252 6556
rect 21308 6554 21314 6556
rect 21068 6502 21070 6554
rect 21250 6502 21252 6554
rect 21006 6500 21012 6502
rect 21068 6500 21092 6502
rect 21148 6500 21172 6502
rect 21228 6500 21252 6502
rect 21308 6500 21314 6502
rect 21006 6491 21314 6500
rect 21362 6352 21418 6361
rect 21560 6322 21588 6802
rect 22112 6322 22140 6886
rect 22928 6870 22980 6876
rect 23400 6798 23428 7482
rect 23492 7002 23520 7822
rect 23676 7806 24256 7834
rect 23480 6996 23532 7002
rect 23480 6938 23532 6944
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 21362 6287 21418 6296
rect 21548 6316 21600 6322
rect 21376 5642 21404 6287
rect 21548 6258 21600 6264
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 21560 5914 21588 6258
rect 21666 6012 21974 6021
rect 21666 6010 21672 6012
rect 21728 6010 21752 6012
rect 21808 6010 21832 6012
rect 21888 6010 21912 6012
rect 21968 6010 21974 6012
rect 21728 5958 21730 6010
rect 21910 5958 21912 6010
rect 21666 5956 21672 5958
rect 21728 5956 21752 5958
rect 21808 5956 21832 5958
rect 21888 5956 21912 5958
rect 21968 5956 21974 5958
rect 21666 5947 21974 5956
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21364 5636 21416 5642
rect 21364 5578 21416 5584
rect 21006 5468 21314 5477
rect 21006 5466 21012 5468
rect 21068 5466 21092 5468
rect 21148 5466 21172 5468
rect 21228 5466 21252 5468
rect 21308 5466 21314 5468
rect 21068 5414 21070 5466
rect 21250 5414 21252 5466
rect 21006 5412 21012 5414
rect 21068 5412 21092 5414
rect 21148 5412 21172 5414
rect 21228 5412 21252 5414
rect 21308 5412 21314 5414
rect 21006 5403 21314 5412
rect 21272 5364 21324 5370
rect 21376 5352 21404 5578
rect 21560 5386 21588 5850
rect 21640 5704 21692 5710
rect 21640 5646 21692 5652
rect 21324 5324 21404 5352
rect 21468 5358 21588 5386
rect 21272 5306 21324 5312
rect 21180 5092 21232 5098
rect 21180 5034 21232 5040
rect 21192 4826 21220 5034
rect 21468 4826 21496 5358
rect 21652 5302 21680 5646
rect 21640 5296 21692 5302
rect 21640 5238 21692 5244
rect 22112 5234 22140 6258
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 22560 5840 22612 5846
rect 22560 5782 22612 5788
rect 22744 5840 22796 5846
rect 22744 5782 22796 5788
rect 22572 5574 22600 5782
rect 22756 5681 22784 5782
rect 22742 5672 22798 5681
rect 22742 5607 22798 5616
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22560 5568 22612 5574
rect 22560 5510 22612 5516
rect 21548 5228 21600 5234
rect 21548 5170 21600 5176
rect 22100 5228 22152 5234
rect 22100 5170 22152 5176
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21456 4820 21508 4826
rect 21456 4762 21508 4768
rect 21560 4690 21588 5170
rect 22388 5166 22416 5510
rect 22008 5160 22060 5166
rect 22008 5102 22060 5108
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 21666 4924 21974 4933
rect 21666 4922 21672 4924
rect 21728 4922 21752 4924
rect 21808 4922 21832 4924
rect 21888 4922 21912 4924
rect 21968 4922 21974 4924
rect 21728 4870 21730 4922
rect 21910 4870 21912 4922
rect 21666 4868 21672 4870
rect 21728 4868 21752 4870
rect 21808 4868 21832 4870
rect 21888 4868 21912 4870
rect 21968 4868 21974 4870
rect 21666 4859 21974 4868
rect 22020 4826 22048 5102
rect 23584 4826 23612 6190
rect 23676 5574 23704 7806
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 24136 7342 24164 7686
rect 24124 7336 24176 7342
rect 24124 7278 24176 7284
rect 24504 7274 24532 7686
rect 24492 7268 24544 7274
rect 24492 7210 24544 7216
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23860 5914 23888 6802
rect 24676 6656 24728 6662
rect 24676 6598 24728 6604
rect 24688 6458 24716 6598
rect 24676 6452 24728 6458
rect 24676 6394 24728 6400
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 23940 6112 23992 6118
rect 23940 6054 23992 6060
rect 24032 6112 24084 6118
rect 24032 6054 24084 6060
rect 23952 5914 23980 6054
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23664 5568 23716 5574
rect 23664 5510 23716 5516
rect 23676 5030 23704 5510
rect 23768 5030 23796 5850
rect 24044 5370 24072 6054
rect 24596 5914 24624 6190
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24492 5568 24544 5574
rect 24492 5510 24544 5516
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24032 5364 24084 5370
rect 24032 5306 24084 5312
rect 23664 5024 23716 5030
rect 23664 4966 23716 4972
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23952 4826 23980 5306
rect 24216 5228 24268 5234
rect 24216 5170 24268 5176
rect 24124 5160 24176 5166
rect 24044 5120 24124 5148
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 23572 4820 23624 4826
rect 23572 4762 23624 4768
rect 23940 4820 23992 4826
rect 23940 4762 23992 4768
rect 23112 4752 23164 4758
rect 23112 4694 23164 4700
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21006 4380 21314 4389
rect 21006 4378 21012 4380
rect 21068 4378 21092 4380
rect 21148 4378 21172 4380
rect 21228 4378 21252 4380
rect 21308 4378 21314 4380
rect 21068 4326 21070 4378
rect 21250 4326 21252 4378
rect 21006 4324 21012 4326
rect 21068 4324 21092 4326
rect 21148 4324 21172 4326
rect 21228 4324 21252 4326
rect 21308 4324 21314 4326
rect 21006 4315 21314 4324
rect 21560 4146 21588 4626
rect 20904 4140 20956 4146
rect 20904 4082 20956 4088
rect 21548 4140 21600 4146
rect 21548 4082 21600 4088
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 20916 3602 20944 4082
rect 21180 4004 21232 4010
rect 21180 3946 21232 3952
rect 21192 3738 21220 3946
rect 21836 3942 21864 4082
rect 21824 3936 21876 3942
rect 21824 3878 21876 3884
rect 22192 3936 22244 3942
rect 22192 3878 22244 3884
rect 21666 3836 21974 3845
rect 21666 3834 21672 3836
rect 21728 3834 21752 3836
rect 21808 3834 21832 3836
rect 21888 3834 21912 3836
rect 21968 3834 21974 3836
rect 21728 3782 21730 3834
rect 21910 3782 21912 3834
rect 21666 3780 21672 3782
rect 21728 3780 21752 3782
rect 21808 3780 21832 3782
rect 21888 3780 21912 3782
rect 21968 3780 21974 3782
rect 21666 3771 21974 3780
rect 22204 3738 22232 3878
rect 23124 3738 23152 4694
rect 23480 4684 23532 4690
rect 23480 4626 23532 4632
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 23400 4282 23428 4422
rect 23388 4276 23440 4282
rect 23388 4218 23440 4224
rect 23492 4162 23520 4626
rect 24044 4622 24072 5120
rect 24124 5102 24176 5108
rect 24228 4706 24256 5170
rect 24136 4690 24256 4706
rect 24504 4690 24532 5510
rect 24780 5302 24808 7890
rect 25332 7206 25360 8366
rect 25780 8288 25832 8294
rect 25780 8230 25832 8236
rect 25792 8022 25820 8230
rect 25780 8016 25832 8022
rect 25884 7993 25912 8366
rect 26436 8090 26464 8978
rect 26620 8362 26648 8978
rect 26896 8566 26924 9318
rect 26884 8560 26936 8566
rect 26884 8502 26936 8508
rect 26988 8430 27016 9386
rect 27068 9376 27120 9382
rect 27068 9318 27120 9324
rect 27080 9178 27108 9318
rect 27264 9178 27292 9658
rect 27448 9654 27476 9862
rect 27816 9722 27844 10134
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 27908 9722 27936 9862
rect 27804 9716 27856 9722
rect 27804 9658 27856 9664
rect 27896 9716 27948 9722
rect 27896 9658 27948 9664
rect 27436 9648 27488 9654
rect 27436 9590 27488 9596
rect 27448 9178 27476 9590
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27526 9480 27582 9489
rect 27724 9466 27752 9522
rect 28000 9466 28028 9998
rect 28184 9586 28212 10134
rect 28276 9926 28304 13144
rect 28448 13126 28500 13132
rect 28724 13184 28776 13190
rect 28724 13126 28776 13132
rect 28366 13084 28674 13093
rect 28366 13082 28372 13084
rect 28428 13082 28452 13084
rect 28508 13082 28532 13084
rect 28588 13082 28612 13084
rect 28668 13082 28674 13084
rect 28428 13030 28430 13082
rect 28610 13030 28612 13082
rect 28366 13028 28372 13030
rect 28428 13028 28452 13030
rect 28508 13028 28532 13030
rect 28588 13028 28612 13030
rect 28668 13028 28674 13030
rect 28366 13019 28674 13028
rect 28356 12776 28408 12782
rect 28356 12718 28408 12724
rect 28368 12374 28396 12718
rect 28632 12640 28684 12646
rect 28632 12582 28684 12588
rect 28644 12442 28672 12582
rect 28632 12436 28684 12442
rect 28632 12378 28684 12384
rect 28736 12374 28764 13126
rect 28906 12880 28962 12889
rect 29104 12850 29132 13382
rect 29472 13138 29500 14062
rect 29552 14010 29604 14016
rect 29550 13832 29606 13841
rect 29550 13767 29606 13776
rect 29288 13110 29500 13138
rect 28906 12815 28962 12824
rect 29092 12844 29144 12850
rect 28816 12708 28868 12714
rect 28816 12650 28868 12656
rect 28356 12368 28408 12374
rect 28356 12310 28408 12316
rect 28724 12368 28776 12374
rect 28724 12310 28776 12316
rect 28828 12102 28856 12650
rect 28920 12434 28948 12815
rect 29092 12786 29144 12792
rect 29288 12714 29316 13110
rect 29460 12980 29512 12986
rect 29460 12922 29512 12928
rect 29276 12708 29328 12714
rect 29276 12650 29328 12656
rect 29026 12540 29334 12549
rect 29026 12538 29032 12540
rect 29088 12538 29112 12540
rect 29168 12538 29192 12540
rect 29248 12538 29272 12540
rect 29328 12538 29334 12540
rect 29088 12486 29090 12538
rect 29270 12486 29272 12538
rect 29026 12484 29032 12486
rect 29088 12484 29112 12486
rect 29168 12484 29192 12486
rect 29248 12484 29272 12486
rect 29328 12484 29334 12486
rect 29026 12475 29334 12484
rect 28920 12406 29224 12434
rect 29196 12306 29224 12406
rect 29184 12300 29236 12306
rect 29184 12242 29236 12248
rect 29196 12102 29224 12242
rect 28816 12096 28868 12102
rect 28816 12038 28868 12044
rect 29184 12096 29236 12102
rect 29184 12038 29236 12044
rect 28366 11996 28674 12005
rect 28366 11994 28372 11996
rect 28428 11994 28452 11996
rect 28508 11994 28532 11996
rect 28588 11994 28612 11996
rect 28668 11994 28674 11996
rect 28428 11942 28430 11994
rect 28610 11942 28612 11994
rect 28366 11940 28372 11942
rect 28428 11940 28452 11942
rect 28508 11940 28532 11942
rect 28588 11940 28612 11942
rect 28668 11940 28674 11942
rect 28366 11931 28674 11940
rect 28828 11778 28856 12038
rect 28644 11750 28856 11778
rect 29472 11762 29500 12922
rect 29564 12374 29592 13767
rect 29656 12714 29684 14214
rect 29748 13297 29776 14894
rect 29840 13682 29868 16050
rect 30196 15972 30248 15978
rect 30196 15914 30248 15920
rect 30208 15706 30236 15914
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 29920 14816 29972 14822
rect 29920 14758 29972 14764
rect 29932 14414 29960 14758
rect 30300 14550 30328 18226
rect 30760 18154 30788 25434
rect 31036 22094 31064 31962
rect 31588 30870 31616 33544
rect 31666 32056 31722 32065
rect 31666 31991 31722 32000
rect 31576 30864 31628 30870
rect 31576 30806 31628 30812
rect 31300 30048 31352 30054
rect 31300 29990 31352 29996
rect 31484 30048 31536 30054
rect 31484 29990 31536 29996
rect 31312 29306 31340 29990
rect 31392 29504 31444 29510
rect 31392 29446 31444 29452
rect 31300 29300 31352 29306
rect 31300 29242 31352 29248
rect 31404 29170 31432 29446
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31300 29028 31352 29034
rect 31300 28970 31352 28976
rect 31116 28756 31168 28762
rect 31116 28698 31168 28704
rect 31128 28150 31156 28698
rect 31208 28552 31260 28558
rect 31208 28494 31260 28500
rect 31116 28144 31168 28150
rect 31116 28086 31168 28092
rect 31220 27878 31248 28494
rect 31208 27872 31260 27878
rect 31208 27814 31260 27820
rect 31116 27600 31168 27606
rect 31116 27542 31168 27548
rect 31128 27441 31156 27542
rect 31312 27538 31340 28970
rect 31300 27532 31352 27538
rect 31300 27474 31352 27480
rect 31114 27432 31170 27441
rect 31114 27367 31170 27376
rect 31312 25294 31340 27474
rect 31404 26790 31432 29106
rect 31392 26784 31444 26790
rect 31392 26726 31444 26732
rect 31404 25498 31432 26726
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31300 25288 31352 25294
rect 31300 25230 31352 25236
rect 31312 23186 31340 25230
rect 31300 23180 31352 23186
rect 31300 23122 31352 23128
rect 31312 22982 31340 23122
rect 31300 22976 31352 22982
rect 31300 22918 31352 22924
rect 30852 22066 31064 22094
rect 30852 19922 30880 22066
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 30840 19916 30892 19922
rect 30840 19858 30892 19864
rect 31220 19786 31248 20198
rect 31496 19854 31524 29990
rect 31680 29782 31708 31991
rect 32600 30938 32628 33646
rect 32862 33544 32918 33646
rect 34150 33544 34206 34344
rect 33138 33416 33194 33425
rect 33138 33351 33194 33360
rect 33152 32026 33180 33351
rect 33140 32020 33192 32026
rect 33140 31962 33192 31968
rect 34164 31346 34192 33544
rect 34152 31340 34204 31346
rect 34152 31282 34204 31288
rect 32588 30932 32640 30938
rect 32588 30874 32640 30880
rect 33046 30696 33102 30705
rect 33046 30631 33102 30640
rect 33060 30258 33088 30631
rect 33048 30252 33100 30258
rect 33048 30194 33100 30200
rect 31668 29776 31720 29782
rect 31668 29718 31720 29724
rect 31668 28960 31720 28966
rect 31668 28902 31720 28908
rect 31680 28694 31708 28902
rect 31668 28688 31720 28694
rect 31668 28630 31720 28636
rect 31852 27872 31904 27878
rect 31852 27814 31904 27820
rect 31864 27606 31892 27814
rect 31852 27600 31904 27606
rect 31852 27542 31904 27548
rect 33138 27296 33194 27305
rect 33138 27231 33194 27240
rect 33152 26926 33180 27231
rect 33140 26920 33192 26926
rect 33140 26862 33192 26868
rect 33140 25288 33192 25294
rect 33138 25256 33140 25265
rect 33192 25256 33194 25265
rect 33138 25191 33194 25200
rect 31576 24200 31628 24206
rect 31576 24142 31628 24148
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 31484 19848 31536 19854
rect 31484 19790 31536 19796
rect 31208 19780 31260 19786
rect 31208 19722 31260 19728
rect 31392 19780 31444 19786
rect 31392 19722 31444 19728
rect 31024 19168 31076 19174
rect 31024 19110 31076 19116
rect 31208 19168 31260 19174
rect 31208 19110 31260 19116
rect 31036 18834 31064 19110
rect 31220 18970 31248 19110
rect 31208 18964 31260 18970
rect 31208 18906 31260 18912
rect 31024 18828 31076 18834
rect 31024 18770 31076 18776
rect 30380 18148 30432 18154
rect 30380 18090 30432 18096
rect 30748 18148 30800 18154
rect 30748 18090 30800 18096
rect 30392 16998 30420 18090
rect 30840 17740 30892 17746
rect 30840 17682 30892 17688
rect 30656 17128 30708 17134
rect 30656 17070 30708 17076
rect 30852 17116 30880 17682
rect 30932 17128 30984 17134
rect 30852 17088 30932 17116
rect 30380 16992 30432 16998
rect 30380 16934 30432 16940
rect 30392 16538 30420 16934
rect 30668 16794 30696 17070
rect 30656 16788 30708 16794
rect 30656 16730 30708 16736
rect 30392 16510 30512 16538
rect 30852 16522 30880 17088
rect 30932 17070 30984 17076
rect 31300 16720 31352 16726
rect 31300 16662 31352 16668
rect 30380 16448 30432 16454
rect 30380 16390 30432 16396
rect 30392 15570 30420 16390
rect 30484 15706 30512 16510
rect 30840 16516 30892 16522
rect 30840 16458 30892 16464
rect 30472 15700 30524 15706
rect 30472 15642 30524 15648
rect 30748 15632 30800 15638
rect 30748 15574 30800 15580
rect 30380 15564 30432 15570
rect 30380 15506 30432 15512
rect 30760 14958 30788 15574
rect 31312 15162 31340 16662
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30748 14952 30800 14958
rect 30748 14894 30800 14900
rect 30840 14884 30892 14890
rect 30840 14826 30892 14832
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 30288 14544 30340 14550
rect 30288 14486 30340 14492
rect 30668 14482 30696 14758
rect 30852 14482 30880 14826
rect 30656 14476 30708 14482
rect 30656 14418 30708 14424
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 29920 14408 29972 14414
rect 29920 14350 29972 14356
rect 29932 13818 29960 14350
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 29932 13790 30144 13818
rect 29840 13654 30052 13682
rect 29734 13288 29790 13297
rect 29734 13223 29790 13232
rect 29644 12708 29696 12714
rect 29644 12650 29696 12656
rect 29748 12442 29776 13223
rect 29828 13184 29880 13190
rect 29828 13126 29880 13132
rect 29840 12714 29868 13126
rect 29828 12708 29880 12714
rect 29828 12650 29880 12656
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29552 12368 29604 12374
rect 29552 12310 29604 12316
rect 29748 12306 29776 12378
rect 29736 12300 29788 12306
rect 29736 12242 29788 12248
rect 29748 11898 29776 12242
rect 29828 12096 29880 12102
rect 29828 12038 29880 12044
rect 29736 11892 29788 11898
rect 29736 11834 29788 11840
rect 29368 11756 29420 11762
rect 28644 11286 28672 11750
rect 29368 11698 29420 11704
rect 29460 11756 29512 11762
rect 29460 11698 29512 11704
rect 28908 11552 28960 11558
rect 28908 11494 28960 11500
rect 28920 11354 28948 11494
rect 29026 11452 29334 11461
rect 29026 11450 29032 11452
rect 29088 11450 29112 11452
rect 29168 11450 29192 11452
rect 29248 11450 29272 11452
rect 29328 11450 29334 11452
rect 29088 11398 29090 11450
rect 29270 11398 29272 11450
rect 29026 11396 29032 11398
rect 29088 11396 29112 11398
rect 29168 11396 29192 11398
rect 29248 11396 29272 11398
rect 29328 11396 29334 11398
rect 29026 11387 29334 11396
rect 29380 11354 29408 11698
rect 28908 11348 28960 11354
rect 28908 11290 28960 11296
rect 29368 11348 29420 11354
rect 29368 11290 29420 11296
rect 28632 11280 28684 11286
rect 28632 11222 28684 11228
rect 29736 11212 29788 11218
rect 29736 11154 29788 11160
rect 28724 11008 28776 11014
rect 28724 10950 28776 10956
rect 28816 11008 28868 11014
rect 28816 10950 28868 10956
rect 28366 10908 28674 10917
rect 28366 10906 28372 10908
rect 28428 10906 28452 10908
rect 28508 10906 28532 10908
rect 28588 10906 28612 10908
rect 28668 10906 28674 10908
rect 28428 10854 28430 10906
rect 28610 10854 28612 10906
rect 28366 10852 28372 10854
rect 28428 10852 28452 10854
rect 28508 10852 28532 10854
rect 28588 10852 28612 10854
rect 28668 10852 28674 10854
rect 28366 10843 28674 10852
rect 28736 10606 28764 10950
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28264 9920 28316 9926
rect 28264 9862 28316 9868
rect 28724 9920 28776 9926
rect 28724 9862 28776 9868
rect 28172 9580 28224 9586
rect 28172 9522 28224 9528
rect 28276 9518 28304 9862
rect 28366 9820 28674 9829
rect 28366 9818 28372 9820
rect 28428 9818 28452 9820
rect 28508 9818 28532 9820
rect 28588 9818 28612 9820
rect 28668 9818 28674 9820
rect 28428 9766 28430 9818
rect 28610 9766 28612 9818
rect 28366 9764 28372 9766
rect 28428 9764 28452 9766
rect 28508 9764 28532 9766
rect 28588 9764 28612 9766
rect 28668 9764 28674 9766
rect 28366 9755 28674 9764
rect 28540 9580 28592 9586
rect 28540 9522 28592 9528
rect 27526 9415 27582 9424
rect 27620 9444 27672 9450
rect 27540 9382 27568 9415
rect 27724 9438 28028 9466
rect 28264 9512 28316 9518
rect 28264 9454 28316 9460
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 27620 9386 27672 9392
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27068 9172 27120 9178
rect 27068 9114 27120 9120
rect 27252 9172 27304 9178
rect 27436 9172 27488 9178
rect 27304 9132 27384 9160
rect 27252 9114 27304 9120
rect 27356 9058 27384 9132
rect 27436 9114 27488 9120
rect 27632 9058 27660 9386
rect 27804 9376 27856 9382
rect 27804 9318 27856 9324
rect 27816 9178 27844 9318
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27896 9172 27948 9178
rect 27896 9114 27948 9120
rect 27356 9030 27660 9058
rect 27908 8922 27936 9114
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 27540 8894 27936 8922
rect 27080 8498 27108 8842
rect 27540 8838 27568 8894
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27528 8560 27580 8566
rect 27528 8502 27580 8508
rect 27068 8492 27120 8498
rect 27068 8434 27120 8440
rect 27540 8430 27568 8502
rect 26976 8424 27028 8430
rect 26976 8366 27028 8372
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 26608 8356 26660 8362
rect 26608 8298 26660 8304
rect 26700 8288 26752 8294
rect 26700 8230 26752 8236
rect 27436 8288 27488 8294
rect 27436 8230 27488 8236
rect 26712 8090 26740 8230
rect 26424 8084 26476 8090
rect 26424 8026 26476 8032
rect 26700 8084 26752 8090
rect 26700 8026 26752 8032
rect 25780 7958 25832 7964
rect 25870 7984 25926 7993
rect 25870 7919 25926 7928
rect 27448 7886 27476 8230
rect 27632 7954 27660 8774
rect 28000 8634 28028 9438
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28368 9178 28396 9318
rect 28460 9178 28488 9454
rect 28356 9172 28408 9178
rect 28356 9114 28408 9120
rect 28448 9172 28500 9178
rect 28448 9114 28500 9120
rect 28080 8968 28132 8974
rect 28080 8910 28132 8916
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 27988 8628 28040 8634
rect 27988 8570 28040 8576
rect 27620 7948 27672 7954
rect 27620 7890 27672 7896
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 26976 7812 27028 7818
rect 26976 7754 27028 7760
rect 26332 7744 26384 7750
rect 26252 7692 26332 7698
rect 26252 7686 26384 7692
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26252 7670 26372 7686
rect 26252 7274 26280 7670
rect 26240 7268 26292 7274
rect 26240 7210 26292 7216
rect 26332 7268 26384 7274
rect 26332 7210 26384 7216
rect 25320 7200 25372 7206
rect 25320 7142 25372 7148
rect 25780 7200 25832 7206
rect 25780 7142 25832 7148
rect 24952 6656 25004 6662
rect 24952 6598 25004 6604
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 24964 5846 24992 6598
rect 25056 5914 25084 6598
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 24952 5840 25004 5846
rect 24952 5782 25004 5788
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25608 5370 25636 5646
rect 25596 5364 25648 5370
rect 25596 5306 25648 5312
rect 24768 5296 24820 5302
rect 24768 5238 24820 5244
rect 24952 5160 25004 5166
rect 24952 5102 25004 5108
rect 24676 5092 24728 5098
rect 24860 5092 24912 5098
rect 24728 5052 24860 5080
rect 24676 5034 24728 5040
rect 24860 5034 24912 5040
rect 24964 4758 24992 5102
rect 24952 4752 25004 4758
rect 24952 4694 25004 4700
rect 24124 4684 24256 4690
rect 24176 4678 24256 4684
rect 24492 4684 24544 4690
rect 24124 4626 24176 4632
rect 24492 4626 24544 4632
rect 24032 4616 24084 4622
rect 24032 4558 24084 4564
rect 23572 4480 23624 4486
rect 23572 4422 23624 4428
rect 23400 4134 23520 4162
rect 23400 3738 23428 4134
rect 23584 3942 23612 4422
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 21180 3732 21232 3738
rect 21180 3674 21232 3680
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 20904 3596 20956 3602
rect 20904 3538 20956 3544
rect 23492 3534 23520 3878
rect 23480 3528 23532 3534
rect 20720 3460 20772 3466
rect 20824 3454 20944 3482
rect 23480 3470 23532 3476
rect 20720 3402 20772 3408
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20916 3194 20944 3454
rect 21006 3292 21314 3301
rect 21006 3290 21012 3292
rect 21068 3290 21092 3292
rect 21148 3290 21172 3292
rect 21228 3290 21252 3292
rect 21308 3290 21314 3292
rect 21068 3238 21070 3290
rect 21250 3238 21252 3290
rect 21006 3236 21012 3238
rect 21068 3236 21092 3238
rect 21148 3236 21172 3238
rect 21228 3236 21252 3238
rect 21308 3236 21314 3238
rect 21006 3227 21314 3236
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19352 1414 19472 1442
rect 19352 800 19380 1414
rect 21284 800 21312 2926
rect 21666 2748 21974 2757
rect 21666 2746 21672 2748
rect 21728 2746 21752 2748
rect 21808 2746 21832 2748
rect 21888 2746 21912 2748
rect 21968 2746 21974 2748
rect 21728 2694 21730 2746
rect 21910 2694 21912 2746
rect 21666 2692 21672 2694
rect 21728 2692 21752 2694
rect 21808 2692 21832 2694
rect 21888 2692 21912 2694
rect 21968 2692 21974 2694
rect 21666 2683 21974 2692
rect 22572 800 22600 2994
rect 23492 2990 23520 3470
rect 23584 2990 23612 3878
rect 24044 3738 24072 4558
rect 25412 4480 25464 4486
rect 25412 4422 25464 4428
rect 25424 4282 25452 4422
rect 25412 4276 25464 4282
rect 25412 4218 25464 4224
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 25792 3602 25820 7142
rect 26252 6322 26280 7210
rect 26344 7002 26372 7210
rect 26896 7002 26924 7686
rect 26988 7206 27016 7754
rect 27632 7274 27660 7890
rect 27712 7880 27764 7886
rect 27712 7822 27764 7828
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27724 7546 27752 7822
rect 27712 7540 27764 7546
rect 27712 7482 27764 7488
rect 27620 7268 27672 7274
rect 27620 7210 27672 7216
rect 26976 7200 27028 7206
rect 26976 7142 27028 7148
rect 27252 7200 27304 7206
rect 27252 7142 27304 7148
rect 26332 6996 26384 7002
rect 26332 6938 26384 6944
rect 26884 6996 26936 7002
rect 26884 6938 26936 6944
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 27264 6186 27292 7142
rect 27632 7002 27660 7210
rect 27816 7002 27844 7822
rect 27620 6996 27672 7002
rect 27620 6938 27672 6944
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 27632 6866 27660 6938
rect 27620 6860 27672 6866
rect 27620 6802 27672 6808
rect 27908 6798 27936 8570
rect 28092 8430 28120 8910
rect 28460 8906 28488 9114
rect 28448 8900 28500 8906
rect 28448 8842 28500 8848
rect 28552 8820 28580 9522
rect 28736 9518 28764 9862
rect 28724 9512 28776 9518
rect 28630 9480 28686 9489
rect 28724 9454 28776 9460
rect 28630 9415 28686 9424
rect 28644 8974 28672 9415
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28552 8792 28764 8820
rect 28366 8732 28674 8741
rect 28366 8730 28372 8732
rect 28428 8730 28452 8732
rect 28508 8730 28532 8732
rect 28588 8730 28612 8732
rect 28668 8730 28674 8732
rect 28428 8678 28430 8730
rect 28610 8678 28612 8730
rect 28366 8676 28372 8678
rect 28428 8676 28452 8678
rect 28508 8676 28532 8678
rect 28588 8676 28612 8678
rect 28668 8676 28674 8678
rect 28366 8667 28674 8676
rect 28446 8528 28502 8537
rect 28446 8463 28502 8472
rect 28460 8430 28488 8463
rect 28736 8430 28764 8792
rect 28828 8634 28856 10950
rect 29460 10804 29512 10810
rect 29460 10746 29512 10752
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29026 10364 29334 10373
rect 29026 10362 29032 10364
rect 29088 10362 29112 10364
rect 29168 10362 29192 10364
rect 29248 10362 29272 10364
rect 29328 10362 29334 10364
rect 29088 10310 29090 10362
rect 29270 10310 29272 10362
rect 29026 10308 29032 10310
rect 29088 10308 29112 10310
rect 29168 10308 29192 10310
rect 29248 10308 29272 10310
rect 29328 10308 29334 10310
rect 29026 10299 29334 10308
rect 28908 10124 28960 10130
rect 28908 10066 28960 10072
rect 29092 10124 29144 10130
rect 29092 10066 29144 10072
rect 28920 9382 28948 10066
rect 29104 9674 29132 10066
rect 29380 10062 29408 10610
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 29000 9648 29052 9654
rect 29104 9646 29224 9674
rect 29000 9590 29052 9596
rect 29012 9382 29040 9590
rect 29196 9489 29224 9646
rect 29182 9480 29238 9489
rect 29182 9415 29184 9424
rect 29236 9415 29238 9424
rect 29184 9386 29236 9392
rect 28908 9376 28960 9382
rect 28908 9318 28960 9324
rect 29000 9376 29052 9382
rect 29000 9318 29052 9324
rect 29026 9276 29334 9285
rect 29026 9274 29032 9276
rect 29088 9274 29112 9276
rect 29168 9274 29192 9276
rect 29248 9274 29272 9276
rect 29328 9274 29334 9276
rect 29088 9222 29090 9274
rect 29270 9222 29272 9274
rect 29026 9220 29032 9222
rect 29088 9220 29112 9222
rect 29168 9220 29192 9222
rect 29248 9220 29272 9222
rect 29328 9220 29334 9222
rect 29026 9211 29334 9220
rect 29380 8974 29408 9998
rect 29472 9722 29500 10746
rect 29552 10600 29604 10606
rect 29552 10542 29604 10548
rect 29564 10266 29592 10542
rect 29644 10532 29696 10538
rect 29644 10474 29696 10480
rect 29552 10260 29604 10266
rect 29552 10202 29604 10208
rect 29656 10062 29684 10474
rect 29748 10470 29776 11154
rect 29736 10464 29788 10470
rect 29736 10406 29788 10412
rect 29644 10056 29696 10062
rect 29644 9998 29696 10004
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29644 9716 29696 9722
rect 29644 9658 29696 9664
rect 29472 9110 29500 9658
rect 29552 9512 29604 9518
rect 29552 9454 29604 9460
rect 29564 9178 29592 9454
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29460 9104 29512 9110
rect 29460 9046 29512 9052
rect 28908 8968 28960 8974
rect 28908 8910 28960 8916
rect 29368 8968 29420 8974
rect 29368 8910 29420 8916
rect 28816 8628 28868 8634
rect 28816 8570 28868 8576
rect 28080 8424 28132 8430
rect 28080 8366 28132 8372
rect 28448 8424 28500 8430
rect 28448 8366 28500 8372
rect 28724 8424 28776 8430
rect 28724 8366 28776 8372
rect 28092 8090 28120 8366
rect 28264 8288 28316 8294
rect 28264 8230 28316 8236
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28816 8288 28868 8294
rect 28920 8242 28948 8910
rect 29276 8832 29328 8838
rect 29276 8774 29328 8780
rect 29288 8430 29316 8774
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 28868 8236 28948 8242
rect 28816 8230 28948 8236
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 28170 7984 28226 7993
rect 28170 7919 28172 7928
rect 28224 7919 28226 7928
rect 28172 7890 28224 7896
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 27620 6316 27672 6322
rect 27620 6258 27672 6264
rect 27252 6180 27304 6186
rect 27252 6122 27304 6128
rect 27632 4146 27660 6258
rect 27712 6180 27764 6186
rect 27712 6122 27764 6128
rect 27724 5914 27752 6122
rect 27712 5908 27764 5914
rect 27712 5850 27764 5856
rect 28184 5778 28212 7890
rect 28276 7426 28304 8230
rect 28736 8090 28764 8230
rect 28828 8214 28948 8230
rect 28724 8084 28776 8090
rect 28724 8026 28776 8032
rect 28724 7744 28776 7750
rect 28724 7686 28776 7692
rect 28366 7644 28674 7653
rect 28366 7642 28372 7644
rect 28428 7642 28452 7644
rect 28508 7642 28532 7644
rect 28588 7642 28612 7644
rect 28668 7642 28674 7644
rect 28428 7590 28430 7642
rect 28610 7590 28612 7642
rect 28366 7588 28372 7590
rect 28428 7588 28452 7590
rect 28508 7588 28532 7590
rect 28588 7588 28612 7590
rect 28668 7588 28674 7590
rect 28366 7579 28674 7588
rect 28736 7546 28764 7686
rect 28920 7546 28948 8214
rect 29026 8188 29334 8197
rect 29026 8186 29032 8188
rect 29088 8186 29112 8188
rect 29168 8186 29192 8188
rect 29248 8186 29272 8188
rect 29328 8186 29334 8188
rect 29088 8134 29090 8186
rect 29270 8134 29272 8186
rect 29026 8132 29032 8134
rect 29088 8132 29112 8134
rect 29168 8132 29192 8134
rect 29248 8132 29272 8134
rect 29328 8132 29334 8134
rect 29026 8123 29334 8132
rect 28724 7540 28776 7546
rect 28724 7482 28776 7488
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 28276 7398 28764 7426
rect 29380 7410 29408 8910
rect 29460 8900 29512 8906
rect 29460 8842 29512 8848
rect 29472 8430 29500 8842
rect 29656 8838 29684 9658
rect 29644 8832 29696 8838
rect 29644 8774 29696 8780
rect 29656 8566 29684 8774
rect 29748 8634 29776 10406
rect 29840 10146 29868 12038
rect 29920 10464 29972 10470
rect 29920 10406 29972 10412
rect 29932 10266 29960 10406
rect 29920 10260 29972 10266
rect 29920 10202 29972 10208
rect 29840 10118 29960 10146
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29644 8560 29696 8566
rect 29644 8502 29696 8508
rect 29460 8424 29512 8430
rect 29460 8366 29512 8372
rect 29828 8424 29880 8430
rect 29828 8366 29880 8372
rect 29644 8356 29696 8362
rect 29644 8298 29696 8304
rect 29460 8288 29512 8294
rect 29460 8230 29512 8236
rect 29472 8022 29500 8230
rect 29460 8016 29512 8022
rect 29460 7958 29512 7964
rect 29458 7848 29514 7857
rect 29458 7783 29514 7792
rect 29472 7750 29500 7783
rect 29656 7750 29684 8298
rect 29736 7948 29788 7954
rect 29736 7890 29788 7896
rect 29460 7744 29512 7750
rect 29460 7686 29512 7692
rect 29644 7744 29696 7750
rect 29644 7686 29696 7692
rect 28264 7336 28316 7342
rect 28264 7278 28316 7284
rect 28448 7336 28500 7342
rect 28448 7278 28500 7284
rect 28276 6866 28304 7278
rect 28460 7018 28488 7278
rect 28736 7274 28764 7398
rect 29368 7404 29420 7410
rect 29368 7346 29420 7352
rect 29000 7336 29052 7342
rect 28920 7284 29000 7290
rect 28920 7278 29052 7284
rect 28724 7268 28776 7274
rect 28724 7210 28776 7216
rect 28920 7262 29040 7278
rect 28368 7002 28488 7018
rect 28736 7002 28764 7210
rect 28356 6996 28488 7002
rect 28408 6990 28488 6996
rect 28724 6996 28776 7002
rect 28356 6938 28408 6944
rect 28724 6938 28776 6944
rect 28264 6860 28316 6866
rect 28264 6802 28316 6808
rect 28276 6458 28304 6802
rect 28736 6798 28764 6938
rect 28724 6792 28776 6798
rect 28724 6734 28776 6740
rect 28816 6656 28868 6662
rect 28816 6598 28868 6604
rect 28366 6556 28674 6565
rect 28366 6554 28372 6556
rect 28428 6554 28452 6556
rect 28508 6554 28532 6556
rect 28588 6554 28612 6556
rect 28668 6554 28674 6556
rect 28428 6502 28430 6554
rect 28610 6502 28612 6554
rect 28366 6500 28372 6502
rect 28428 6500 28452 6502
rect 28508 6500 28532 6502
rect 28588 6500 28612 6502
rect 28668 6500 28674 6502
rect 28366 6491 28674 6500
rect 28264 6452 28316 6458
rect 28264 6394 28316 6400
rect 28828 5914 28856 6598
rect 28920 6322 28948 7262
rect 29748 7206 29776 7890
rect 29368 7200 29420 7206
rect 29368 7142 29420 7148
rect 29736 7200 29788 7206
rect 29736 7142 29788 7148
rect 29026 7100 29334 7109
rect 29026 7098 29032 7100
rect 29088 7098 29112 7100
rect 29168 7098 29192 7100
rect 29248 7098 29272 7100
rect 29328 7098 29334 7100
rect 29088 7046 29090 7098
rect 29270 7046 29272 7098
rect 29026 7044 29032 7046
rect 29088 7044 29112 7046
rect 29168 7044 29192 7046
rect 29248 7044 29272 7046
rect 29328 7044 29334 7046
rect 29026 7035 29334 7044
rect 28908 6316 28960 6322
rect 28908 6258 28960 6264
rect 29026 6012 29334 6021
rect 29026 6010 29032 6012
rect 29088 6010 29112 6012
rect 29168 6010 29192 6012
rect 29248 6010 29272 6012
rect 29328 6010 29334 6012
rect 29088 5958 29090 6010
rect 29270 5958 29272 6010
rect 29026 5956 29032 5958
rect 29088 5956 29112 5958
rect 29168 5956 29192 5958
rect 29248 5956 29272 5958
rect 29328 5956 29334 5958
rect 29026 5947 29334 5956
rect 28816 5908 28868 5914
rect 28816 5850 28868 5856
rect 28172 5772 28224 5778
rect 28172 5714 28224 5720
rect 28724 5772 28776 5778
rect 28724 5714 28776 5720
rect 27620 4140 27672 4146
rect 27620 4082 27672 4088
rect 28184 3942 28212 5714
rect 28736 5574 28764 5714
rect 29380 5710 29408 7142
rect 29840 6798 29868 8366
rect 29932 8090 29960 10118
rect 29920 8084 29972 8090
rect 29920 8026 29972 8032
rect 29828 6792 29880 6798
rect 29828 6734 29880 6740
rect 29840 6390 29868 6734
rect 29828 6384 29880 6390
rect 29828 6326 29880 6332
rect 29552 6180 29604 6186
rect 29552 6122 29604 6128
rect 29460 6112 29512 6118
rect 29460 6054 29512 6060
rect 29472 5778 29500 6054
rect 29564 5914 29592 6122
rect 29552 5908 29604 5914
rect 29552 5850 29604 5856
rect 29460 5772 29512 5778
rect 29460 5714 29512 5720
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 29734 5672 29790 5681
rect 29734 5607 29790 5616
rect 28724 5568 28776 5574
rect 28724 5510 28776 5516
rect 28366 5468 28674 5477
rect 28366 5466 28372 5468
rect 28428 5466 28452 5468
rect 28508 5466 28532 5468
rect 28588 5466 28612 5468
rect 28668 5466 28674 5468
rect 28428 5414 28430 5466
rect 28610 5414 28612 5466
rect 28366 5412 28372 5414
rect 28428 5412 28452 5414
rect 28508 5412 28532 5414
rect 28588 5412 28612 5414
rect 28668 5412 28674 5414
rect 28366 5403 28674 5412
rect 28540 5024 28592 5030
rect 28540 4966 28592 4972
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 28552 4690 28580 4966
rect 29026 4924 29334 4933
rect 29026 4922 29032 4924
rect 29088 4922 29112 4924
rect 29168 4922 29192 4924
rect 29248 4922 29272 4924
rect 29328 4922 29334 4924
rect 29088 4870 29090 4922
rect 29270 4870 29272 4922
rect 29026 4868 29032 4870
rect 29088 4868 29112 4870
rect 29168 4868 29192 4870
rect 29248 4868 29272 4870
rect 29328 4868 29334 4870
rect 29026 4859 29334 4868
rect 29472 4826 29500 4966
rect 29748 4826 29776 5607
rect 29932 5574 29960 8026
rect 30024 6322 30052 13654
rect 30116 12850 30144 13790
rect 30104 12844 30156 12850
rect 30104 12786 30156 12792
rect 30116 12374 30144 12786
rect 30104 12368 30156 12374
rect 30104 12310 30156 12316
rect 30208 12306 30236 14010
rect 30288 13728 30340 13734
rect 30288 13670 30340 13676
rect 30196 12300 30248 12306
rect 30196 12242 30248 12248
rect 30208 11558 30236 12242
rect 30300 11830 30328 13670
rect 30564 13456 30616 13462
rect 30562 13424 30564 13433
rect 30616 13424 30618 13433
rect 30562 13359 30618 13368
rect 30668 12986 30696 14418
rect 30748 14272 30800 14278
rect 30748 14214 30800 14220
rect 30760 14074 30788 14214
rect 30748 14068 30800 14074
rect 30748 14010 30800 14016
rect 30852 13954 30880 14418
rect 30760 13926 30880 13954
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30656 12640 30708 12646
rect 30484 12588 30656 12594
rect 30484 12582 30708 12588
rect 30484 12566 30696 12582
rect 30288 11824 30340 11830
rect 30288 11766 30340 11772
rect 30484 11626 30512 12566
rect 30472 11620 30524 11626
rect 30472 11562 30524 11568
rect 30196 11552 30248 11558
rect 30196 11494 30248 11500
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30104 11212 30156 11218
rect 30104 11154 30156 11160
rect 30116 10810 30144 11154
rect 30208 10810 30236 11494
rect 30392 11354 30420 11494
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30288 11212 30340 11218
rect 30288 11154 30340 11160
rect 30300 10810 30328 11154
rect 30104 10804 30156 10810
rect 30104 10746 30156 10752
rect 30196 10804 30248 10810
rect 30196 10746 30248 10752
rect 30288 10804 30340 10810
rect 30288 10746 30340 10752
rect 30208 10062 30236 10746
rect 30300 10538 30328 10746
rect 30288 10532 30340 10538
rect 30288 10474 30340 10480
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 30300 9450 30328 10474
rect 30484 9586 30512 11562
rect 30760 11354 30788 13926
rect 30840 13796 30892 13802
rect 30840 13738 30892 13744
rect 30852 13326 30880 13738
rect 30944 13530 30972 15030
rect 31404 14804 31432 19722
rect 31588 17218 31616 24142
rect 33152 23905 33180 24142
rect 33138 23896 33194 23905
rect 33138 23831 33194 23840
rect 31666 22536 31722 22545
rect 31666 22471 31722 22480
rect 31680 22098 31708 22471
rect 31668 22092 31720 22098
rect 31668 22034 31720 22040
rect 33048 20936 33100 20942
rect 33048 20878 33100 20884
rect 33060 20505 33088 20878
rect 33046 20496 33102 20505
rect 33046 20431 33102 20440
rect 33138 19136 33194 19145
rect 33138 19071 33194 19080
rect 33152 18902 33180 19071
rect 33140 18896 33192 18902
rect 33140 18838 33192 18844
rect 33140 17672 33192 17678
rect 33140 17614 33192 17620
rect 31128 14776 31432 14804
rect 31496 17190 31616 17218
rect 31024 14408 31076 14414
rect 31024 14350 31076 14356
rect 31036 14074 31064 14350
rect 31024 14068 31076 14074
rect 31024 14010 31076 14016
rect 31022 13832 31078 13841
rect 31022 13767 31078 13776
rect 30932 13524 30984 13530
rect 30932 13466 30984 13472
rect 31036 13462 31064 13767
rect 31024 13456 31076 13462
rect 31024 13398 31076 13404
rect 30840 13320 30892 13326
rect 30840 13262 30892 13268
rect 30932 13320 30984 13326
rect 30932 13262 30984 13268
rect 30944 11898 30972 13262
rect 31128 12434 31156 14776
rect 31300 14408 31352 14414
rect 31300 14350 31352 14356
rect 31128 12406 31248 12434
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 30840 11824 30892 11830
rect 30840 11766 30892 11772
rect 30852 11354 30880 11766
rect 30748 11348 30800 11354
rect 30748 11290 30800 11296
rect 30840 11348 30892 11354
rect 30840 11290 30892 11296
rect 30760 10606 30788 11290
rect 31024 11008 31076 11014
rect 31024 10950 31076 10956
rect 30748 10600 30800 10606
rect 30748 10542 30800 10548
rect 30932 10600 30984 10606
rect 30932 10542 30984 10548
rect 30944 10266 30972 10542
rect 30932 10260 30984 10266
rect 30932 10202 30984 10208
rect 30472 9580 30524 9586
rect 30472 9522 30524 9528
rect 30380 9512 30432 9518
rect 30380 9454 30432 9460
rect 30656 9512 30708 9518
rect 30656 9454 30708 9460
rect 30288 9444 30340 9450
rect 30288 9386 30340 9392
rect 30104 9376 30156 9382
rect 30104 9318 30156 9324
rect 30116 9178 30144 9318
rect 30104 9172 30156 9178
rect 30104 9114 30156 9120
rect 30288 8832 30340 8838
rect 30288 8774 30340 8780
rect 30300 8430 30328 8774
rect 30288 8424 30340 8430
rect 30288 8366 30340 8372
rect 30392 8022 30420 9454
rect 30668 8634 30696 9454
rect 30656 8628 30708 8634
rect 30656 8570 30708 8576
rect 30656 8424 30708 8430
rect 30484 8384 30656 8412
rect 30484 8294 30512 8384
rect 30840 8424 30892 8430
rect 30656 8366 30708 8372
rect 30760 8384 30840 8412
rect 30472 8288 30524 8294
rect 30472 8230 30524 8236
rect 30564 8288 30616 8294
rect 30564 8230 30616 8236
rect 30576 8090 30604 8230
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 30380 8016 30432 8022
rect 30380 7958 30432 7964
rect 30760 7954 30788 8384
rect 30840 8366 30892 8372
rect 30748 7948 30800 7954
rect 30748 7890 30800 7896
rect 30840 7948 30892 7954
rect 30840 7890 30892 7896
rect 30104 7744 30156 7750
rect 30104 7686 30156 7692
rect 30116 7546 30144 7686
rect 30852 7546 30880 7890
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 30840 7540 30892 7546
rect 30840 7482 30892 7488
rect 30472 7336 30524 7342
rect 30472 7278 30524 7284
rect 30104 6656 30156 6662
rect 30104 6598 30156 6604
rect 30116 6458 30144 6598
rect 30484 6458 30512 7278
rect 30656 6792 30708 6798
rect 30656 6734 30708 6740
rect 30104 6452 30156 6458
rect 30104 6394 30156 6400
rect 30472 6452 30524 6458
rect 30472 6394 30524 6400
rect 30012 6316 30064 6322
rect 30012 6258 30064 6264
rect 30668 5914 30696 6734
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 29920 5568 29972 5574
rect 29920 5510 29972 5516
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29736 4820 29788 4826
rect 29736 4762 29788 4768
rect 28540 4684 28592 4690
rect 28540 4626 28592 4632
rect 28264 4480 28316 4486
rect 28264 4422 28316 4428
rect 28276 4010 28304 4422
rect 28366 4380 28674 4389
rect 28366 4378 28372 4380
rect 28428 4378 28452 4380
rect 28508 4378 28532 4380
rect 28588 4378 28612 4380
rect 28668 4378 28674 4380
rect 28428 4326 28430 4378
rect 28610 4326 28612 4378
rect 28366 4324 28372 4326
rect 28428 4324 28452 4326
rect 28508 4324 28532 4326
rect 28588 4324 28612 4326
rect 28668 4324 28674 4326
rect 28366 4315 28674 4324
rect 30024 4282 30052 5102
rect 31036 4706 31064 10950
rect 31220 9602 31248 12406
rect 31312 11354 31340 14350
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31496 11234 31524 17190
rect 33152 17105 33180 17614
rect 33138 17096 33194 17105
rect 33138 17031 33194 17040
rect 31852 16584 31904 16590
rect 31852 16526 31904 16532
rect 31864 16250 31892 16526
rect 31852 16244 31904 16250
rect 31852 16186 31904 16192
rect 33138 15736 33194 15745
rect 33138 15671 33194 15680
rect 33152 15638 33180 15671
rect 33140 15632 33192 15638
rect 33140 15574 33192 15580
rect 31668 14884 31720 14890
rect 31668 14826 31720 14832
rect 31576 13796 31628 13802
rect 31576 13738 31628 13744
rect 31588 11354 31616 13738
rect 31680 13394 31708 14826
rect 33140 14408 33192 14414
rect 33138 14376 33140 14385
rect 33192 14376 33194 14385
rect 33138 14311 33194 14320
rect 31760 13864 31812 13870
rect 31760 13806 31812 13812
rect 31772 13530 31800 13806
rect 31760 13524 31812 13530
rect 31760 13466 31812 13472
rect 31758 13424 31814 13433
rect 31668 13388 31720 13394
rect 31758 13359 31814 13368
rect 31668 13330 31720 13336
rect 31576 11348 31628 11354
rect 31576 11290 31628 11296
rect 31392 11212 31444 11218
rect 31496 11206 31616 11234
rect 31680 11218 31708 13330
rect 31772 13326 31800 13359
rect 31760 13320 31812 13326
rect 31760 13262 31812 13268
rect 31760 13184 31812 13190
rect 31760 13126 31812 13132
rect 31772 11762 31800 13126
rect 33138 12336 33194 12345
rect 33138 12271 33140 12280
rect 33192 12271 33194 12280
rect 33140 12242 33192 12248
rect 31760 11756 31812 11762
rect 31760 11698 31812 11704
rect 31392 11154 31444 11160
rect 31404 10985 31432 11154
rect 31484 11076 31536 11082
rect 31484 11018 31536 11024
rect 31390 10976 31446 10985
rect 31390 10911 31446 10920
rect 31392 10532 31444 10538
rect 31392 10474 31444 10480
rect 31404 10130 31432 10474
rect 31496 10130 31524 11018
rect 31392 10124 31444 10130
rect 31392 10066 31444 10072
rect 31484 10124 31536 10130
rect 31484 10066 31536 10072
rect 31220 9574 31340 9602
rect 31208 9512 31260 9518
rect 31208 9454 31260 9460
rect 31220 9178 31248 9454
rect 31208 9172 31260 9178
rect 31208 9114 31260 9120
rect 31116 9104 31168 9110
rect 31116 9046 31168 9052
rect 31128 8634 31156 9046
rect 31116 8628 31168 8634
rect 31116 8570 31168 8576
rect 31116 8424 31168 8430
rect 31116 8366 31168 8372
rect 31208 8424 31260 8430
rect 31208 8366 31260 8372
rect 31128 8090 31156 8366
rect 31116 8084 31168 8090
rect 31116 8026 31168 8032
rect 31220 6254 31248 8366
rect 31208 6248 31260 6254
rect 31208 6190 31260 6196
rect 30852 4690 31064 4706
rect 30840 4684 31064 4690
rect 30892 4678 31064 4684
rect 30840 4626 30892 4632
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30932 4616 30984 4622
rect 30932 4558 30984 4564
rect 30012 4276 30064 4282
rect 30012 4218 30064 4224
rect 28264 4004 28316 4010
rect 28264 3946 28316 3952
rect 28172 3936 28224 3942
rect 28172 3878 28224 3884
rect 29026 3836 29334 3845
rect 29026 3834 29032 3836
rect 29088 3834 29112 3836
rect 29168 3834 29192 3836
rect 29248 3834 29272 3836
rect 29328 3834 29334 3836
rect 29088 3782 29090 3834
rect 29270 3782 29272 3834
rect 29026 3780 29032 3782
rect 29088 3780 29112 3782
rect 29168 3780 29192 3782
rect 29248 3780 29272 3782
rect 29328 3780 29334 3782
rect 29026 3771 29334 3780
rect 30024 3602 30052 4218
rect 30484 4214 30512 4558
rect 30472 4208 30524 4214
rect 30472 4150 30524 4156
rect 25780 3596 25832 3602
rect 25780 3538 25832 3544
rect 30012 3596 30064 3602
rect 30012 3538 30064 3544
rect 24492 3528 24544 3534
rect 24492 3470 24544 3476
rect 30288 3528 30340 3534
rect 30288 3470 30340 3476
rect 23480 2984 23532 2990
rect 23480 2926 23532 2932
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 24504 800 24532 3470
rect 28366 3292 28674 3301
rect 28366 3290 28372 3292
rect 28428 3290 28452 3292
rect 28508 3290 28532 3292
rect 28588 3290 28612 3292
rect 28668 3290 28674 3292
rect 28428 3238 28430 3290
rect 28610 3238 28612 3290
rect 28366 3236 28372 3238
rect 28428 3236 28452 3238
rect 28508 3236 28532 3238
rect 28588 3236 28612 3238
rect 28668 3236 28674 3238
rect 28366 3227 28674 3236
rect 25780 3052 25832 3058
rect 25780 2994 25832 3000
rect 25792 800 25820 2994
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 29368 2984 29420 2990
rect 29368 2926 29420 2932
rect 27080 800 27108 2926
rect 29026 2748 29334 2757
rect 29026 2746 29032 2748
rect 29088 2746 29112 2748
rect 29168 2746 29192 2748
rect 29248 2746 29272 2748
rect 29328 2746 29334 2748
rect 29088 2694 29090 2746
rect 29270 2694 29272 2746
rect 29026 2692 29032 2694
rect 29088 2692 29112 2694
rect 29168 2692 29192 2694
rect 29248 2692 29272 2694
rect 29328 2692 29334 2694
rect 29026 2683 29334 2692
rect 29012 870 29132 898
rect 29012 800 29040 870
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28998 0 29054 800
rect 29104 762 29132 870
rect 29380 762 29408 2926
rect 30300 800 30328 3470
rect 30944 3194 30972 4558
rect 31312 3942 31340 9574
rect 31404 8430 31432 10066
rect 31484 8832 31536 8838
rect 31484 8774 31536 8780
rect 31496 8430 31524 8774
rect 31392 8424 31444 8430
rect 31392 8366 31444 8372
rect 31484 8424 31536 8430
rect 31484 8366 31536 8372
rect 31588 7857 31616 11206
rect 31668 11212 31720 11218
rect 31668 11154 31720 11160
rect 33138 9616 33194 9625
rect 33138 9551 33194 9560
rect 33152 9110 33180 9551
rect 33140 9104 33192 9110
rect 31666 9072 31722 9081
rect 33140 9046 33192 9052
rect 31666 9007 31722 9016
rect 31680 8906 31708 9007
rect 31668 8900 31720 8906
rect 31668 8842 31720 8848
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 31574 7848 31630 7857
rect 31574 7783 31630 7792
rect 31668 7744 31720 7750
rect 31668 7686 31720 7692
rect 31680 5273 31708 7686
rect 33152 7585 33180 7890
rect 33138 7576 33194 7585
rect 33138 7511 33194 7520
rect 33140 6248 33192 6254
rect 33138 6216 33140 6225
rect 33192 6216 33194 6225
rect 33138 6151 33194 6160
rect 31666 5264 31722 5273
rect 31666 5199 31722 5208
rect 31668 4616 31720 4622
rect 31668 4558 31720 4564
rect 31852 4616 31904 4622
rect 31852 4558 31904 4564
rect 31680 4282 31708 4558
rect 31668 4276 31720 4282
rect 31668 4218 31720 4224
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31668 3664 31720 3670
rect 31668 3606 31720 3612
rect 30932 3188 30984 3194
rect 30932 3130 30984 3136
rect 31680 1465 31708 3606
rect 31864 3194 31892 4558
rect 33046 4176 33102 4185
rect 33046 4111 33048 4120
rect 33100 4111 33102 4120
rect 33048 4082 33100 4088
rect 33508 4004 33560 4010
rect 33508 3946 33560 3952
rect 31852 3188 31904 3194
rect 31852 3130 31904 3136
rect 32220 3052 32272 3058
rect 32220 2994 32272 3000
rect 31666 1456 31722 1465
rect 31666 1391 31722 1400
rect 32232 800 32260 2994
rect 33140 2916 33192 2922
rect 33140 2858 33192 2864
rect 33152 2825 33180 2858
rect 33138 2816 33194 2825
rect 33138 2751 33194 2760
rect 33520 800 33548 3946
rect 34796 2848 34848 2854
rect 34796 2790 34848 2796
rect 34808 800 34836 2790
rect 29104 734 29408 762
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 33506 0 33562 800
rect 34794 0 34850 800
<< via2 >>
rect 4526 34040 4582 34096
rect 2778 32000 2834 32056
rect 1306 30676 1308 30696
rect 1308 30676 1360 30696
rect 1360 30676 1362 30696
rect 1306 30640 1362 30676
rect 1306 27240 1362 27296
rect 1306 23840 1362 23896
rect 1306 22500 1362 22536
rect 1306 22480 1308 22500
rect 1308 22480 1360 22500
rect 1360 22480 1362 22500
rect 3514 28600 3570 28656
rect 3238 25880 3294 25936
rect 6952 32122 7008 32124
rect 7032 32122 7088 32124
rect 7112 32122 7168 32124
rect 7192 32122 7248 32124
rect 6952 32070 6998 32122
rect 6998 32070 7008 32122
rect 7032 32070 7062 32122
rect 7062 32070 7074 32122
rect 7074 32070 7088 32122
rect 7112 32070 7126 32122
rect 7126 32070 7138 32122
rect 7138 32070 7168 32122
rect 7192 32070 7202 32122
rect 7202 32070 7248 32122
rect 6952 32068 7008 32070
rect 7032 32068 7088 32070
rect 7112 32068 7168 32070
rect 7192 32068 7248 32070
rect 6292 31578 6348 31580
rect 6372 31578 6428 31580
rect 6452 31578 6508 31580
rect 6532 31578 6588 31580
rect 6292 31526 6338 31578
rect 6338 31526 6348 31578
rect 6372 31526 6402 31578
rect 6402 31526 6414 31578
rect 6414 31526 6428 31578
rect 6452 31526 6466 31578
rect 6466 31526 6478 31578
rect 6478 31526 6508 31578
rect 6532 31526 6542 31578
rect 6542 31526 6588 31578
rect 6292 31524 6348 31526
rect 6372 31524 6428 31526
rect 6452 31524 6508 31526
rect 6532 31524 6588 31526
rect 3330 21004 3386 21040
rect 3330 20984 3332 21004
rect 3332 20984 3384 21004
rect 3384 20984 3386 21004
rect 3054 20440 3110 20496
rect 1306 19080 1362 19136
rect 1306 15680 1362 15736
rect 1306 14320 1362 14376
rect 1306 12960 1362 13016
rect 4066 17720 4122 17776
rect 3238 10920 3294 10976
rect 3054 9560 3110 9616
rect 1306 7520 1362 7576
rect 1306 6196 1308 6216
rect 1308 6196 1360 6216
rect 1360 6196 1362 6216
rect 1306 6160 1362 6196
rect 1306 4800 1362 4856
rect 6292 30490 6348 30492
rect 6372 30490 6428 30492
rect 6452 30490 6508 30492
rect 6532 30490 6588 30492
rect 6292 30438 6338 30490
rect 6338 30438 6348 30490
rect 6372 30438 6402 30490
rect 6402 30438 6414 30490
rect 6414 30438 6428 30490
rect 6452 30438 6466 30490
rect 6466 30438 6478 30490
rect 6478 30438 6508 30490
rect 6532 30438 6542 30490
rect 6542 30438 6588 30490
rect 6292 30436 6348 30438
rect 6372 30436 6428 30438
rect 6452 30436 6508 30438
rect 6532 30436 6588 30438
rect 6292 29402 6348 29404
rect 6372 29402 6428 29404
rect 6452 29402 6508 29404
rect 6532 29402 6588 29404
rect 6292 29350 6338 29402
rect 6338 29350 6348 29402
rect 6372 29350 6402 29402
rect 6402 29350 6414 29402
rect 6414 29350 6428 29402
rect 6452 29350 6466 29402
rect 6466 29350 6478 29402
rect 6478 29350 6508 29402
rect 6532 29350 6542 29402
rect 6542 29350 6588 29402
rect 6292 29348 6348 29350
rect 6372 29348 6428 29350
rect 6452 29348 6508 29350
rect 6532 29348 6588 29350
rect 6952 31034 7008 31036
rect 7032 31034 7088 31036
rect 7112 31034 7168 31036
rect 7192 31034 7248 31036
rect 6952 30982 6998 31034
rect 6998 30982 7008 31034
rect 7032 30982 7062 31034
rect 7062 30982 7074 31034
rect 7074 30982 7088 31034
rect 7112 30982 7126 31034
rect 7126 30982 7138 31034
rect 7138 30982 7168 31034
rect 7192 30982 7202 31034
rect 7202 30982 7248 31034
rect 6952 30980 7008 30982
rect 7032 30980 7088 30982
rect 7112 30980 7168 30982
rect 7192 30980 7248 30982
rect 6952 29946 7008 29948
rect 7032 29946 7088 29948
rect 7112 29946 7168 29948
rect 7192 29946 7248 29948
rect 6952 29894 6998 29946
rect 6998 29894 7008 29946
rect 7032 29894 7062 29946
rect 7062 29894 7074 29946
rect 7074 29894 7088 29946
rect 7112 29894 7126 29946
rect 7126 29894 7138 29946
rect 7138 29894 7168 29946
rect 7192 29894 7202 29946
rect 7202 29894 7248 29946
rect 6952 29892 7008 29894
rect 7032 29892 7088 29894
rect 7112 29892 7168 29894
rect 7192 29892 7248 29894
rect 6292 28314 6348 28316
rect 6372 28314 6428 28316
rect 6452 28314 6508 28316
rect 6532 28314 6588 28316
rect 6292 28262 6338 28314
rect 6338 28262 6348 28314
rect 6372 28262 6402 28314
rect 6402 28262 6414 28314
rect 6414 28262 6428 28314
rect 6452 28262 6466 28314
rect 6466 28262 6478 28314
rect 6478 28262 6508 28314
rect 6532 28262 6542 28314
rect 6542 28262 6588 28314
rect 6292 28260 6348 28262
rect 6372 28260 6428 28262
rect 6452 28260 6508 28262
rect 6532 28260 6588 28262
rect 6952 28858 7008 28860
rect 7032 28858 7088 28860
rect 7112 28858 7168 28860
rect 7192 28858 7248 28860
rect 6952 28806 6998 28858
rect 6998 28806 7008 28858
rect 7032 28806 7062 28858
rect 7062 28806 7074 28858
rect 7074 28806 7088 28858
rect 7112 28806 7126 28858
rect 7126 28806 7138 28858
rect 7138 28806 7168 28858
rect 7192 28806 7202 28858
rect 7202 28806 7248 28858
rect 6952 28804 7008 28806
rect 7032 28804 7088 28806
rect 7112 28804 7168 28806
rect 7192 28804 7248 28806
rect 6952 27770 7008 27772
rect 7032 27770 7088 27772
rect 7112 27770 7168 27772
rect 7192 27770 7248 27772
rect 6952 27718 6998 27770
rect 6998 27718 7008 27770
rect 7032 27718 7062 27770
rect 7062 27718 7074 27770
rect 7074 27718 7088 27770
rect 7112 27718 7126 27770
rect 7126 27718 7138 27770
rect 7138 27718 7168 27770
rect 7192 27718 7202 27770
rect 7202 27718 7248 27770
rect 6952 27716 7008 27718
rect 7032 27716 7088 27718
rect 7112 27716 7168 27718
rect 7192 27716 7248 27718
rect 6826 27532 6882 27568
rect 6826 27512 6828 27532
rect 6828 27512 6880 27532
rect 6880 27512 6882 27532
rect 6292 27226 6348 27228
rect 6372 27226 6428 27228
rect 6452 27226 6508 27228
rect 6532 27226 6588 27228
rect 6292 27174 6338 27226
rect 6338 27174 6348 27226
rect 6372 27174 6402 27226
rect 6402 27174 6414 27226
rect 6414 27174 6428 27226
rect 6452 27174 6466 27226
rect 6466 27174 6478 27226
rect 6478 27174 6508 27226
rect 6532 27174 6542 27226
rect 6542 27174 6588 27226
rect 6292 27172 6348 27174
rect 6372 27172 6428 27174
rect 6452 27172 6508 27174
rect 6532 27172 6588 27174
rect 6952 26682 7008 26684
rect 7032 26682 7088 26684
rect 7112 26682 7168 26684
rect 7192 26682 7248 26684
rect 6952 26630 6998 26682
rect 6998 26630 7008 26682
rect 7032 26630 7062 26682
rect 7062 26630 7074 26682
rect 7074 26630 7088 26682
rect 7112 26630 7126 26682
rect 7126 26630 7138 26682
rect 7138 26630 7168 26682
rect 7192 26630 7202 26682
rect 7202 26630 7248 26682
rect 6952 26628 7008 26630
rect 7032 26628 7088 26630
rect 7112 26628 7168 26630
rect 7192 26628 7248 26630
rect 6292 26138 6348 26140
rect 6372 26138 6428 26140
rect 6452 26138 6508 26140
rect 6532 26138 6588 26140
rect 6292 26086 6338 26138
rect 6338 26086 6348 26138
rect 6372 26086 6402 26138
rect 6402 26086 6414 26138
rect 6414 26086 6428 26138
rect 6452 26086 6466 26138
rect 6466 26086 6478 26138
rect 6478 26086 6508 26138
rect 6532 26086 6542 26138
rect 6542 26086 6588 26138
rect 6292 26084 6348 26086
rect 6372 26084 6428 26086
rect 6452 26084 6508 26086
rect 6532 26084 6588 26086
rect 6952 25594 7008 25596
rect 7032 25594 7088 25596
rect 7112 25594 7168 25596
rect 7192 25594 7248 25596
rect 6952 25542 6998 25594
rect 6998 25542 7008 25594
rect 7032 25542 7062 25594
rect 7062 25542 7074 25594
rect 7074 25542 7088 25594
rect 7112 25542 7126 25594
rect 7126 25542 7138 25594
rect 7138 25542 7168 25594
rect 7192 25542 7202 25594
rect 7202 25542 7248 25594
rect 6952 25540 7008 25542
rect 7032 25540 7088 25542
rect 7112 25540 7168 25542
rect 7192 25540 7248 25542
rect 6292 25050 6348 25052
rect 6372 25050 6428 25052
rect 6452 25050 6508 25052
rect 6532 25050 6588 25052
rect 6292 24998 6338 25050
rect 6338 24998 6348 25050
rect 6372 24998 6402 25050
rect 6402 24998 6414 25050
rect 6414 24998 6428 25050
rect 6452 24998 6466 25050
rect 6466 24998 6478 25050
rect 6478 24998 6508 25050
rect 6532 24998 6542 25050
rect 6542 24998 6588 25050
rect 6292 24996 6348 24998
rect 6372 24996 6428 24998
rect 6452 24996 6508 24998
rect 6532 24996 6588 24998
rect 6952 24506 7008 24508
rect 7032 24506 7088 24508
rect 7112 24506 7168 24508
rect 7192 24506 7248 24508
rect 6952 24454 6998 24506
rect 6998 24454 7008 24506
rect 7032 24454 7062 24506
rect 7062 24454 7074 24506
rect 7074 24454 7088 24506
rect 7112 24454 7126 24506
rect 7126 24454 7138 24506
rect 7138 24454 7168 24506
rect 7192 24454 7202 24506
rect 7202 24454 7248 24506
rect 6952 24452 7008 24454
rect 7032 24452 7088 24454
rect 7112 24452 7168 24454
rect 7192 24452 7248 24454
rect 6292 23962 6348 23964
rect 6372 23962 6428 23964
rect 6452 23962 6508 23964
rect 6532 23962 6588 23964
rect 6292 23910 6338 23962
rect 6338 23910 6348 23962
rect 6372 23910 6402 23962
rect 6402 23910 6414 23962
rect 6414 23910 6428 23962
rect 6452 23910 6466 23962
rect 6466 23910 6478 23962
rect 6478 23910 6508 23962
rect 6532 23910 6542 23962
rect 6542 23910 6588 23962
rect 6292 23908 6348 23910
rect 6372 23908 6428 23910
rect 6452 23908 6508 23910
rect 6532 23908 6588 23910
rect 6952 23418 7008 23420
rect 7032 23418 7088 23420
rect 7112 23418 7168 23420
rect 7192 23418 7248 23420
rect 6952 23366 6998 23418
rect 6998 23366 7008 23418
rect 7032 23366 7062 23418
rect 7062 23366 7074 23418
rect 7074 23366 7088 23418
rect 7112 23366 7126 23418
rect 7126 23366 7138 23418
rect 7138 23366 7168 23418
rect 7192 23366 7202 23418
rect 7202 23366 7248 23418
rect 6952 23364 7008 23366
rect 7032 23364 7088 23366
rect 7112 23364 7168 23366
rect 7192 23364 7248 23366
rect 6292 22874 6348 22876
rect 6372 22874 6428 22876
rect 6452 22874 6508 22876
rect 6532 22874 6588 22876
rect 6292 22822 6338 22874
rect 6338 22822 6348 22874
rect 6372 22822 6402 22874
rect 6402 22822 6414 22874
rect 6414 22822 6428 22874
rect 6452 22822 6466 22874
rect 6466 22822 6478 22874
rect 6478 22822 6508 22874
rect 6532 22822 6542 22874
rect 6542 22822 6588 22874
rect 6292 22820 6348 22822
rect 6372 22820 6428 22822
rect 6452 22820 6508 22822
rect 6532 22820 6588 22822
rect 6292 21786 6348 21788
rect 6372 21786 6428 21788
rect 6452 21786 6508 21788
rect 6532 21786 6588 21788
rect 6292 21734 6338 21786
rect 6338 21734 6348 21786
rect 6372 21734 6402 21786
rect 6402 21734 6414 21786
rect 6414 21734 6428 21786
rect 6452 21734 6466 21786
rect 6466 21734 6478 21786
rect 6478 21734 6508 21786
rect 6532 21734 6542 21786
rect 6542 21734 6588 21786
rect 6292 21732 6348 21734
rect 6372 21732 6428 21734
rect 6452 21732 6508 21734
rect 6532 21732 6588 21734
rect 6292 20698 6348 20700
rect 6372 20698 6428 20700
rect 6452 20698 6508 20700
rect 6532 20698 6588 20700
rect 6292 20646 6338 20698
rect 6338 20646 6348 20698
rect 6372 20646 6402 20698
rect 6402 20646 6414 20698
rect 6414 20646 6428 20698
rect 6452 20646 6466 20698
rect 6466 20646 6478 20698
rect 6478 20646 6508 20698
rect 6532 20646 6542 20698
rect 6542 20646 6588 20698
rect 6292 20644 6348 20646
rect 6372 20644 6428 20646
rect 6452 20644 6508 20646
rect 6532 20644 6588 20646
rect 6292 19610 6348 19612
rect 6372 19610 6428 19612
rect 6452 19610 6508 19612
rect 6532 19610 6588 19612
rect 6292 19558 6338 19610
rect 6338 19558 6348 19610
rect 6372 19558 6402 19610
rect 6402 19558 6414 19610
rect 6414 19558 6428 19610
rect 6452 19558 6466 19610
rect 6466 19558 6478 19610
rect 6478 19558 6508 19610
rect 6532 19558 6542 19610
rect 6542 19558 6588 19610
rect 6292 19556 6348 19558
rect 6372 19556 6428 19558
rect 6452 19556 6508 19558
rect 6532 19556 6588 19558
rect 6292 18522 6348 18524
rect 6372 18522 6428 18524
rect 6452 18522 6508 18524
rect 6532 18522 6588 18524
rect 6292 18470 6338 18522
rect 6338 18470 6348 18522
rect 6372 18470 6402 18522
rect 6402 18470 6414 18522
rect 6414 18470 6428 18522
rect 6452 18470 6466 18522
rect 6466 18470 6478 18522
rect 6478 18470 6508 18522
rect 6532 18470 6542 18522
rect 6542 18470 6588 18522
rect 6292 18468 6348 18470
rect 6372 18468 6428 18470
rect 6452 18468 6508 18470
rect 6532 18468 6588 18470
rect 6292 17434 6348 17436
rect 6372 17434 6428 17436
rect 6452 17434 6508 17436
rect 6532 17434 6588 17436
rect 6292 17382 6338 17434
rect 6338 17382 6348 17434
rect 6372 17382 6402 17434
rect 6402 17382 6414 17434
rect 6414 17382 6428 17434
rect 6452 17382 6466 17434
rect 6466 17382 6478 17434
rect 6478 17382 6508 17434
rect 6532 17382 6542 17434
rect 6542 17382 6588 17434
rect 6292 17380 6348 17382
rect 6372 17380 6428 17382
rect 6452 17380 6508 17382
rect 6532 17380 6588 17382
rect 6292 16346 6348 16348
rect 6372 16346 6428 16348
rect 6452 16346 6508 16348
rect 6532 16346 6588 16348
rect 6292 16294 6338 16346
rect 6338 16294 6348 16346
rect 6372 16294 6402 16346
rect 6402 16294 6414 16346
rect 6414 16294 6428 16346
rect 6452 16294 6466 16346
rect 6466 16294 6478 16346
rect 6478 16294 6508 16346
rect 6532 16294 6542 16346
rect 6542 16294 6588 16346
rect 6292 16292 6348 16294
rect 6372 16292 6428 16294
rect 6452 16292 6508 16294
rect 6532 16292 6588 16294
rect 6952 22330 7008 22332
rect 7032 22330 7088 22332
rect 7112 22330 7168 22332
rect 7192 22330 7248 22332
rect 6952 22278 6998 22330
rect 6998 22278 7008 22330
rect 7032 22278 7062 22330
rect 7062 22278 7074 22330
rect 7074 22278 7088 22330
rect 7112 22278 7126 22330
rect 7126 22278 7138 22330
rect 7138 22278 7168 22330
rect 7192 22278 7202 22330
rect 7202 22278 7248 22330
rect 6952 22276 7008 22278
rect 7032 22276 7088 22278
rect 7112 22276 7168 22278
rect 7192 22276 7248 22278
rect 6952 21242 7008 21244
rect 7032 21242 7088 21244
rect 7112 21242 7168 21244
rect 7192 21242 7248 21244
rect 6952 21190 6998 21242
rect 6998 21190 7008 21242
rect 7032 21190 7062 21242
rect 7062 21190 7074 21242
rect 7074 21190 7088 21242
rect 7112 21190 7126 21242
rect 7126 21190 7138 21242
rect 7138 21190 7168 21242
rect 7192 21190 7202 21242
rect 7202 21190 7248 21242
rect 6952 21188 7008 21190
rect 7032 21188 7088 21190
rect 7112 21188 7168 21190
rect 7192 21188 7248 21190
rect 6952 20154 7008 20156
rect 7032 20154 7088 20156
rect 7112 20154 7168 20156
rect 7192 20154 7248 20156
rect 6952 20102 6998 20154
rect 6998 20102 7008 20154
rect 7032 20102 7062 20154
rect 7062 20102 7074 20154
rect 7074 20102 7088 20154
rect 7112 20102 7126 20154
rect 7126 20102 7138 20154
rect 7138 20102 7168 20154
rect 7192 20102 7202 20154
rect 7202 20102 7248 20154
rect 6952 20100 7008 20102
rect 7032 20100 7088 20102
rect 7112 20100 7168 20102
rect 7192 20100 7248 20102
rect 6952 19066 7008 19068
rect 7032 19066 7088 19068
rect 7112 19066 7168 19068
rect 7192 19066 7248 19068
rect 6952 19014 6998 19066
rect 6998 19014 7008 19066
rect 7032 19014 7062 19066
rect 7062 19014 7074 19066
rect 7074 19014 7088 19066
rect 7112 19014 7126 19066
rect 7126 19014 7138 19066
rect 7138 19014 7168 19066
rect 7192 19014 7202 19066
rect 7202 19014 7248 19066
rect 6952 19012 7008 19014
rect 7032 19012 7088 19014
rect 7112 19012 7168 19014
rect 7192 19012 7248 19014
rect 6952 17978 7008 17980
rect 7032 17978 7088 17980
rect 7112 17978 7168 17980
rect 7192 17978 7248 17980
rect 6952 17926 6998 17978
rect 6998 17926 7008 17978
rect 7032 17926 7062 17978
rect 7062 17926 7074 17978
rect 7074 17926 7088 17978
rect 7112 17926 7126 17978
rect 7126 17926 7138 17978
rect 7138 17926 7168 17978
rect 7192 17926 7202 17978
rect 7202 17926 7248 17978
rect 6952 17924 7008 17926
rect 7032 17924 7088 17926
rect 7112 17924 7168 17926
rect 7192 17924 7248 17926
rect 6952 16890 7008 16892
rect 7032 16890 7088 16892
rect 7112 16890 7168 16892
rect 7192 16890 7248 16892
rect 6952 16838 6998 16890
rect 6998 16838 7008 16890
rect 7032 16838 7062 16890
rect 7062 16838 7074 16890
rect 7074 16838 7088 16890
rect 7112 16838 7126 16890
rect 7126 16838 7138 16890
rect 7138 16838 7168 16890
rect 7192 16838 7202 16890
rect 7202 16838 7248 16890
rect 6952 16836 7008 16838
rect 7032 16836 7088 16838
rect 7112 16836 7168 16838
rect 7192 16836 7248 16838
rect 6952 15802 7008 15804
rect 7032 15802 7088 15804
rect 7112 15802 7168 15804
rect 7192 15802 7248 15804
rect 6952 15750 6998 15802
rect 6998 15750 7008 15802
rect 7032 15750 7062 15802
rect 7062 15750 7074 15802
rect 7074 15750 7088 15802
rect 7112 15750 7126 15802
rect 7126 15750 7138 15802
rect 7138 15750 7168 15802
rect 7192 15750 7202 15802
rect 7202 15750 7248 15802
rect 6952 15748 7008 15750
rect 7032 15748 7088 15750
rect 7112 15748 7168 15750
rect 7192 15748 7248 15750
rect 6292 15258 6348 15260
rect 6372 15258 6428 15260
rect 6452 15258 6508 15260
rect 6532 15258 6588 15260
rect 6292 15206 6338 15258
rect 6338 15206 6348 15258
rect 6372 15206 6402 15258
rect 6402 15206 6414 15258
rect 6414 15206 6428 15258
rect 6452 15206 6466 15258
rect 6466 15206 6478 15258
rect 6478 15206 6508 15258
rect 6532 15206 6542 15258
rect 6542 15206 6588 15258
rect 6292 15204 6348 15206
rect 6372 15204 6428 15206
rect 6452 15204 6508 15206
rect 6532 15204 6588 15206
rect 9218 27512 9274 27568
rect 11058 27648 11114 27704
rect 9862 24656 9918 24712
rect 6952 14714 7008 14716
rect 7032 14714 7088 14716
rect 7112 14714 7168 14716
rect 7192 14714 7248 14716
rect 6952 14662 6998 14714
rect 6998 14662 7008 14714
rect 7032 14662 7062 14714
rect 7062 14662 7074 14714
rect 7074 14662 7088 14714
rect 7112 14662 7126 14714
rect 7126 14662 7138 14714
rect 7138 14662 7168 14714
rect 7192 14662 7202 14714
rect 7202 14662 7248 14714
rect 6952 14660 7008 14662
rect 7032 14660 7088 14662
rect 7112 14660 7168 14662
rect 7192 14660 7248 14662
rect 6292 14170 6348 14172
rect 6372 14170 6428 14172
rect 6452 14170 6508 14172
rect 6532 14170 6588 14172
rect 6292 14118 6338 14170
rect 6338 14118 6348 14170
rect 6372 14118 6402 14170
rect 6402 14118 6414 14170
rect 6414 14118 6428 14170
rect 6452 14118 6466 14170
rect 6466 14118 6478 14170
rect 6478 14118 6508 14170
rect 6532 14118 6542 14170
rect 6542 14118 6588 14170
rect 6292 14116 6348 14118
rect 6372 14116 6428 14118
rect 6452 14116 6508 14118
rect 6532 14116 6588 14118
rect 6292 13082 6348 13084
rect 6372 13082 6428 13084
rect 6452 13082 6508 13084
rect 6532 13082 6588 13084
rect 6292 13030 6338 13082
rect 6338 13030 6348 13082
rect 6372 13030 6402 13082
rect 6402 13030 6414 13082
rect 6414 13030 6428 13082
rect 6452 13030 6466 13082
rect 6466 13030 6478 13082
rect 6478 13030 6508 13082
rect 6532 13030 6542 13082
rect 6542 13030 6588 13082
rect 6292 13028 6348 13030
rect 6372 13028 6428 13030
rect 6452 13028 6508 13030
rect 6532 13028 6588 13030
rect 6952 13626 7008 13628
rect 7032 13626 7088 13628
rect 7112 13626 7168 13628
rect 7192 13626 7248 13628
rect 6952 13574 6998 13626
rect 6998 13574 7008 13626
rect 7032 13574 7062 13626
rect 7062 13574 7074 13626
rect 7074 13574 7088 13626
rect 7112 13574 7126 13626
rect 7126 13574 7138 13626
rect 7138 13574 7168 13626
rect 7192 13574 7202 13626
rect 7202 13574 7248 13626
rect 6952 13572 7008 13574
rect 7032 13572 7088 13574
rect 7112 13572 7168 13574
rect 7192 13572 7248 13574
rect 6952 12538 7008 12540
rect 7032 12538 7088 12540
rect 7112 12538 7168 12540
rect 7192 12538 7248 12540
rect 6952 12486 6998 12538
rect 6998 12486 7008 12538
rect 7032 12486 7062 12538
rect 7062 12486 7074 12538
rect 7074 12486 7088 12538
rect 7112 12486 7126 12538
rect 7126 12486 7138 12538
rect 7138 12486 7168 12538
rect 7192 12486 7202 12538
rect 7202 12486 7248 12538
rect 6952 12484 7008 12486
rect 7032 12484 7088 12486
rect 7112 12484 7168 12486
rect 7192 12484 7248 12486
rect 6918 12316 6920 12336
rect 6920 12316 6972 12336
rect 6972 12316 6974 12336
rect 6918 12280 6974 12316
rect 6292 11994 6348 11996
rect 6372 11994 6428 11996
rect 6452 11994 6508 11996
rect 6532 11994 6588 11996
rect 6292 11942 6338 11994
rect 6338 11942 6348 11994
rect 6372 11942 6402 11994
rect 6402 11942 6414 11994
rect 6414 11942 6428 11994
rect 6452 11942 6466 11994
rect 6466 11942 6478 11994
rect 6478 11942 6508 11994
rect 6532 11942 6542 11994
rect 6542 11942 6588 11994
rect 6292 11940 6348 11942
rect 6372 11940 6428 11942
rect 6452 11940 6508 11942
rect 6532 11940 6588 11942
rect 6952 11450 7008 11452
rect 7032 11450 7088 11452
rect 7112 11450 7168 11452
rect 7192 11450 7248 11452
rect 6952 11398 6998 11450
rect 6998 11398 7008 11450
rect 7032 11398 7062 11450
rect 7062 11398 7074 11450
rect 7074 11398 7088 11450
rect 7112 11398 7126 11450
rect 7126 11398 7138 11450
rect 7138 11398 7168 11450
rect 7192 11398 7202 11450
rect 7202 11398 7248 11450
rect 6952 11396 7008 11398
rect 7032 11396 7088 11398
rect 7112 11396 7168 11398
rect 7192 11396 7248 11398
rect 6292 10906 6348 10908
rect 6372 10906 6428 10908
rect 6452 10906 6508 10908
rect 6532 10906 6588 10908
rect 6292 10854 6338 10906
rect 6338 10854 6348 10906
rect 6372 10854 6402 10906
rect 6402 10854 6414 10906
rect 6414 10854 6428 10906
rect 6452 10854 6466 10906
rect 6466 10854 6478 10906
rect 6478 10854 6508 10906
rect 6532 10854 6542 10906
rect 6542 10854 6588 10906
rect 6292 10852 6348 10854
rect 6372 10852 6428 10854
rect 6452 10852 6508 10854
rect 6532 10852 6588 10854
rect 6292 9818 6348 9820
rect 6372 9818 6428 9820
rect 6452 9818 6508 9820
rect 6532 9818 6588 9820
rect 6292 9766 6338 9818
rect 6338 9766 6348 9818
rect 6372 9766 6402 9818
rect 6402 9766 6414 9818
rect 6414 9766 6428 9818
rect 6452 9766 6466 9818
rect 6466 9766 6478 9818
rect 6478 9766 6508 9818
rect 6532 9766 6542 9818
rect 6542 9766 6588 9818
rect 6292 9764 6348 9766
rect 6372 9764 6428 9766
rect 6452 9764 6508 9766
rect 6532 9764 6588 9766
rect 6952 10362 7008 10364
rect 7032 10362 7088 10364
rect 7112 10362 7168 10364
rect 7192 10362 7248 10364
rect 6952 10310 6998 10362
rect 6998 10310 7008 10362
rect 7032 10310 7062 10362
rect 7062 10310 7074 10362
rect 7074 10310 7088 10362
rect 7112 10310 7126 10362
rect 7126 10310 7138 10362
rect 7138 10310 7168 10362
rect 7192 10310 7202 10362
rect 7202 10310 7248 10362
rect 6952 10308 7008 10310
rect 7032 10308 7088 10310
rect 7112 10308 7168 10310
rect 7192 10308 7248 10310
rect 6952 9274 7008 9276
rect 7032 9274 7088 9276
rect 7112 9274 7168 9276
rect 7192 9274 7248 9276
rect 6952 9222 6998 9274
rect 6998 9222 7008 9274
rect 7032 9222 7062 9274
rect 7062 9222 7074 9274
rect 7074 9222 7088 9274
rect 7112 9222 7126 9274
rect 7126 9222 7138 9274
rect 7138 9222 7168 9274
rect 7192 9222 7202 9274
rect 7202 9222 7248 9274
rect 6952 9220 7008 9222
rect 7032 9220 7088 9222
rect 7112 9220 7168 9222
rect 7192 9220 7248 9222
rect 9678 20440 9734 20496
rect 9954 23160 10010 23216
rect 9862 19216 9918 19272
rect 7746 14340 7802 14376
rect 7746 14320 7748 14340
rect 7748 14320 7800 14340
rect 7800 14320 7802 14340
rect 8114 12436 8170 12472
rect 8114 12416 8116 12436
rect 8116 12416 8168 12436
rect 8168 12416 8170 12436
rect 6292 8730 6348 8732
rect 6372 8730 6428 8732
rect 6452 8730 6508 8732
rect 6532 8730 6588 8732
rect 6292 8678 6338 8730
rect 6338 8678 6348 8730
rect 6372 8678 6402 8730
rect 6402 8678 6414 8730
rect 6414 8678 6428 8730
rect 6452 8678 6466 8730
rect 6466 8678 6478 8730
rect 6478 8678 6508 8730
rect 6532 8678 6542 8730
rect 6542 8678 6588 8730
rect 6292 8676 6348 8678
rect 6372 8676 6428 8678
rect 6452 8676 6508 8678
rect 6532 8676 6588 8678
rect 6292 7642 6348 7644
rect 6372 7642 6428 7644
rect 6452 7642 6508 7644
rect 6532 7642 6588 7644
rect 6292 7590 6338 7642
rect 6338 7590 6348 7642
rect 6372 7590 6402 7642
rect 6402 7590 6414 7642
rect 6414 7590 6428 7642
rect 6452 7590 6466 7642
rect 6466 7590 6478 7642
rect 6478 7590 6508 7642
rect 6532 7590 6542 7642
rect 6542 7590 6588 7642
rect 6292 7588 6348 7590
rect 6372 7588 6428 7590
rect 6452 7588 6508 7590
rect 6532 7588 6588 7590
rect 6292 6554 6348 6556
rect 6372 6554 6428 6556
rect 6452 6554 6508 6556
rect 6532 6554 6588 6556
rect 6292 6502 6338 6554
rect 6338 6502 6348 6554
rect 6372 6502 6402 6554
rect 6402 6502 6414 6554
rect 6414 6502 6428 6554
rect 6452 6502 6466 6554
rect 6466 6502 6478 6554
rect 6478 6502 6508 6554
rect 6532 6502 6542 6554
rect 6542 6502 6588 6554
rect 6292 6500 6348 6502
rect 6372 6500 6428 6502
rect 6452 6500 6508 6502
rect 6532 6500 6588 6502
rect 6292 5466 6348 5468
rect 6372 5466 6428 5468
rect 6452 5466 6508 5468
rect 6532 5466 6588 5468
rect 6292 5414 6338 5466
rect 6338 5414 6348 5466
rect 6372 5414 6402 5466
rect 6402 5414 6414 5466
rect 6414 5414 6428 5466
rect 6452 5414 6466 5466
rect 6466 5414 6478 5466
rect 6478 5414 6508 5466
rect 6532 5414 6542 5466
rect 6542 5414 6588 5466
rect 6292 5412 6348 5414
rect 6372 5412 6428 5414
rect 6452 5412 6508 5414
rect 6532 5412 6588 5414
rect 6952 8186 7008 8188
rect 7032 8186 7088 8188
rect 7112 8186 7168 8188
rect 7192 8186 7248 8188
rect 6952 8134 6998 8186
rect 6998 8134 7008 8186
rect 7032 8134 7062 8186
rect 7062 8134 7074 8186
rect 7074 8134 7088 8186
rect 7112 8134 7126 8186
rect 7126 8134 7138 8186
rect 7138 8134 7168 8186
rect 7192 8134 7202 8186
rect 7202 8134 7248 8186
rect 6952 8132 7008 8134
rect 7032 8132 7088 8134
rect 7112 8132 7168 8134
rect 7192 8132 7248 8134
rect 6952 7098 7008 7100
rect 7032 7098 7088 7100
rect 7112 7098 7168 7100
rect 7192 7098 7248 7100
rect 6952 7046 6998 7098
rect 6998 7046 7008 7098
rect 7032 7046 7062 7098
rect 7062 7046 7074 7098
rect 7074 7046 7088 7098
rect 7112 7046 7126 7098
rect 7126 7046 7138 7098
rect 7138 7046 7168 7098
rect 7192 7046 7202 7098
rect 7202 7046 7248 7098
rect 6952 7044 7008 7046
rect 7032 7044 7088 7046
rect 7112 7044 7168 7046
rect 7192 7044 7248 7046
rect 6952 6010 7008 6012
rect 7032 6010 7088 6012
rect 7112 6010 7168 6012
rect 7192 6010 7248 6012
rect 6952 5958 6998 6010
rect 6998 5958 7008 6010
rect 7032 5958 7062 6010
rect 7062 5958 7074 6010
rect 7074 5958 7088 6010
rect 7112 5958 7126 6010
rect 7126 5958 7138 6010
rect 7138 5958 7168 6010
rect 7192 5958 7202 6010
rect 7202 5958 7248 6010
rect 6952 5956 7008 5958
rect 7032 5956 7088 5958
rect 7112 5956 7168 5958
rect 7192 5956 7248 5958
rect 6292 4378 6348 4380
rect 6372 4378 6428 4380
rect 6452 4378 6508 4380
rect 6532 4378 6588 4380
rect 6292 4326 6338 4378
rect 6338 4326 6348 4378
rect 6372 4326 6402 4378
rect 6402 4326 6414 4378
rect 6414 4326 6428 4378
rect 6452 4326 6466 4378
rect 6466 4326 6478 4378
rect 6478 4326 6508 4378
rect 6532 4326 6542 4378
rect 6542 4326 6588 4378
rect 6292 4324 6348 4326
rect 6372 4324 6428 4326
rect 6452 4324 6508 4326
rect 6532 4324 6588 4326
rect 6952 4922 7008 4924
rect 7032 4922 7088 4924
rect 7112 4922 7168 4924
rect 7192 4922 7248 4924
rect 6952 4870 6998 4922
rect 6998 4870 7008 4922
rect 7032 4870 7062 4922
rect 7062 4870 7074 4922
rect 7074 4870 7088 4922
rect 7112 4870 7126 4922
rect 7126 4870 7138 4922
rect 7138 4870 7168 4922
rect 7192 4870 7202 4922
rect 7202 4870 7248 4922
rect 6952 4868 7008 4870
rect 7032 4868 7088 4870
rect 7112 4868 7168 4870
rect 7192 4868 7248 4870
rect 6952 3834 7008 3836
rect 7032 3834 7088 3836
rect 7112 3834 7168 3836
rect 7192 3834 7248 3836
rect 6952 3782 6998 3834
rect 6998 3782 7008 3834
rect 7032 3782 7062 3834
rect 7062 3782 7074 3834
rect 7074 3782 7088 3834
rect 7112 3782 7126 3834
rect 7126 3782 7138 3834
rect 7138 3782 7168 3834
rect 7192 3782 7202 3834
rect 7202 3782 7248 3834
rect 6952 3780 7008 3782
rect 7032 3780 7088 3782
rect 7112 3780 7168 3782
rect 7192 3780 7248 3782
rect 3606 2760 3662 2816
rect 3054 1400 3110 1456
rect 6292 3290 6348 3292
rect 6372 3290 6428 3292
rect 6452 3290 6508 3292
rect 6532 3290 6588 3292
rect 6292 3238 6338 3290
rect 6338 3238 6348 3290
rect 6372 3238 6402 3290
rect 6402 3238 6414 3290
rect 6414 3238 6428 3290
rect 6452 3238 6466 3290
rect 6466 3238 6478 3290
rect 6478 3238 6508 3290
rect 6532 3238 6542 3290
rect 6542 3238 6588 3290
rect 6292 3236 6348 3238
rect 6372 3236 6428 3238
rect 6452 3236 6508 3238
rect 6532 3236 6588 3238
rect 14312 32122 14368 32124
rect 14392 32122 14448 32124
rect 14472 32122 14528 32124
rect 14552 32122 14608 32124
rect 14312 32070 14358 32122
rect 14358 32070 14368 32122
rect 14392 32070 14422 32122
rect 14422 32070 14434 32122
rect 14434 32070 14448 32122
rect 14472 32070 14486 32122
rect 14486 32070 14498 32122
rect 14498 32070 14528 32122
rect 14552 32070 14562 32122
rect 14562 32070 14608 32122
rect 14312 32068 14368 32070
rect 14392 32068 14448 32070
rect 14472 32068 14528 32070
rect 14552 32068 14608 32070
rect 13652 31578 13708 31580
rect 13732 31578 13788 31580
rect 13812 31578 13868 31580
rect 13892 31578 13948 31580
rect 13652 31526 13698 31578
rect 13698 31526 13708 31578
rect 13732 31526 13762 31578
rect 13762 31526 13774 31578
rect 13774 31526 13788 31578
rect 13812 31526 13826 31578
rect 13826 31526 13838 31578
rect 13838 31526 13868 31578
rect 13892 31526 13902 31578
rect 13902 31526 13948 31578
rect 13652 31524 13708 31526
rect 13732 31524 13788 31526
rect 13812 31524 13868 31526
rect 13892 31524 13948 31526
rect 11334 25744 11390 25800
rect 11058 24112 11114 24168
rect 10966 16652 11022 16688
rect 10966 16632 10968 16652
rect 10968 16632 11020 16652
rect 11020 16632 11022 16652
rect 10414 16516 10470 16552
rect 10414 16496 10416 16516
rect 10416 16496 10468 16516
rect 10468 16496 10470 16516
rect 11610 23704 11666 23760
rect 11794 24112 11850 24168
rect 12254 24676 12310 24712
rect 12254 24656 12256 24676
rect 12256 24656 12308 24676
rect 12308 24656 12310 24676
rect 11610 19896 11666 19952
rect 12162 22480 12218 22536
rect 11518 14900 11520 14920
rect 11520 14900 11572 14920
rect 11572 14900 11574 14920
rect 11518 14864 11574 14900
rect 13652 30490 13708 30492
rect 13732 30490 13788 30492
rect 13812 30490 13868 30492
rect 13892 30490 13948 30492
rect 13652 30438 13698 30490
rect 13698 30438 13708 30490
rect 13732 30438 13762 30490
rect 13762 30438 13774 30490
rect 13774 30438 13788 30490
rect 13812 30438 13826 30490
rect 13826 30438 13838 30490
rect 13838 30438 13868 30490
rect 13892 30438 13902 30490
rect 13902 30438 13948 30490
rect 13652 30436 13708 30438
rect 13732 30436 13788 30438
rect 13812 30436 13868 30438
rect 13892 30436 13948 30438
rect 14554 31340 14610 31376
rect 14554 31320 14556 31340
rect 14556 31320 14608 31340
rect 14608 31320 14610 31340
rect 14312 31034 14368 31036
rect 14392 31034 14448 31036
rect 14472 31034 14528 31036
rect 14552 31034 14608 31036
rect 14312 30982 14358 31034
rect 14358 30982 14368 31034
rect 14392 30982 14422 31034
rect 14422 30982 14434 31034
rect 14434 30982 14448 31034
rect 14472 30982 14486 31034
rect 14486 30982 14498 31034
rect 14498 30982 14528 31034
rect 14552 30982 14562 31034
rect 14562 30982 14608 31034
rect 14312 30980 14368 30982
rect 14392 30980 14448 30982
rect 14472 30980 14528 30982
rect 14552 30980 14608 30982
rect 14312 29946 14368 29948
rect 14392 29946 14448 29948
rect 14472 29946 14528 29948
rect 14552 29946 14608 29948
rect 14312 29894 14358 29946
rect 14358 29894 14368 29946
rect 14392 29894 14422 29946
rect 14422 29894 14434 29946
rect 14434 29894 14448 29946
rect 14472 29894 14486 29946
rect 14486 29894 14498 29946
rect 14498 29894 14528 29946
rect 14552 29894 14562 29946
rect 14562 29894 14608 29946
rect 14312 29892 14368 29894
rect 14392 29892 14448 29894
rect 14472 29892 14528 29894
rect 14552 29892 14608 29894
rect 13652 29402 13708 29404
rect 13732 29402 13788 29404
rect 13812 29402 13868 29404
rect 13892 29402 13948 29404
rect 13652 29350 13698 29402
rect 13698 29350 13708 29402
rect 13732 29350 13762 29402
rect 13762 29350 13774 29402
rect 13774 29350 13788 29402
rect 13812 29350 13826 29402
rect 13826 29350 13838 29402
rect 13838 29350 13868 29402
rect 13892 29350 13902 29402
rect 13902 29350 13948 29402
rect 13652 29348 13708 29350
rect 13732 29348 13788 29350
rect 13812 29348 13868 29350
rect 13892 29348 13948 29350
rect 13652 28314 13708 28316
rect 13732 28314 13788 28316
rect 13812 28314 13868 28316
rect 13892 28314 13948 28316
rect 13652 28262 13698 28314
rect 13698 28262 13708 28314
rect 13732 28262 13762 28314
rect 13762 28262 13774 28314
rect 13774 28262 13788 28314
rect 13812 28262 13826 28314
rect 13826 28262 13838 28314
rect 13838 28262 13868 28314
rect 13892 28262 13902 28314
rect 13902 28262 13948 28314
rect 13652 28260 13708 28262
rect 13732 28260 13788 28262
rect 13812 28260 13868 28262
rect 13892 28260 13948 28262
rect 14312 28858 14368 28860
rect 14392 28858 14448 28860
rect 14472 28858 14528 28860
rect 14552 28858 14608 28860
rect 14312 28806 14358 28858
rect 14358 28806 14368 28858
rect 14392 28806 14422 28858
rect 14422 28806 14434 28858
rect 14434 28806 14448 28858
rect 14472 28806 14486 28858
rect 14486 28806 14498 28858
rect 14498 28806 14528 28858
rect 14552 28806 14562 28858
rect 14562 28806 14608 28858
rect 14312 28804 14368 28806
rect 14392 28804 14448 28806
rect 14472 28804 14528 28806
rect 14552 28804 14608 28806
rect 14312 27770 14368 27772
rect 14392 27770 14448 27772
rect 14472 27770 14528 27772
rect 14552 27770 14608 27772
rect 14312 27718 14358 27770
rect 14358 27718 14368 27770
rect 14392 27718 14422 27770
rect 14422 27718 14434 27770
rect 14434 27718 14448 27770
rect 14472 27718 14486 27770
rect 14486 27718 14498 27770
rect 14498 27718 14528 27770
rect 14552 27718 14562 27770
rect 14562 27718 14608 27770
rect 14312 27716 14368 27718
rect 14392 27716 14448 27718
rect 14472 27716 14528 27718
rect 14552 27716 14608 27718
rect 13652 27226 13708 27228
rect 13732 27226 13788 27228
rect 13812 27226 13868 27228
rect 13892 27226 13948 27228
rect 13652 27174 13698 27226
rect 13698 27174 13708 27226
rect 13732 27174 13762 27226
rect 13762 27174 13774 27226
rect 13774 27174 13788 27226
rect 13812 27174 13826 27226
rect 13826 27174 13838 27226
rect 13838 27174 13868 27226
rect 13892 27174 13902 27226
rect 13902 27174 13948 27226
rect 13652 27172 13708 27174
rect 13732 27172 13788 27174
rect 13812 27172 13868 27174
rect 13892 27172 13948 27174
rect 13652 26138 13708 26140
rect 13732 26138 13788 26140
rect 13812 26138 13868 26140
rect 13892 26138 13948 26140
rect 13652 26086 13698 26138
rect 13698 26086 13708 26138
rect 13732 26086 13762 26138
rect 13762 26086 13774 26138
rect 13774 26086 13788 26138
rect 13812 26086 13826 26138
rect 13826 26086 13838 26138
rect 13838 26086 13868 26138
rect 13892 26086 13902 26138
rect 13902 26086 13948 26138
rect 13652 26084 13708 26086
rect 13732 26084 13788 26086
rect 13812 26084 13868 26086
rect 13892 26084 13948 26086
rect 14312 26682 14368 26684
rect 14392 26682 14448 26684
rect 14472 26682 14528 26684
rect 14552 26682 14608 26684
rect 14312 26630 14358 26682
rect 14358 26630 14368 26682
rect 14392 26630 14422 26682
rect 14422 26630 14434 26682
rect 14434 26630 14448 26682
rect 14472 26630 14486 26682
rect 14486 26630 14498 26682
rect 14498 26630 14528 26682
rect 14552 26630 14562 26682
rect 14562 26630 14608 26682
rect 14312 26628 14368 26630
rect 14392 26628 14448 26630
rect 14472 26628 14528 26630
rect 14552 26628 14608 26630
rect 13652 25050 13708 25052
rect 13732 25050 13788 25052
rect 13812 25050 13868 25052
rect 13892 25050 13948 25052
rect 13652 24998 13698 25050
rect 13698 24998 13708 25050
rect 13732 24998 13762 25050
rect 13762 24998 13774 25050
rect 13774 24998 13788 25050
rect 13812 24998 13826 25050
rect 13826 24998 13838 25050
rect 13838 24998 13868 25050
rect 13892 24998 13902 25050
rect 13902 24998 13948 25050
rect 13652 24996 13708 24998
rect 13732 24996 13788 24998
rect 13812 24996 13868 24998
rect 13892 24996 13948 24998
rect 13652 23962 13708 23964
rect 13732 23962 13788 23964
rect 13812 23962 13868 23964
rect 13892 23962 13948 23964
rect 13652 23910 13698 23962
rect 13698 23910 13708 23962
rect 13732 23910 13762 23962
rect 13762 23910 13774 23962
rect 13774 23910 13788 23962
rect 13812 23910 13826 23962
rect 13826 23910 13838 23962
rect 13838 23910 13868 23962
rect 13892 23910 13902 23962
rect 13902 23910 13948 23962
rect 13652 23908 13708 23910
rect 13732 23908 13788 23910
rect 13812 23908 13868 23910
rect 13892 23908 13948 23910
rect 13542 23024 13598 23080
rect 13652 22874 13708 22876
rect 13732 22874 13788 22876
rect 13812 22874 13868 22876
rect 13892 22874 13948 22876
rect 13652 22822 13698 22874
rect 13698 22822 13708 22874
rect 13732 22822 13762 22874
rect 13762 22822 13774 22874
rect 13774 22822 13788 22874
rect 13812 22822 13826 22874
rect 13826 22822 13838 22874
rect 13838 22822 13868 22874
rect 13892 22822 13902 22874
rect 13902 22822 13948 22874
rect 13652 22820 13708 22822
rect 13732 22820 13788 22822
rect 13812 22820 13868 22822
rect 13892 22820 13948 22822
rect 12990 19760 13046 19816
rect 13082 19352 13138 19408
rect 11794 15000 11850 15056
rect 13652 21786 13708 21788
rect 13732 21786 13788 21788
rect 13812 21786 13868 21788
rect 13892 21786 13948 21788
rect 13652 21734 13698 21786
rect 13698 21734 13708 21786
rect 13732 21734 13762 21786
rect 13762 21734 13774 21786
rect 13774 21734 13788 21786
rect 13812 21734 13826 21786
rect 13826 21734 13838 21786
rect 13838 21734 13868 21786
rect 13892 21734 13902 21786
rect 13902 21734 13948 21786
rect 13652 21732 13708 21734
rect 13732 21732 13788 21734
rect 13812 21732 13868 21734
rect 13892 21732 13948 21734
rect 14312 25594 14368 25596
rect 14392 25594 14448 25596
rect 14472 25594 14528 25596
rect 14552 25594 14608 25596
rect 14312 25542 14358 25594
rect 14358 25542 14368 25594
rect 14392 25542 14422 25594
rect 14422 25542 14434 25594
rect 14434 25542 14448 25594
rect 14472 25542 14486 25594
rect 14486 25542 14498 25594
rect 14498 25542 14528 25594
rect 14552 25542 14562 25594
rect 14562 25542 14608 25594
rect 14312 25540 14368 25542
rect 14392 25540 14448 25542
rect 14472 25540 14528 25542
rect 14552 25540 14608 25542
rect 14312 24506 14368 24508
rect 14392 24506 14448 24508
rect 14472 24506 14528 24508
rect 14552 24506 14608 24508
rect 14312 24454 14358 24506
rect 14358 24454 14368 24506
rect 14392 24454 14422 24506
rect 14422 24454 14434 24506
rect 14434 24454 14448 24506
rect 14472 24454 14486 24506
rect 14486 24454 14498 24506
rect 14498 24454 14528 24506
rect 14552 24454 14562 24506
rect 14562 24454 14608 24506
rect 14312 24452 14368 24454
rect 14392 24452 14448 24454
rect 14472 24452 14528 24454
rect 14552 24452 14608 24454
rect 15106 26288 15162 26344
rect 16578 28056 16634 28112
rect 14312 23418 14368 23420
rect 14392 23418 14448 23420
rect 14472 23418 14528 23420
rect 14552 23418 14608 23420
rect 14312 23366 14358 23418
rect 14358 23366 14368 23418
rect 14392 23366 14422 23418
rect 14422 23366 14434 23418
rect 14434 23366 14448 23418
rect 14472 23366 14486 23418
rect 14486 23366 14498 23418
rect 14498 23366 14528 23418
rect 14552 23366 14562 23418
rect 14562 23366 14608 23418
rect 14312 23364 14368 23366
rect 14392 23364 14448 23366
rect 14472 23364 14528 23366
rect 14552 23364 14608 23366
rect 14370 23180 14426 23216
rect 14370 23160 14372 23180
rect 14372 23160 14424 23180
rect 14424 23160 14426 23180
rect 15198 24112 15254 24168
rect 14462 22480 14518 22536
rect 14312 22330 14368 22332
rect 14392 22330 14448 22332
rect 14472 22330 14528 22332
rect 14552 22330 14608 22332
rect 14312 22278 14358 22330
rect 14358 22278 14368 22330
rect 14392 22278 14422 22330
rect 14422 22278 14434 22330
rect 14434 22278 14448 22330
rect 14472 22278 14486 22330
rect 14486 22278 14498 22330
rect 14498 22278 14528 22330
rect 14552 22278 14562 22330
rect 14562 22278 14608 22330
rect 14312 22276 14368 22278
rect 14392 22276 14448 22278
rect 14472 22276 14528 22278
rect 14552 22276 14608 22278
rect 14312 21242 14368 21244
rect 14392 21242 14448 21244
rect 14472 21242 14528 21244
rect 14552 21242 14608 21244
rect 14312 21190 14358 21242
rect 14358 21190 14368 21242
rect 14392 21190 14422 21242
rect 14422 21190 14434 21242
rect 14434 21190 14448 21242
rect 14472 21190 14486 21242
rect 14486 21190 14498 21242
rect 14498 21190 14528 21242
rect 14552 21190 14562 21242
rect 14562 21190 14608 21242
rect 14312 21188 14368 21190
rect 14392 21188 14448 21190
rect 14472 21188 14528 21190
rect 14552 21188 14608 21190
rect 13818 20884 13820 20904
rect 13820 20884 13872 20904
rect 13872 20884 13874 20904
rect 13818 20848 13874 20884
rect 13652 20698 13708 20700
rect 13732 20698 13788 20700
rect 13812 20698 13868 20700
rect 13892 20698 13948 20700
rect 13652 20646 13698 20698
rect 13698 20646 13708 20698
rect 13732 20646 13762 20698
rect 13762 20646 13774 20698
rect 13774 20646 13788 20698
rect 13812 20646 13826 20698
rect 13826 20646 13838 20698
rect 13838 20646 13868 20698
rect 13892 20646 13902 20698
rect 13902 20646 13948 20698
rect 13652 20644 13708 20646
rect 13732 20644 13788 20646
rect 13812 20644 13868 20646
rect 13892 20644 13948 20646
rect 13652 19610 13708 19612
rect 13732 19610 13788 19612
rect 13812 19610 13868 19612
rect 13892 19610 13948 19612
rect 13652 19558 13698 19610
rect 13698 19558 13708 19610
rect 13732 19558 13762 19610
rect 13762 19558 13774 19610
rect 13774 19558 13788 19610
rect 13812 19558 13826 19610
rect 13826 19558 13838 19610
rect 13838 19558 13868 19610
rect 13892 19558 13902 19610
rect 13902 19558 13948 19610
rect 13652 19556 13708 19558
rect 13732 19556 13788 19558
rect 13812 19556 13868 19558
rect 13892 19556 13948 19558
rect 13542 19352 13598 19408
rect 13082 17176 13138 17232
rect 11058 12416 11114 12472
rect 12530 16496 12586 16552
rect 15106 22208 15162 22264
rect 14738 20712 14794 20768
rect 14312 20154 14368 20156
rect 14392 20154 14448 20156
rect 14472 20154 14528 20156
rect 14552 20154 14608 20156
rect 14312 20102 14358 20154
rect 14358 20102 14368 20154
rect 14392 20102 14422 20154
rect 14422 20102 14434 20154
rect 14434 20102 14448 20154
rect 14472 20102 14486 20154
rect 14486 20102 14498 20154
rect 14498 20102 14528 20154
rect 14552 20102 14562 20154
rect 14562 20102 14608 20154
rect 14312 20100 14368 20102
rect 14392 20100 14448 20102
rect 14472 20100 14528 20102
rect 14552 20100 14608 20102
rect 14738 19352 14794 19408
rect 14554 19216 14610 19272
rect 14738 19252 14740 19272
rect 14740 19252 14792 19272
rect 14792 19252 14794 19272
rect 14738 19216 14794 19252
rect 14312 19066 14368 19068
rect 14392 19066 14448 19068
rect 14472 19066 14528 19068
rect 14552 19066 14608 19068
rect 14312 19014 14358 19066
rect 14358 19014 14368 19066
rect 14392 19014 14422 19066
rect 14422 19014 14434 19066
rect 14434 19014 14448 19066
rect 14472 19014 14486 19066
rect 14486 19014 14498 19066
rect 14498 19014 14528 19066
rect 14552 19014 14562 19066
rect 14562 19014 14608 19066
rect 14312 19012 14368 19014
rect 14392 19012 14448 19014
rect 14472 19012 14528 19014
rect 14552 19012 14608 19014
rect 14370 18808 14426 18864
rect 13652 18522 13708 18524
rect 13732 18522 13788 18524
rect 13812 18522 13868 18524
rect 13892 18522 13948 18524
rect 13652 18470 13698 18522
rect 13698 18470 13708 18522
rect 13732 18470 13762 18522
rect 13762 18470 13774 18522
rect 13774 18470 13788 18522
rect 13812 18470 13826 18522
rect 13826 18470 13838 18522
rect 13838 18470 13868 18522
rect 13892 18470 13902 18522
rect 13902 18470 13948 18522
rect 13652 18468 13708 18470
rect 13732 18468 13788 18470
rect 13812 18468 13868 18470
rect 13892 18468 13948 18470
rect 14002 17720 14058 17776
rect 14370 18128 14426 18184
rect 14312 17978 14368 17980
rect 14392 17978 14448 17980
rect 14472 17978 14528 17980
rect 14552 17978 14608 17980
rect 14312 17926 14358 17978
rect 14358 17926 14368 17978
rect 14392 17926 14422 17978
rect 14422 17926 14434 17978
rect 14434 17926 14448 17978
rect 14472 17926 14486 17978
rect 14486 17926 14498 17978
rect 14498 17926 14528 17978
rect 14552 17926 14562 17978
rect 14562 17926 14608 17978
rect 14312 17924 14368 17926
rect 14392 17924 14448 17926
rect 14472 17924 14528 17926
rect 14552 17924 14608 17926
rect 13652 17434 13708 17436
rect 13732 17434 13788 17436
rect 13812 17434 13868 17436
rect 13892 17434 13948 17436
rect 13652 17382 13698 17434
rect 13698 17382 13708 17434
rect 13732 17382 13762 17434
rect 13762 17382 13774 17434
rect 13774 17382 13788 17434
rect 13812 17382 13826 17434
rect 13826 17382 13838 17434
rect 13838 17382 13868 17434
rect 13892 17382 13902 17434
rect 13902 17382 13948 17434
rect 13652 17380 13708 17382
rect 13732 17380 13788 17382
rect 13812 17380 13868 17382
rect 13892 17380 13948 17382
rect 14094 17312 14150 17368
rect 13358 17076 13360 17096
rect 13360 17076 13412 17096
rect 13412 17076 13414 17096
rect 13358 17040 13414 17076
rect 12254 14184 12310 14240
rect 13652 16346 13708 16348
rect 13732 16346 13788 16348
rect 13812 16346 13868 16348
rect 13892 16346 13948 16348
rect 13652 16294 13698 16346
rect 13698 16294 13708 16346
rect 13732 16294 13762 16346
rect 13762 16294 13774 16346
rect 13774 16294 13788 16346
rect 13812 16294 13826 16346
rect 13826 16294 13838 16346
rect 13838 16294 13868 16346
rect 13892 16294 13902 16346
rect 13902 16294 13948 16346
rect 13652 16292 13708 16294
rect 13732 16292 13788 16294
rect 13812 16292 13868 16294
rect 13892 16292 13948 16294
rect 14554 17312 14610 17368
rect 15290 21120 15346 21176
rect 16118 23704 16174 23760
rect 16394 22208 16450 22264
rect 15198 19896 15254 19952
rect 15106 18264 15162 18320
rect 14312 16890 14368 16892
rect 14392 16890 14448 16892
rect 14472 16890 14528 16892
rect 14552 16890 14608 16892
rect 14312 16838 14358 16890
rect 14358 16838 14368 16890
rect 14392 16838 14422 16890
rect 14422 16838 14434 16890
rect 14434 16838 14448 16890
rect 14472 16838 14486 16890
rect 14486 16838 14498 16890
rect 14498 16838 14528 16890
rect 14552 16838 14562 16890
rect 14562 16838 14608 16890
rect 14312 16836 14368 16838
rect 14392 16836 14448 16838
rect 14472 16836 14528 16838
rect 14552 16836 14608 16838
rect 12806 14764 12808 14784
rect 12808 14764 12860 14784
rect 12860 14764 12862 14784
rect 12806 14728 12862 14764
rect 14094 16088 14150 16144
rect 14312 15802 14368 15804
rect 14392 15802 14448 15804
rect 14472 15802 14528 15804
rect 14552 15802 14608 15804
rect 14312 15750 14358 15802
rect 14358 15750 14368 15802
rect 14392 15750 14422 15802
rect 14422 15750 14434 15802
rect 14434 15750 14448 15802
rect 14472 15750 14486 15802
rect 14486 15750 14498 15802
rect 14498 15750 14528 15802
rect 14552 15750 14562 15802
rect 14562 15750 14608 15802
rect 14312 15748 14368 15750
rect 14392 15748 14448 15750
rect 14472 15748 14528 15750
rect 14552 15748 14608 15750
rect 13358 15000 13414 15056
rect 13358 14728 13414 14784
rect 13652 15258 13708 15260
rect 13732 15258 13788 15260
rect 13812 15258 13868 15260
rect 13892 15258 13948 15260
rect 13652 15206 13698 15258
rect 13698 15206 13708 15258
rect 13732 15206 13762 15258
rect 13762 15206 13774 15258
rect 13774 15206 13788 15258
rect 13812 15206 13826 15258
rect 13826 15206 13838 15258
rect 13838 15206 13868 15258
rect 13892 15206 13902 15258
rect 13902 15206 13948 15258
rect 13652 15204 13708 15206
rect 13732 15204 13788 15206
rect 13812 15204 13868 15206
rect 13892 15204 13948 15206
rect 14094 14864 14150 14920
rect 14312 14714 14368 14716
rect 14392 14714 14448 14716
rect 14472 14714 14528 14716
rect 14552 14714 14608 14716
rect 14312 14662 14358 14714
rect 14358 14662 14368 14714
rect 14392 14662 14422 14714
rect 14422 14662 14434 14714
rect 14434 14662 14448 14714
rect 14472 14662 14486 14714
rect 14486 14662 14498 14714
rect 14498 14662 14528 14714
rect 14552 14662 14562 14714
rect 14562 14662 14608 14714
rect 14312 14660 14368 14662
rect 14392 14660 14448 14662
rect 14472 14660 14528 14662
rect 14552 14660 14608 14662
rect 13652 14170 13708 14172
rect 13732 14170 13788 14172
rect 13812 14170 13868 14172
rect 13892 14170 13948 14172
rect 13652 14118 13698 14170
rect 13698 14118 13708 14170
rect 13732 14118 13762 14170
rect 13762 14118 13774 14170
rect 13774 14118 13788 14170
rect 13812 14118 13826 14170
rect 13826 14118 13838 14170
rect 13838 14118 13868 14170
rect 13892 14118 13902 14170
rect 13902 14118 13948 14170
rect 13652 14116 13708 14118
rect 13732 14116 13788 14118
rect 13812 14116 13868 14118
rect 13892 14116 13948 14118
rect 11150 12316 11152 12336
rect 11152 12316 11204 12336
rect 11204 12316 11206 12336
rect 11150 12280 11206 12316
rect 10874 9036 10930 9072
rect 10874 9016 10876 9036
rect 10876 9016 10928 9036
rect 10928 9016 10930 9036
rect 6952 2746 7008 2748
rect 7032 2746 7088 2748
rect 7112 2746 7168 2748
rect 7192 2746 7248 2748
rect 6952 2694 6998 2746
rect 6998 2694 7008 2746
rect 7032 2694 7062 2746
rect 7062 2694 7074 2746
rect 7074 2694 7088 2746
rect 7112 2694 7126 2746
rect 7126 2694 7138 2746
rect 7138 2694 7168 2746
rect 7192 2694 7202 2746
rect 7202 2694 7248 2746
rect 6952 2692 7008 2694
rect 7032 2692 7088 2694
rect 7112 2692 7168 2694
rect 7192 2692 7248 2694
rect 15014 17312 15070 17368
rect 15290 17176 15346 17232
rect 15658 19932 15660 19952
rect 15660 19932 15712 19952
rect 15712 19932 15714 19952
rect 15658 19896 15714 19932
rect 14312 13626 14368 13628
rect 14392 13626 14448 13628
rect 14472 13626 14528 13628
rect 14552 13626 14608 13628
rect 14312 13574 14358 13626
rect 14358 13574 14368 13626
rect 14392 13574 14422 13626
rect 14422 13574 14434 13626
rect 14434 13574 14448 13626
rect 14472 13574 14486 13626
rect 14486 13574 14498 13626
rect 14498 13574 14528 13626
rect 14552 13574 14562 13626
rect 14562 13574 14608 13626
rect 14312 13572 14368 13574
rect 14392 13572 14448 13574
rect 14472 13572 14528 13574
rect 14552 13572 14608 13574
rect 13652 13082 13708 13084
rect 13732 13082 13788 13084
rect 13812 13082 13868 13084
rect 13892 13082 13948 13084
rect 13652 13030 13698 13082
rect 13698 13030 13708 13082
rect 13732 13030 13762 13082
rect 13762 13030 13774 13082
rect 13774 13030 13788 13082
rect 13812 13030 13826 13082
rect 13826 13030 13838 13082
rect 13838 13030 13868 13082
rect 13892 13030 13902 13082
rect 13902 13030 13948 13082
rect 13652 13028 13708 13030
rect 13732 13028 13788 13030
rect 13812 13028 13868 13030
rect 13892 13028 13948 13030
rect 13652 11994 13708 11996
rect 13732 11994 13788 11996
rect 13812 11994 13868 11996
rect 13892 11994 13948 11996
rect 13652 11942 13698 11994
rect 13698 11942 13708 11994
rect 13732 11942 13762 11994
rect 13762 11942 13774 11994
rect 13774 11942 13788 11994
rect 13812 11942 13826 11994
rect 13826 11942 13838 11994
rect 13838 11942 13868 11994
rect 13892 11942 13902 11994
rect 13902 11942 13948 11994
rect 13652 11940 13708 11942
rect 13732 11940 13788 11942
rect 13812 11940 13868 11942
rect 13892 11940 13948 11942
rect 16026 20712 16082 20768
rect 15934 19896 15990 19952
rect 15842 18264 15898 18320
rect 15750 18128 15806 18184
rect 16670 21120 16726 21176
rect 18786 31864 18842 31920
rect 17866 31728 17922 31784
rect 18142 23024 18198 23080
rect 16486 17856 16542 17912
rect 15658 16632 15714 16688
rect 15474 16088 15530 16144
rect 15382 15156 15438 15192
rect 15382 15136 15384 15156
rect 15384 15136 15436 15156
rect 15436 15136 15438 15156
rect 14312 12538 14368 12540
rect 14392 12538 14448 12540
rect 14472 12538 14528 12540
rect 14552 12538 14608 12540
rect 14312 12486 14358 12538
rect 14358 12486 14368 12538
rect 14392 12486 14422 12538
rect 14422 12486 14434 12538
rect 14434 12486 14448 12538
rect 14472 12486 14486 12538
rect 14486 12486 14498 12538
rect 14498 12486 14528 12538
rect 14552 12486 14562 12538
rect 14562 12486 14608 12538
rect 14312 12484 14368 12486
rect 14392 12484 14448 12486
rect 14472 12484 14528 12486
rect 14552 12484 14608 12486
rect 14312 11450 14368 11452
rect 14392 11450 14448 11452
rect 14472 11450 14528 11452
rect 14552 11450 14608 11452
rect 14312 11398 14358 11450
rect 14358 11398 14368 11450
rect 14392 11398 14422 11450
rect 14422 11398 14434 11450
rect 14434 11398 14448 11450
rect 14472 11398 14486 11450
rect 14486 11398 14498 11450
rect 14498 11398 14528 11450
rect 14552 11398 14562 11450
rect 14562 11398 14608 11450
rect 14312 11396 14368 11398
rect 14392 11396 14448 11398
rect 14472 11396 14528 11398
rect 14552 11396 14608 11398
rect 14002 11212 14058 11248
rect 14002 11192 14004 11212
rect 14004 11192 14056 11212
rect 14056 11192 14058 11212
rect 13652 10906 13708 10908
rect 13732 10906 13788 10908
rect 13812 10906 13868 10908
rect 13892 10906 13948 10908
rect 13652 10854 13698 10906
rect 13698 10854 13708 10906
rect 13732 10854 13762 10906
rect 13762 10854 13774 10906
rect 13774 10854 13788 10906
rect 13812 10854 13826 10906
rect 13826 10854 13838 10906
rect 13838 10854 13868 10906
rect 13892 10854 13902 10906
rect 13902 10854 13948 10906
rect 13652 10852 13708 10854
rect 13732 10852 13788 10854
rect 13812 10852 13868 10854
rect 13892 10852 13948 10854
rect 13652 9818 13708 9820
rect 13732 9818 13788 9820
rect 13812 9818 13868 9820
rect 13892 9818 13948 9820
rect 13652 9766 13698 9818
rect 13698 9766 13708 9818
rect 13732 9766 13762 9818
rect 13762 9766 13774 9818
rect 13774 9766 13788 9818
rect 13812 9766 13826 9818
rect 13826 9766 13838 9818
rect 13838 9766 13868 9818
rect 13892 9766 13902 9818
rect 13902 9766 13948 9818
rect 13652 9764 13708 9766
rect 13732 9764 13788 9766
rect 13812 9764 13868 9766
rect 13892 9764 13948 9766
rect 14312 10362 14368 10364
rect 14392 10362 14448 10364
rect 14472 10362 14528 10364
rect 14552 10362 14608 10364
rect 14312 10310 14358 10362
rect 14358 10310 14368 10362
rect 14392 10310 14422 10362
rect 14422 10310 14434 10362
rect 14434 10310 14448 10362
rect 14472 10310 14486 10362
rect 14486 10310 14498 10362
rect 14498 10310 14528 10362
rect 14552 10310 14562 10362
rect 14562 10310 14608 10362
rect 14312 10308 14368 10310
rect 14392 10308 14448 10310
rect 14472 10308 14528 10310
rect 14552 10308 14608 10310
rect 16486 17040 16542 17096
rect 16854 18028 16856 18048
rect 16856 18028 16908 18048
rect 16908 18028 16910 18048
rect 16854 17992 16910 18028
rect 17406 17992 17462 18048
rect 17038 17060 17094 17096
rect 17038 17040 17040 17060
rect 17040 17040 17092 17060
rect 17092 17040 17094 17060
rect 17590 19760 17646 19816
rect 21012 31578 21068 31580
rect 21092 31578 21148 31580
rect 21172 31578 21228 31580
rect 21252 31578 21308 31580
rect 21012 31526 21058 31578
rect 21058 31526 21068 31578
rect 21092 31526 21122 31578
rect 21122 31526 21134 31578
rect 21134 31526 21148 31578
rect 21172 31526 21186 31578
rect 21186 31526 21198 31578
rect 21198 31526 21228 31578
rect 21252 31526 21262 31578
rect 21262 31526 21308 31578
rect 21012 31524 21068 31526
rect 21092 31524 21148 31526
rect 21172 31524 21228 31526
rect 21252 31524 21308 31526
rect 19154 26288 19210 26344
rect 18602 19896 18658 19952
rect 18878 19760 18934 19816
rect 17774 17176 17830 17232
rect 16670 14320 16726 14376
rect 17130 13640 17186 13696
rect 14312 9274 14368 9276
rect 14392 9274 14448 9276
rect 14472 9274 14528 9276
rect 14552 9274 14608 9276
rect 14312 9222 14358 9274
rect 14358 9222 14368 9274
rect 14392 9222 14422 9274
rect 14422 9222 14434 9274
rect 14434 9222 14448 9274
rect 14472 9222 14486 9274
rect 14486 9222 14498 9274
rect 14498 9222 14528 9274
rect 14552 9222 14562 9274
rect 14562 9222 14608 9274
rect 14312 9220 14368 9222
rect 14392 9220 14448 9222
rect 14472 9220 14528 9222
rect 14552 9220 14608 9222
rect 13652 8730 13708 8732
rect 13732 8730 13788 8732
rect 13812 8730 13868 8732
rect 13892 8730 13948 8732
rect 13652 8678 13698 8730
rect 13698 8678 13708 8730
rect 13732 8678 13762 8730
rect 13762 8678 13774 8730
rect 13774 8678 13788 8730
rect 13812 8678 13826 8730
rect 13826 8678 13838 8730
rect 13838 8678 13868 8730
rect 13892 8678 13902 8730
rect 13902 8678 13948 8730
rect 13652 8676 13708 8678
rect 13732 8676 13788 8678
rect 13812 8676 13868 8678
rect 13892 8676 13948 8678
rect 13266 8200 13322 8256
rect 12990 6840 13046 6896
rect 12990 5480 13046 5536
rect 13652 7642 13708 7644
rect 13732 7642 13788 7644
rect 13812 7642 13868 7644
rect 13892 7642 13948 7644
rect 13652 7590 13698 7642
rect 13698 7590 13708 7642
rect 13732 7590 13762 7642
rect 13762 7590 13774 7642
rect 13774 7590 13788 7642
rect 13812 7590 13826 7642
rect 13826 7590 13838 7642
rect 13838 7590 13868 7642
rect 13892 7590 13902 7642
rect 13902 7590 13948 7642
rect 13652 7588 13708 7590
rect 13732 7588 13788 7590
rect 13812 7588 13868 7590
rect 13892 7588 13948 7590
rect 13652 6554 13708 6556
rect 13732 6554 13788 6556
rect 13812 6554 13868 6556
rect 13892 6554 13948 6556
rect 13652 6502 13698 6554
rect 13698 6502 13708 6554
rect 13732 6502 13762 6554
rect 13762 6502 13774 6554
rect 13774 6502 13788 6554
rect 13812 6502 13826 6554
rect 13826 6502 13838 6554
rect 13838 6502 13868 6554
rect 13892 6502 13902 6554
rect 13902 6502 13948 6554
rect 13652 6500 13708 6502
rect 13732 6500 13788 6502
rect 13812 6500 13868 6502
rect 13892 6500 13948 6502
rect 13652 5466 13708 5468
rect 13732 5466 13788 5468
rect 13812 5466 13868 5468
rect 13892 5466 13948 5468
rect 13652 5414 13698 5466
rect 13698 5414 13708 5466
rect 13732 5414 13762 5466
rect 13762 5414 13774 5466
rect 13774 5414 13788 5466
rect 13812 5414 13826 5466
rect 13826 5414 13838 5466
rect 13838 5414 13868 5466
rect 13892 5414 13902 5466
rect 13902 5414 13948 5466
rect 13652 5412 13708 5414
rect 13732 5412 13788 5414
rect 13812 5412 13868 5414
rect 13892 5412 13948 5414
rect 14312 8186 14368 8188
rect 14392 8186 14448 8188
rect 14472 8186 14528 8188
rect 14552 8186 14608 8188
rect 14312 8134 14358 8186
rect 14358 8134 14368 8186
rect 14392 8134 14422 8186
rect 14422 8134 14434 8186
rect 14434 8134 14448 8186
rect 14472 8134 14486 8186
rect 14486 8134 14498 8186
rect 14498 8134 14528 8186
rect 14552 8134 14562 8186
rect 14562 8134 14608 8186
rect 14312 8132 14368 8134
rect 14392 8132 14448 8134
rect 14472 8132 14528 8134
rect 14552 8132 14608 8134
rect 13652 4378 13708 4380
rect 13732 4378 13788 4380
rect 13812 4378 13868 4380
rect 13892 4378 13948 4380
rect 13652 4326 13698 4378
rect 13698 4326 13708 4378
rect 13732 4326 13762 4378
rect 13762 4326 13774 4378
rect 13774 4326 13788 4378
rect 13812 4326 13826 4378
rect 13826 4326 13838 4378
rect 13838 4326 13868 4378
rect 13892 4326 13902 4378
rect 13902 4326 13948 4378
rect 13652 4324 13708 4326
rect 13732 4324 13788 4326
rect 13812 4324 13868 4326
rect 13892 4324 13948 4326
rect 14312 7098 14368 7100
rect 14392 7098 14448 7100
rect 14472 7098 14528 7100
rect 14552 7098 14608 7100
rect 14312 7046 14358 7098
rect 14358 7046 14368 7098
rect 14392 7046 14422 7098
rect 14422 7046 14434 7098
rect 14434 7046 14448 7098
rect 14472 7046 14486 7098
rect 14486 7046 14498 7098
rect 14498 7046 14528 7098
rect 14552 7046 14562 7098
rect 14562 7046 14608 7098
rect 14312 7044 14368 7046
rect 14392 7044 14448 7046
rect 14472 7044 14528 7046
rect 14552 7044 14608 7046
rect 14312 6010 14368 6012
rect 14392 6010 14448 6012
rect 14472 6010 14528 6012
rect 14552 6010 14608 6012
rect 14312 5958 14358 6010
rect 14358 5958 14368 6010
rect 14392 5958 14422 6010
rect 14422 5958 14434 6010
rect 14434 5958 14448 6010
rect 14472 5958 14486 6010
rect 14486 5958 14498 6010
rect 14498 5958 14528 6010
rect 14552 5958 14562 6010
rect 14562 5958 14608 6010
rect 14312 5956 14368 5958
rect 14392 5956 14448 5958
rect 14472 5956 14528 5958
rect 14552 5956 14608 5958
rect 14312 4922 14368 4924
rect 14392 4922 14448 4924
rect 14472 4922 14528 4924
rect 14552 4922 14608 4924
rect 14312 4870 14358 4922
rect 14358 4870 14368 4922
rect 14392 4870 14422 4922
rect 14422 4870 14434 4922
rect 14434 4870 14448 4922
rect 14472 4870 14486 4922
rect 14486 4870 14498 4922
rect 14498 4870 14528 4922
rect 14552 4870 14562 4922
rect 14562 4870 14608 4922
rect 14312 4868 14368 4870
rect 14392 4868 14448 4870
rect 14472 4868 14528 4870
rect 14552 4868 14608 4870
rect 13652 3290 13708 3292
rect 13732 3290 13788 3292
rect 13812 3290 13868 3292
rect 13892 3290 13948 3292
rect 13652 3238 13698 3290
rect 13698 3238 13708 3290
rect 13732 3238 13762 3290
rect 13762 3238 13774 3290
rect 13774 3238 13788 3290
rect 13812 3238 13826 3290
rect 13826 3238 13838 3290
rect 13838 3238 13868 3290
rect 13892 3238 13902 3290
rect 13902 3238 13948 3290
rect 13652 3236 13708 3238
rect 13732 3236 13788 3238
rect 13812 3236 13868 3238
rect 13892 3236 13948 3238
rect 14312 3834 14368 3836
rect 14392 3834 14448 3836
rect 14472 3834 14528 3836
rect 14552 3834 14608 3836
rect 14312 3782 14358 3834
rect 14358 3782 14368 3834
rect 14392 3782 14422 3834
rect 14422 3782 14434 3834
rect 14434 3782 14448 3834
rect 14472 3782 14486 3834
rect 14486 3782 14498 3834
rect 14498 3782 14528 3834
rect 14552 3782 14562 3834
rect 14562 3782 14608 3834
rect 14312 3780 14368 3782
rect 14392 3780 14448 3782
rect 14472 3780 14528 3782
rect 14552 3780 14608 3782
rect 15290 6296 15346 6352
rect 15750 5228 15806 5264
rect 15750 5208 15752 5228
rect 15752 5208 15804 5228
rect 15804 5208 15806 5228
rect 14312 2746 14368 2748
rect 14392 2746 14448 2748
rect 14472 2746 14528 2748
rect 14552 2746 14608 2748
rect 14312 2694 14358 2746
rect 14358 2694 14368 2746
rect 14392 2694 14422 2746
rect 14422 2694 14434 2746
rect 14434 2694 14448 2746
rect 14472 2694 14486 2746
rect 14486 2694 14498 2746
rect 14498 2694 14528 2746
rect 14552 2694 14562 2746
rect 14562 2694 14608 2746
rect 14312 2692 14368 2694
rect 14392 2692 14448 2694
rect 14472 2692 14528 2694
rect 14552 2692 14608 2694
rect 21012 30490 21068 30492
rect 21092 30490 21148 30492
rect 21172 30490 21228 30492
rect 21252 30490 21308 30492
rect 21012 30438 21058 30490
rect 21058 30438 21068 30490
rect 21092 30438 21122 30490
rect 21122 30438 21134 30490
rect 21134 30438 21148 30490
rect 21172 30438 21186 30490
rect 21186 30438 21198 30490
rect 21198 30438 21228 30490
rect 21252 30438 21262 30490
rect 21262 30438 21308 30490
rect 21012 30436 21068 30438
rect 21092 30436 21148 30438
rect 21172 30436 21228 30438
rect 21252 30436 21308 30438
rect 21672 32122 21728 32124
rect 21752 32122 21808 32124
rect 21832 32122 21888 32124
rect 21912 32122 21968 32124
rect 21672 32070 21718 32122
rect 21718 32070 21728 32122
rect 21752 32070 21782 32122
rect 21782 32070 21794 32122
rect 21794 32070 21808 32122
rect 21832 32070 21846 32122
rect 21846 32070 21858 32122
rect 21858 32070 21888 32122
rect 21912 32070 21922 32122
rect 21922 32070 21968 32122
rect 21672 32068 21728 32070
rect 21752 32068 21808 32070
rect 21832 32068 21888 32070
rect 21912 32068 21968 32070
rect 21672 31034 21728 31036
rect 21752 31034 21808 31036
rect 21832 31034 21888 31036
rect 21912 31034 21968 31036
rect 21672 30982 21718 31034
rect 21718 30982 21728 31034
rect 21752 30982 21782 31034
rect 21782 30982 21794 31034
rect 21794 30982 21808 31034
rect 21832 30982 21846 31034
rect 21846 30982 21858 31034
rect 21858 30982 21888 31034
rect 21912 30982 21922 31034
rect 21922 30982 21968 31034
rect 21672 30980 21728 30982
rect 21752 30980 21808 30982
rect 21832 30980 21888 30982
rect 21912 30980 21968 30982
rect 21672 29946 21728 29948
rect 21752 29946 21808 29948
rect 21832 29946 21888 29948
rect 21912 29946 21968 29948
rect 21672 29894 21718 29946
rect 21718 29894 21728 29946
rect 21752 29894 21782 29946
rect 21782 29894 21794 29946
rect 21794 29894 21808 29946
rect 21832 29894 21846 29946
rect 21846 29894 21858 29946
rect 21858 29894 21888 29946
rect 21912 29894 21922 29946
rect 21922 29894 21968 29946
rect 21672 29892 21728 29894
rect 21752 29892 21808 29894
rect 21832 29892 21888 29894
rect 21912 29892 21968 29894
rect 21012 29402 21068 29404
rect 21092 29402 21148 29404
rect 21172 29402 21228 29404
rect 21252 29402 21308 29404
rect 21012 29350 21058 29402
rect 21058 29350 21068 29402
rect 21092 29350 21122 29402
rect 21122 29350 21134 29402
rect 21134 29350 21148 29402
rect 21172 29350 21186 29402
rect 21186 29350 21198 29402
rect 21198 29350 21228 29402
rect 21252 29350 21262 29402
rect 21262 29350 21308 29402
rect 21012 29348 21068 29350
rect 21092 29348 21148 29350
rect 21172 29348 21228 29350
rect 21252 29348 21308 29350
rect 21672 28858 21728 28860
rect 21752 28858 21808 28860
rect 21832 28858 21888 28860
rect 21912 28858 21968 28860
rect 21672 28806 21718 28858
rect 21718 28806 21728 28858
rect 21752 28806 21782 28858
rect 21782 28806 21794 28858
rect 21794 28806 21808 28858
rect 21832 28806 21846 28858
rect 21846 28806 21858 28858
rect 21858 28806 21888 28858
rect 21912 28806 21922 28858
rect 21922 28806 21968 28858
rect 21672 28804 21728 28806
rect 21752 28804 21808 28806
rect 21832 28804 21888 28806
rect 21912 28804 21968 28806
rect 21012 28314 21068 28316
rect 21092 28314 21148 28316
rect 21172 28314 21228 28316
rect 21252 28314 21308 28316
rect 21012 28262 21058 28314
rect 21058 28262 21068 28314
rect 21092 28262 21122 28314
rect 21122 28262 21134 28314
rect 21134 28262 21148 28314
rect 21172 28262 21186 28314
rect 21186 28262 21198 28314
rect 21198 28262 21228 28314
rect 21252 28262 21262 28314
rect 21262 28262 21308 28314
rect 21012 28260 21068 28262
rect 21092 28260 21148 28262
rect 21172 28260 21228 28262
rect 21252 28260 21308 28262
rect 21012 27226 21068 27228
rect 21092 27226 21148 27228
rect 21172 27226 21228 27228
rect 21252 27226 21308 27228
rect 21012 27174 21058 27226
rect 21058 27174 21068 27226
rect 21092 27174 21122 27226
rect 21122 27174 21134 27226
rect 21134 27174 21148 27226
rect 21172 27174 21186 27226
rect 21186 27174 21198 27226
rect 21198 27174 21228 27226
rect 21252 27174 21262 27226
rect 21262 27174 21308 27226
rect 21012 27172 21068 27174
rect 21092 27172 21148 27174
rect 21172 27172 21228 27174
rect 21252 27172 21308 27174
rect 21672 27770 21728 27772
rect 21752 27770 21808 27772
rect 21832 27770 21888 27772
rect 21912 27770 21968 27772
rect 21672 27718 21718 27770
rect 21718 27718 21728 27770
rect 21752 27718 21782 27770
rect 21782 27718 21794 27770
rect 21794 27718 21808 27770
rect 21832 27718 21846 27770
rect 21846 27718 21858 27770
rect 21858 27718 21888 27770
rect 21912 27718 21922 27770
rect 21922 27718 21968 27770
rect 21672 27716 21728 27718
rect 21752 27716 21808 27718
rect 21832 27716 21888 27718
rect 21912 27716 21968 27718
rect 19062 17992 19118 18048
rect 18970 17856 19026 17912
rect 18878 17720 18934 17776
rect 19614 18400 19670 18456
rect 19522 18264 19578 18320
rect 18326 17040 18382 17096
rect 21672 26682 21728 26684
rect 21752 26682 21808 26684
rect 21832 26682 21888 26684
rect 21912 26682 21968 26684
rect 21672 26630 21718 26682
rect 21718 26630 21728 26682
rect 21752 26630 21782 26682
rect 21782 26630 21794 26682
rect 21794 26630 21808 26682
rect 21832 26630 21846 26682
rect 21846 26630 21858 26682
rect 21858 26630 21888 26682
rect 21912 26630 21922 26682
rect 21922 26630 21968 26682
rect 21672 26628 21728 26630
rect 21752 26628 21808 26630
rect 21832 26628 21888 26630
rect 21912 26628 21968 26630
rect 21012 26138 21068 26140
rect 21092 26138 21148 26140
rect 21172 26138 21228 26140
rect 21252 26138 21308 26140
rect 21012 26086 21058 26138
rect 21058 26086 21068 26138
rect 21092 26086 21122 26138
rect 21122 26086 21134 26138
rect 21134 26086 21148 26138
rect 21172 26086 21186 26138
rect 21186 26086 21198 26138
rect 21198 26086 21228 26138
rect 21252 26086 21262 26138
rect 21262 26086 21308 26138
rect 21012 26084 21068 26086
rect 21092 26084 21148 26086
rect 21172 26084 21228 26086
rect 21252 26084 21308 26086
rect 21012 25050 21068 25052
rect 21092 25050 21148 25052
rect 21172 25050 21228 25052
rect 21252 25050 21308 25052
rect 21012 24998 21058 25050
rect 21058 24998 21068 25050
rect 21092 24998 21122 25050
rect 21122 24998 21134 25050
rect 21134 24998 21148 25050
rect 21172 24998 21186 25050
rect 21186 24998 21198 25050
rect 21198 24998 21228 25050
rect 21252 24998 21262 25050
rect 21262 24998 21308 25050
rect 21012 24996 21068 24998
rect 21092 24996 21148 24998
rect 21172 24996 21228 24998
rect 21252 24996 21308 24998
rect 21672 25594 21728 25596
rect 21752 25594 21808 25596
rect 21832 25594 21888 25596
rect 21912 25594 21968 25596
rect 21672 25542 21718 25594
rect 21718 25542 21728 25594
rect 21752 25542 21782 25594
rect 21782 25542 21794 25594
rect 21794 25542 21808 25594
rect 21832 25542 21846 25594
rect 21846 25542 21858 25594
rect 21858 25542 21888 25594
rect 21912 25542 21922 25594
rect 21922 25542 21968 25594
rect 21672 25540 21728 25542
rect 21752 25540 21808 25542
rect 21832 25540 21888 25542
rect 21912 25540 21968 25542
rect 21672 24506 21728 24508
rect 21752 24506 21808 24508
rect 21832 24506 21888 24508
rect 21912 24506 21968 24508
rect 21672 24454 21718 24506
rect 21718 24454 21728 24506
rect 21752 24454 21782 24506
rect 21782 24454 21794 24506
rect 21794 24454 21808 24506
rect 21832 24454 21846 24506
rect 21846 24454 21858 24506
rect 21858 24454 21888 24506
rect 21912 24454 21922 24506
rect 21922 24454 21968 24506
rect 21672 24452 21728 24454
rect 21752 24452 21808 24454
rect 21832 24452 21888 24454
rect 21912 24452 21968 24454
rect 21012 23962 21068 23964
rect 21092 23962 21148 23964
rect 21172 23962 21228 23964
rect 21252 23962 21308 23964
rect 21012 23910 21058 23962
rect 21058 23910 21068 23962
rect 21092 23910 21122 23962
rect 21122 23910 21134 23962
rect 21134 23910 21148 23962
rect 21172 23910 21186 23962
rect 21186 23910 21198 23962
rect 21198 23910 21228 23962
rect 21252 23910 21262 23962
rect 21262 23910 21308 23962
rect 21012 23908 21068 23910
rect 21092 23908 21148 23910
rect 21172 23908 21228 23910
rect 21252 23908 21308 23910
rect 21012 22874 21068 22876
rect 21092 22874 21148 22876
rect 21172 22874 21228 22876
rect 21252 22874 21308 22876
rect 21012 22822 21058 22874
rect 21058 22822 21068 22874
rect 21092 22822 21122 22874
rect 21122 22822 21134 22874
rect 21134 22822 21148 22874
rect 21172 22822 21186 22874
rect 21186 22822 21198 22874
rect 21198 22822 21228 22874
rect 21252 22822 21262 22874
rect 21262 22822 21308 22874
rect 21012 22820 21068 22822
rect 21092 22820 21148 22822
rect 21172 22820 21228 22822
rect 21252 22820 21308 22822
rect 21672 23418 21728 23420
rect 21752 23418 21808 23420
rect 21832 23418 21888 23420
rect 21912 23418 21968 23420
rect 21672 23366 21718 23418
rect 21718 23366 21728 23418
rect 21752 23366 21782 23418
rect 21782 23366 21794 23418
rect 21794 23366 21808 23418
rect 21832 23366 21846 23418
rect 21846 23366 21858 23418
rect 21858 23366 21888 23418
rect 21912 23366 21922 23418
rect 21922 23366 21968 23418
rect 21672 23364 21728 23366
rect 21752 23364 21808 23366
rect 21832 23364 21888 23366
rect 21912 23364 21968 23366
rect 21546 22616 21602 22672
rect 21012 21786 21068 21788
rect 21092 21786 21148 21788
rect 21172 21786 21228 21788
rect 21252 21786 21308 21788
rect 21012 21734 21058 21786
rect 21058 21734 21068 21786
rect 21092 21734 21122 21786
rect 21122 21734 21134 21786
rect 21134 21734 21148 21786
rect 21172 21734 21186 21786
rect 21186 21734 21198 21786
rect 21198 21734 21228 21786
rect 21252 21734 21262 21786
rect 21262 21734 21308 21786
rect 21012 21732 21068 21734
rect 21092 21732 21148 21734
rect 21172 21732 21228 21734
rect 21252 21732 21308 21734
rect 23570 26968 23626 27024
rect 24490 31048 24546 31104
rect 25226 31084 25228 31104
rect 25228 31084 25280 31104
rect 25280 31084 25282 31104
rect 25226 31048 25282 31084
rect 25594 31048 25650 31104
rect 25778 30096 25834 30152
rect 26606 31084 26608 31104
rect 26608 31084 26660 31104
rect 26660 31084 26662 31104
rect 26606 31048 26662 31084
rect 26146 28600 26202 28656
rect 24398 26968 24454 27024
rect 21638 22480 21694 22536
rect 21672 22330 21728 22332
rect 21752 22330 21808 22332
rect 21832 22330 21888 22332
rect 21912 22330 21968 22332
rect 21672 22278 21718 22330
rect 21718 22278 21728 22330
rect 21752 22278 21782 22330
rect 21782 22278 21794 22330
rect 21794 22278 21808 22330
rect 21832 22278 21846 22330
rect 21846 22278 21858 22330
rect 21858 22278 21888 22330
rect 21912 22278 21922 22330
rect 21922 22278 21968 22330
rect 21672 22276 21728 22278
rect 21752 22276 21808 22278
rect 21832 22276 21888 22278
rect 21912 22276 21968 22278
rect 21672 21242 21728 21244
rect 21752 21242 21808 21244
rect 21832 21242 21888 21244
rect 21912 21242 21968 21244
rect 21672 21190 21718 21242
rect 21718 21190 21728 21242
rect 21752 21190 21782 21242
rect 21782 21190 21794 21242
rect 21794 21190 21808 21242
rect 21832 21190 21846 21242
rect 21846 21190 21858 21242
rect 21858 21190 21888 21242
rect 21912 21190 21922 21242
rect 21922 21190 21968 21242
rect 21672 21188 21728 21190
rect 21752 21188 21808 21190
rect 21832 21188 21888 21190
rect 21912 21188 21968 21190
rect 20442 20304 20498 20360
rect 20442 18264 20498 18320
rect 19798 18164 19800 18184
rect 19800 18164 19852 18184
rect 19852 18164 19854 18184
rect 19798 18128 19854 18164
rect 20074 14220 20076 14240
rect 20076 14220 20128 14240
rect 20128 14220 20130 14240
rect 20074 14184 20130 14220
rect 21012 20698 21068 20700
rect 21092 20698 21148 20700
rect 21172 20698 21228 20700
rect 21252 20698 21308 20700
rect 21012 20646 21058 20698
rect 21058 20646 21068 20698
rect 21092 20646 21122 20698
rect 21122 20646 21134 20698
rect 21134 20646 21148 20698
rect 21172 20646 21186 20698
rect 21186 20646 21198 20698
rect 21198 20646 21228 20698
rect 21252 20646 21262 20698
rect 21262 20646 21308 20698
rect 21012 20644 21068 20646
rect 21092 20644 21148 20646
rect 21172 20644 21228 20646
rect 21252 20644 21308 20646
rect 20902 20440 20958 20496
rect 21012 19610 21068 19612
rect 21092 19610 21148 19612
rect 21172 19610 21228 19612
rect 21252 19610 21308 19612
rect 21012 19558 21058 19610
rect 21058 19558 21068 19610
rect 21092 19558 21122 19610
rect 21122 19558 21134 19610
rect 21134 19558 21148 19610
rect 21172 19558 21186 19610
rect 21186 19558 21198 19610
rect 21198 19558 21228 19610
rect 21252 19558 21262 19610
rect 21262 19558 21308 19610
rect 21012 19556 21068 19558
rect 21092 19556 21148 19558
rect 21172 19556 21228 19558
rect 21252 19556 21308 19558
rect 21672 20154 21728 20156
rect 21752 20154 21808 20156
rect 21832 20154 21888 20156
rect 21912 20154 21968 20156
rect 21672 20102 21718 20154
rect 21718 20102 21728 20154
rect 21752 20102 21782 20154
rect 21782 20102 21794 20154
rect 21794 20102 21808 20154
rect 21832 20102 21846 20154
rect 21846 20102 21858 20154
rect 21858 20102 21888 20154
rect 21912 20102 21922 20154
rect 21922 20102 21968 20154
rect 21672 20100 21728 20102
rect 21752 20100 21808 20102
rect 21832 20100 21888 20102
rect 21912 20100 21968 20102
rect 21672 19066 21728 19068
rect 21752 19066 21808 19068
rect 21832 19066 21888 19068
rect 21912 19066 21968 19068
rect 21672 19014 21718 19066
rect 21718 19014 21728 19066
rect 21752 19014 21782 19066
rect 21782 19014 21794 19066
rect 21794 19014 21808 19066
rect 21832 19014 21846 19066
rect 21846 19014 21858 19066
rect 21858 19014 21888 19066
rect 21912 19014 21922 19066
rect 21922 19014 21968 19066
rect 21672 19012 21728 19014
rect 21752 19012 21808 19014
rect 21832 19012 21888 19014
rect 21912 19012 21968 19014
rect 21362 18808 21418 18864
rect 21362 18672 21418 18728
rect 21012 18522 21068 18524
rect 21092 18522 21148 18524
rect 21172 18522 21228 18524
rect 21252 18522 21308 18524
rect 21012 18470 21058 18522
rect 21058 18470 21068 18522
rect 21092 18470 21122 18522
rect 21122 18470 21134 18522
rect 21134 18470 21148 18522
rect 21172 18470 21186 18522
rect 21186 18470 21198 18522
rect 21198 18470 21228 18522
rect 21252 18470 21262 18522
rect 21262 18470 21308 18522
rect 21012 18468 21068 18470
rect 21092 18468 21148 18470
rect 21172 18468 21228 18470
rect 21252 18468 21308 18470
rect 20810 18400 20866 18456
rect 20626 18128 20682 18184
rect 21012 17434 21068 17436
rect 21092 17434 21148 17436
rect 21172 17434 21228 17436
rect 21252 17434 21308 17436
rect 21012 17382 21058 17434
rect 21058 17382 21068 17434
rect 21092 17382 21122 17434
rect 21122 17382 21134 17434
rect 21134 17382 21148 17434
rect 21172 17382 21186 17434
rect 21186 17382 21198 17434
rect 21198 17382 21228 17434
rect 21252 17382 21262 17434
rect 21262 17382 21308 17434
rect 21012 17380 21068 17382
rect 21092 17380 21148 17382
rect 21172 17380 21228 17382
rect 21252 17380 21308 17382
rect 21672 17978 21728 17980
rect 21752 17978 21808 17980
rect 21832 17978 21888 17980
rect 21912 17978 21968 17980
rect 21672 17926 21718 17978
rect 21718 17926 21728 17978
rect 21752 17926 21782 17978
rect 21782 17926 21794 17978
rect 21794 17926 21808 17978
rect 21832 17926 21846 17978
rect 21846 17926 21858 17978
rect 21858 17926 21888 17978
rect 21912 17926 21922 17978
rect 21922 17926 21968 17978
rect 21672 17924 21728 17926
rect 21752 17924 21808 17926
rect 21832 17924 21888 17926
rect 21912 17924 21968 17926
rect 24582 23296 24638 23352
rect 25778 27004 25780 27024
rect 25780 27004 25832 27024
rect 25832 27004 25834 27024
rect 25778 26968 25834 27004
rect 24674 22108 24676 22128
rect 24676 22108 24728 22128
rect 24728 22108 24730 22128
rect 24674 22072 24730 22108
rect 23754 19624 23810 19680
rect 21672 16890 21728 16892
rect 21752 16890 21808 16892
rect 21832 16890 21888 16892
rect 21912 16890 21968 16892
rect 21672 16838 21718 16890
rect 21718 16838 21728 16890
rect 21752 16838 21782 16890
rect 21782 16838 21794 16890
rect 21794 16838 21808 16890
rect 21832 16838 21846 16890
rect 21846 16838 21858 16890
rect 21858 16838 21888 16890
rect 21912 16838 21922 16890
rect 21922 16838 21968 16890
rect 21672 16836 21728 16838
rect 21752 16836 21808 16838
rect 21832 16836 21888 16838
rect 21912 16836 21968 16838
rect 24398 20304 24454 20360
rect 25502 23568 25558 23624
rect 25318 22344 25374 22400
rect 26974 30096 27030 30152
rect 29032 32122 29088 32124
rect 29112 32122 29168 32124
rect 29192 32122 29248 32124
rect 29272 32122 29328 32124
rect 29032 32070 29078 32122
rect 29078 32070 29088 32122
rect 29112 32070 29142 32122
rect 29142 32070 29154 32122
rect 29154 32070 29168 32122
rect 29192 32070 29206 32122
rect 29206 32070 29218 32122
rect 29218 32070 29248 32122
rect 29272 32070 29282 32122
rect 29282 32070 29328 32122
rect 29032 32068 29088 32070
rect 29112 32068 29168 32070
rect 29192 32068 29248 32070
rect 29272 32068 29328 32070
rect 28372 31578 28428 31580
rect 28452 31578 28508 31580
rect 28532 31578 28588 31580
rect 28612 31578 28668 31580
rect 28372 31526 28418 31578
rect 28418 31526 28428 31578
rect 28452 31526 28482 31578
rect 28482 31526 28494 31578
rect 28494 31526 28508 31578
rect 28532 31526 28546 31578
rect 28546 31526 28558 31578
rect 28558 31526 28588 31578
rect 28612 31526 28622 31578
rect 28622 31526 28668 31578
rect 28372 31524 28428 31526
rect 28452 31524 28508 31526
rect 28532 31524 28588 31526
rect 28612 31524 28668 31526
rect 29642 31320 29698 31376
rect 29032 31034 29088 31036
rect 29112 31034 29168 31036
rect 29192 31034 29248 31036
rect 29272 31034 29328 31036
rect 29032 30982 29078 31034
rect 29078 30982 29088 31034
rect 29112 30982 29142 31034
rect 29142 30982 29154 31034
rect 29154 30982 29168 31034
rect 29192 30982 29206 31034
rect 29206 30982 29218 31034
rect 29218 30982 29248 31034
rect 29272 30982 29282 31034
rect 29282 30982 29328 31034
rect 29032 30980 29088 30982
rect 29112 30980 29168 30982
rect 29192 30980 29248 30982
rect 29272 30980 29328 30982
rect 28372 30490 28428 30492
rect 28452 30490 28508 30492
rect 28532 30490 28588 30492
rect 28612 30490 28668 30492
rect 28372 30438 28418 30490
rect 28418 30438 28428 30490
rect 28452 30438 28482 30490
rect 28482 30438 28494 30490
rect 28494 30438 28508 30490
rect 28532 30438 28546 30490
rect 28546 30438 28558 30490
rect 28558 30438 28588 30490
rect 28612 30438 28622 30490
rect 28622 30438 28668 30490
rect 28372 30436 28428 30438
rect 28452 30436 28508 30438
rect 28532 30436 28588 30438
rect 28612 30436 28668 30438
rect 28372 29402 28428 29404
rect 28452 29402 28508 29404
rect 28532 29402 28588 29404
rect 28612 29402 28668 29404
rect 28372 29350 28418 29402
rect 28418 29350 28428 29402
rect 28452 29350 28482 29402
rect 28482 29350 28494 29402
rect 28494 29350 28508 29402
rect 28532 29350 28546 29402
rect 28546 29350 28558 29402
rect 28558 29350 28588 29402
rect 28612 29350 28622 29402
rect 28622 29350 28668 29402
rect 28372 29348 28428 29350
rect 28452 29348 28508 29350
rect 28532 29348 28588 29350
rect 28612 29348 28668 29350
rect 29032 29946 29088 29948
rect 29112 29946 29168 29948
rect 29192 29946 29248 29948
rect 29272 29946 29328 29948
rect 29032 29894 29078 29946
rect 29078 29894 29088 29946
rect 29112 29894 29142 29946
rect 29142 29894 29154 29946
rect 29154 29894 29168 29946
rect 29192 29894 29206 29946
rect 29206 29894 29218 29946
rect 29218 29894 29248 29946
rect 29272 29894 29282 29946
rect 29282 29894 29328 29946
rect 29032 29892 29088 29894
rect 29112 29892 29168 29894
rect 29192 29892 29248 29894
rect 29272 29892 29328 29894
rect 27526 26968 27582 27024
rect 28372 28314 28428 28316
rect 28452 28314 28508 28316
rect 28532 28314 28588 28316
rect 28612 28314 28668 28316
rect 28372 28262 28418 28314
rect 28418 28262 28428 28314
rect 28452 28262 28482 28314
rect 28482 28262 28494 28314
rect 28494 28262 28508 28314
rect 28532 28262 28546 28314
rect 28546 28262 28558 28314
rect 28558 28262 28588 28314
rect 28612 28262 28622 28314
rect 28622 28262 28668 28314
rect 28372 28260 28428 28262
rect 28452 28260 28508 28262
rect 28532 28260 28588 28262
rect 28612 28260 28668 28262
rect 29032 28858 29088 28860
rect 29112 28858 29168 28860
rect 29192 28858 29248 28860
rect 29272 28858 29328 28860
rect 29032 28806 29078 28858
rect 29078 28806 29088 28858
rect 29112 28806 29142 28858
rect 29142 28806 29154 28858
rect 29154 28806 29168 28858
rect 29192 28806 29206 28858
rect 29206 28806 29218 28858
rect 29218 28806 29248 28858
rect 29272 28806 29282 28858
rect 29282 28806 29328 28858
rect 29032 28804 29088 28806
rect 29112 28804 29168 28806
rect 29192 28804 29248 28806
rect 29272 28804 29328 28806
rect 28906 28600 28962 28656
rect 26054 23296 26110 23352
rect 26054 22616 26110 22672
rect 29458 28056 29514 28112
rect 29366 27920 29422 27976
rect 29032 27770 29088 27772
rect 29112 27770 29168 27772
rect 29192 27770 29248 27772
rect 29272 27770 29328 27772
rect 29032 27718 29078 27770
rect 29078 27718 29088 27770
rect 29112 27718 29142 27770
rect 29142 27718 29154 27770
rect 29154 27718 29168 27770
rect 29192 27718 29206 27770
rect 29206 27718 29218 27770
rect 29218 27718 29248 27770
rect 29272 27718 29282 27770
rect 29282 27718 29328 27770
rect 29032 27716 29088 27718
rect 29112 27716 29168 27718
rect 29192 27716 29248 27718
rect 29272 27716 29328 27718
rect 28372 27226 28428 27228
rect 28452 27226 28508 27228
rect 28532 27226 28588 27228
rect 28612 27226 28668 27228
rect 28372 27174 28418 27226
rect 28418 27174 28428 27226
rect 28452 27174 28482 27226
rect 28482 27174 28494 27226
rect 28494 27174 28508 27226
rect 28532 27174 28546 27226
rect 28546 27174 28558 27226
rect 28558 27174 28588 27226
rect 28612 27174 28622 27226
rect 28622 27174 28668 27226
rect 28372 27172 28428 27174
rect 28452 27172 28508 27174
rect 28532 27172 28588 27174
rect 28612 27172 28668 27174
rect 29550 27396 29606 27432
rect 29550 27376 29552 27396
rect 29552 27376 29604 27396
rect 29604 27376 29606 27396
rect 29032 26682 29088 26684
rect 29112 26682 29168 26684
rect 29192 26682 29248 26684
rect 29272 26682 29328 26684
rect 29032 26630 29078 26682
rect 29078 26630 29088 26682
rect 29112 26630 29142 26682
rect 29142 26630 29154 26682
rect 29154 26630 29168 26682
rect 29192 26630 29206 26682
rect 29206 26630 29218 26682
rect 29218 26630 29248 26682
rect 29272 26630 29282 26682
rect 29282 26630 29328 26682
rect 29032 26628 29088 26630
rect 29112 26628 29168 26630
rect 29192 26628 29248 26630
rect 29272 26628 29328 26630
rect 28372 26138 28428 26140
rect 28452 26138 28508 26140
rect 28532 26138 28588 26140
rect 28612 26138 28668 26140
rect 28372 26086 28418 26138
rect 28418 26086 28428 26138
rect 28452 26086 28482 26138
rect 28482 26086 28494 26138
rect 28494 26086 28508 26138
rect 28532 26086 28546 26138
rect 28546 26086 28558 26138
rect 28558 26086 28588 26138
rect 28612 26086 28622 26138
rect 28622 26086 28668 26138
rect 28372 26084 28428 26086
rect 28452 26084 28508 26086
rect 28532 26084 28588 26086
rect 28612 26084 28668 26086
rect 29032 25594 29088 25596
rect 29112 25594 29168 25596
rect 29192 25594 29248 25596
rect 29272 25594 29328 25596
rect 29032 25542 29078 25594
rect 29078 25542 29088 25594
rect 29112 25542 29142 25594
rect 29142 25542 29154 25594
rect 29154 25542 29168 25594
rect 29192 25542 29206 25594
rect 29206 25542 29218 25594
rect 29218 25542 29248 25594
rect 29272 25542 29282 25594
rect 29282 25542 29328 25594
rect 29032 25540 29088 25542
rect 29112 25540 29168 25542
rect 29192 25540 29248 25542
rect 29272 25540 29328 25542
rect 28372 25050 28428 25052
rect 28452 25050 28508 25052
rect 28532 25050 28588 25052
rect 28612 25050 28668 25052
rect 28372 24998 28418 25050
rect 28418 24998 28428 25050
rect 28452 24998 28482 25050
rect 28482 24998 28494 25050
rect 28494 24998 28508 25050
rect 28532 24998 28546 25050
rect 28546 24998 28558 25050
rect 28558 24998 28588 25050
rect 28612 24998 28622 25050
rect 28622 24998 28668 25050
rect 28372 24996 28428 24998
rect 28452 24996 28508 24998
rect 28532 24996 28588 24998
rect 28612 24996 28668 24998
rect 26790 23568 26846 23624
rect 25318 19624 25374 19680
rect 27250 23296 27306 23352
rect 26698 22480 26754 22536
rect 26974 22344 27030 22400
rect 27434 22480 27490 22536
rect 27342 22108 27344 22128
rect 27344 22108 27396 22128
rect 27396 22108 27398 22128
rect 27342 22072 27398 22108
rect 26882 18808 26938 18864
rect 29032 24506 29088 24508
rect 29112 24506 29168 24508
rect 29192 24506 29248 24508
rect 29272 24506 29328 24508
rect 29032 24454 29078 24506
rect 29078 24454 29088 24506
rect 29112 24454 29142 24506
rect 29142 24454 29154 24506
rect 29154 24454 29168 24506
rect 29192 24454 29206 24506
rect 29206 24454 29218 24506
rect 29218 24454 29248 24506
rect 29272 24454 29282 24506
rect 29282 24454 29328 24506
rect 29032 24452 29088 24454
rect 29112 24452 29168 24454
rect 29192 24452 29248 24454
rect 29272 24452 29328 24454
rect 28372 23962 28428 23964
rect 28452 23962 28508 23964
rect 28532 23962 28588 23964
rect 28612 23962 28668 23964
rect 28372 23910 28418 23962
rect 28418 23910 28428 23962
rect 28452 23910 28482 23962
rect 28482 23910 28494 23962
rect 28494 23910 28508 23962
rect 28532 23910 28546 23962
rect 28546 23910 28558 23962
rect 28558 23910 28588 23962
rect 28612 23910 28622 23962
rect 28622 23910 28668 23962
rect 28372 23908 28428 23910
rect 28452 23908 28508 23910
rect 28532 23908 28588 23910
rect 28612 23908 28668 23910
rect 28372 22874 28428 22876
rect 28452 22874 28508 22876
rect 28532 22874 28588 22876
rect 28612 22874 28668 22876
rect 28372 22822 28418 22874
rect 28418 22822 28428 22874
rect 28452 22822 28482 22874
rect 28482 22822 28494 22874
rect 28494 22822 28508 22874
rect 28532 22822 28546 22874
rect 28546 22822 28558 22874
rect 28558 22822 28588 22874
rect 28612 22822 28622 22874
rect 28622 22822 28668 22874
rect 28372 22820 28428 22822
rect 28452 22820 28508 22822
rect 28532 22820 28588 22822
rect 28612 22820 28668 22822
rect 28372 21786 28428 21788
rect 28452 21786 28508 21788
rect 28532 21786 28588 21788
rect 28612 21786 28668 21788
rect 28372 21734 28418 21786
rect 28418 21734 28428 21786
rect 28452 21734 28482 21786
rect 28482 21734 28494 21786
rect 28494 21734 28508 21786
rect 28532 21734 28546 21786
rect 28546 21734 28558 21786
rect 28558 21734 28588 21786
rect 28612 21734 28622 21786
rect 28622 21734 28668 21786
rect 28372 21732 28428 21734
rect 28452 21732 28508 21734
rect 28532 21732 28588 21734
rect 28612 21732 28668 21734
rect 29032 23418 29088 23420
rect 29112 23418 29168 23420
rect 29192 23418 29248 23420
rect 29272 23418 29328 23420
rect 29032 23366 29078 23418
rect 29078 23366 29088 23418
rect 29112 23366 29142 23418
rect 29142 23366 29154 23418
rect 29154 23366 29168 23418
rect 29192 23366 29206 23418
rect 29206 23366 29218 23418
rect 29218 23366 29248 23418
rect 29272 23366 29282 23418
rect 29282 23366 29328 23418
rect 29032 23364 29088 23366
rect 29112 23364 29168 23366
rect 29192 23364 29248 23366
rect 29272 23364 29328 23366
rect 30378 28600 30434 28656
rect 30194 28076 30250 28112
rect 30194 28056 30196 28076
rect 30196 28056 30248 28076
rect 30248 28056 30250 28076
rect 30746 27920 30802 27976
rect 30102 27376 30158 27432
rect 29032 22330 29088 22332
rect 29112 22330 29168 22332
rect 29192 22330 29248 22332
rect 29272 22330 29328 22332
rect 29032 22278 29078 22330
rect 29078 22278 29088 22330
rect 29112 22278 29142 22330
rect 29142 22278 29154 22330
rect 29154 22278 29168 22330
rect 29192 22278 29206 22330
rect 29206 22278 29218 22330
rect 29218 22278 29248 22330
rect 29272 22278 29282 22330
rect 29282 22278 29328 22330
rect 29032 22276 29088 22278
rect 29112 22276 29168 22278
rect 29192 22276 29248 22278
rect 29272 22276 29328 22278
rect 28372 20698 28428 20700
rect 28452 20698 28508 20700
rect 28532 20698 28588 20700
rect 28612 20698 28668 20700
rect 28372 20646 28418 20698
rect 28418 20646 28428 20698
rect 28452 20646 28482 20698
rect 28482 20646 28494 20698
rect 28494 20646 28508 20698
rect 28532 20646 28546 20698
rect 28546 20646 28558 20698
rect 28558 20646 28588 20698
rect 28612 20646 28622 20698
rect 28622 20646 28668 20698
rect 28372 20644 28428 20646
rect 28452 20644 28508 20646
rect 28532 20644 28588 20646
rect 28612 20644 28668 20646
rect 28078 20440 28134 20496
rect 29032 21242 29088 21244
rect 29112 21242 29168 21244
rect 29192 21242 29248 21244
rect 29272 21242 29328 21244
rect 29032 21190 29078 21242
rect 29078 21190 29088 21242
rect 29112 21190 29142 21242
rect 29142 21190 29154 21242
rect 29154 21190 29168 21242
rect 29192 21190 29206 21242
rect 29206 21190 29218 21242
rect 29218 21190 29248 21242
rect 29272 21190 29282 21242
rect 29282 21190 29328 21242
rect 29032 21188 29088 21190
rect 29112 21188 29168 21190
rect 29192 21188 29248 21190
rect 29272 21188 29328 21190
rect 29734 20984 29790 21040
rect 29032 20154 29088 20156
rect 29112 20154 29168 20156
rect 29192 20154 29248 20156
rect 29272 20154 29328 20156
rect 29032 20102 29078 20154
rect 29078 20102 29088 20154
rect 29112 20102 29142 20154
rect 29142 20102 29154 20154
rect 29154 20102 29168 20154
rect 29192 20102 29206 20154
rect 29206 20102 29218 20154
rect 29218 20102 29248 20154
rect 29272 20102 29282 20154
rect 29282 20102 29328 20154
rect 29032 20100 29088 20102
rect 29112 20100 29168 20102
rect 29192 20100 29248 20102
rect 29272 20100 29328 20102
rect 28372 19610 28428 19612
rect 28452 19610 28508 19612
rect 28532 19610 28588 19612
rect 28612 19610 28668 19612
rect 28372 19558 28418 19610
rect 28418 19558 28428 19610
rect 28452 19558 28482 19610
rect 28482 19558 28494 19610
rect 28494 19558 28508 19610
rect 28532 19558 28546 19610
rect 28546 19558 28558 19610
rect 28558 19558 28588 19610
rect 28612 19558 28622 19610
rect 28622 19558 28668 19610
rect 28372 19556 28428 19558
rect 28452 19556 28508 19558
rect 28532 19556 28588 19558
rect 28612 19556 28668 19558
rect 29032 19066 29088 19068
rect 29112 19066 29168 19068
rect 29192 19066 29248 19068
rect 29272 19066 29328 19068
rect 29032 19014 29078 19066
rect 29078 19014 29088 19066
rect 29112 19014 29142 19066
rect 29142 19014 29154 19066
rect 29154 19014 29168 19066
rect 29192 19014 29206 19066
rect 29206 19014 29218 19066
rect 29218 19014 29248 19066
rect 29272 19014 29282 19066
rect 29282 19014 29328 19066
rect 29032 19012 29088 19014
rect 29112 19012 29168 19014
rect 29192 19012 29248 19014
rect 29272 19012 29328 19014
rect 28814 18672 28870 18728
rect 21012 16346 21068 16348
rect 21092 16346 21148 16348
rect 21172 16346 21228 16348
rect 21252 16346 21308 16348
rect 21012 16294 21058 16346
rect 21058 16294 21068 16346
rect 21092 16294 21122 16346
rect 21122 16294 21134 16346
rect 21134 16294 21148 16346
rect 21172 16294 21186 16346
rect 21186 16294 21198 16346
rect 21198 16294 21228 16346
rect 21252 16294 21262 16346
rect 21262 16294 21308 16346
rect 21012 16292 21068 16294
rect 21092 16292 21148 16294
rect 21172 16292 21228 16294
rect 21252 16292 21308 16294
rect 21672 15802 21728 15804
rect 21752 15802 21808 15804
rect 21832 15802 21888 15804
rect 21912 15802 21968 15804
rect 21672 15750 21718 15802
rect 21718 15750 21728 15802
rect 21752 15750 21782 15802
rect 21782 15750 21794 15802
rect 21794 15750 21808 15802
rect 21832 15750 21846 15802
rect 21846 15750 21858 15802
rect 21858 15750 21888 15802
rect 21912 15750 21922 15802
rect 21922 15750 21968 15802
rect 21672 15748 21728 15750
rect 21752 15748 21808 15750
rect 21832 15748 21888 15750
rect 21912 15748 21968 15750
rect 21012 15258 21068 15260
rect 21092 15258 21148 15260
rect 21172 15258 21228 15260
rect 21252 15258 21308 15260
rect 21012 15206 21058 15258
rect 21058 15206 21068 15258
rect 21092 15206 21122 15258
rect 21122 15206 21134 15258
rect 21134 15206 21148 15258
rect 21172 15206 21186 15258
rect 21186 15206 21198 15258
rect 21198 15206 21228 15258
rect 21252 15206 21262 15258
rect 21262 15206 21308 15258
rect 21012 15204 21068 15206
rect 21092 15204 21148 15206
rect 21172 15204 21228 15206
rect 21252 15204 21308 15206
rect 21012 14170 21068 14172
rect 21092 14170 21148 14172
rect 21172 14170 21228 14172
rect 21252 14170 21308 14172
rect 21012 14118 21058 14170
rect 21058 14118 21068 14170
rect 21092 14118 21122 14170
rect 21122 14118 21134 14170
rect 21134 14118 21148 14170
rect 21172 14118 21186 14170
rect 21186 14118 21198 14170
rect 21198 14118 21228 14170
rect 21252 14118 21262 14170
rect 21262 14118 21308 14170
rect 21012 14116 21068 14118
rect 21092 14116 21148 14118
rect 21172 14116 21228 14118
rect 21252 14116 21308 14118
rect 21672 14714 21728 14716
rect 21752 14714 21808 14716
rect 21832 14714 21888 14716
rect 21912 14714 21968 14716
rect 21672 14662 21718 14714
rect 21718 14662 21728 14714
rect 21752 14662 21782 14714
rect 21782 14662 21794 14714
rect 21794 14662 21808 14714
rect 21832 14662 21846 14714
rect 21846 14662 21858 14714
rect 21858 14662 21888 14714
rect 21912 14662 21922 14714
rect 21922 14662 21968 14714
rect 21672 14660 21728 14662
rect 21752 14660 21808 14662
rect 21832 14660 21888 14662
rect 21912 14660 21968 14662
rect 21012 13082 21068 13084
rect 21092 13082 21148 13084
rect 21172 13082 21228 13084
rect 21252 13082 21308 13084
rect 21012 13030 21058 13082
rect 21058 13030 21068 13082
rect 21092 13030 21122 13082
rect 21122 13030 21134 13082
rect 21134 13030 21148 13082
rect 21172 13030 21186 13082
rect 21186 13030 21198 13082
rect 21198 13030 21228 13082
rect 21252 13030 21262 13082
rect 21262 13030 21308 13082
rect 21012 13028 21068 13030
rect 21092 13028 21148 13030
rect 21172 13028 21228 13030
rect 21252 13028 21308 13030
rect 21672 13626 21728 13628
rect 21752 13626 21808 13628
rect 21832 13626 21888 13628
rect 21912 13626 21968 13628
rect 21672 13574 21718 13626
rect 21718 13574 21728 13626
rect 21752 13574 21782 13626
rect 21782 13574 21794 13626
rect 21794 13574 21808 13626
rect 21832 13574 21846 13626
rect 21846 13574 21858 13626
rect 21858 13574 21888 13626
rect 21912 13574 21922 13626
rect 21922 13574 21968 13626
rect 21672 13572 21728 13574
rect 21752 13572 21808 13574
rect 21832 13572 21888 13574
rect 21912 13572 21968 13574
rect 20258 9580 20314 9616
rect 20258 9560 20260 9580
rect 20260 9560 20312 9580
rect 20312 9560 20314 9580
rect 18602 6840 18658 6896
rect 18050 5208 18106 5264
rect 18602 5072 18658 5128
rect 19246 5228 19302 5264
rect 19246 5208 19248 5228
rect 19248 5208 19300 5228
rect 19300 5208 19302 5228
rect 21012 11994 21068 11996
rect 21092 11994 21148 11996
rect 21172 11994 21228 11996
rect 21252 11994 21308 11996
rect 21012 11942 21058 11994
rect 21058 11942 21068 11994
rect 21092 11942 21122 11994
rect 21122 11942 21134 11994
rect 21134 11942 21148 11994
rect 21172 11942 21186 11994
rect 21186 11942 21198 11994
rect 21198 11942 21228 11994
rect 21252 11942 21262 11994
rect 21262 11942 21308 11994
rect 21012 11940 21068 11942
rect 21092 11940 21148 11942
rect 21172 11940 21228 11942
rect 21252 11940 21308 11942
rect 21012 10906 21068 10908
rect 21092 10906 21148 10908
rect 21172 10906 21228 10908
rect 21252 10906 21308 10908
rect 21012 10854 21058 10906
rect 21058 10854 21068 10906
rect 21092 10854 21122 10906
rect 21122 10854 21134 10906
rect 21134 10854 21148 10906
rect 21172 10854 21186 10906
rect 21186 10854 21198 10906
rect 21198 10854 21228 10906
rect 21252 10854 21262 10906
rect 21262 10854 21308 10906
rect 21012 10852 21068 10854
rect 21092 10852 21148 10854
rect 21172 10852 21228 10854
rect 21252 10852 21308 10854
rect 21012 9818 21068 9820
rect 21092 9818 21148 9820
rect 21172 9818 21228 9820
rect 21252 9818 21308 9820
rect 21012 9766 21058 9818
rect 21058 9766 21068 9818
rect 21092 9766 21122 9818
rect 21122 9766 21134 9818
rect 21134 9766 21148 9818
rect 21172 9766 21186 9818
rect 21186 9766 21198 9818
rect 21198 9766 21228 9818
rect 21252 9766 21262 9818
rect 21262 9766 21308 9818
rect 21012 9764 21068 9766
rect 21092 9764 21148 9766
rect 21172 9764 21228 9766
rect 21252 9764 21308 9766
rect 20718 5108 20720 5128
rect 20720 5108 20772 5128
rect 20772 5108 20774 5128
rect 20718 5072 20774 5108
rect 21012 8730 21068 8732
rect 21092 8730 21148 8732
rect 21172 8730 21228 8732
rect 21252 8730 21308 8732
rect 21012 8678 21058 8730
rect 21058 8678 21068 8730
rect 21092 8678 21122 8730
rect 21122 8678 21134 8730
rect 21134 8678 21148 8730
rect 21172 8678 21186 8730
rect 21186 8678 21198 8730
rect 21198 8678 21228 8730
rect 21252 8678 21262 8730
rect 21262 8678 21308 8730
rect 21012 8676 21068 8678
rect 21092 8676 21148 8678
rect 21172 8676 21228 8678
rect 21252 8676 21308 8678
rect 21012 7642 21068 7644
rect 21092 7642 21148 7644
rect 21172 7642 21228 7644
rect 21252 7642 21308 7644
rect 21012 7590 21058 7642
rect 21058 7590 21068 7642
rect 21092 7590 21122 7642
rect 21122 7590 21134 7642
rect 21134 7590 21148 7642
rect 21172 7590 21186 7642
rect 21186 7590 21198 7642
rect 21198 7590 21228 7642
rect 21252 7590 21262 7642
rect 21262 7590 21308 7642
rect 21012 7588 21068 7590
rect 21092 7588 21148 7590
rect 21172 7588 21228 7590
rect 21252 7588 21308 7590
rect 21672 12538 21728 12540
rect 21752 12538 21808 12540
rect 21832 12538 21888 12540
rect 21912 12538 21968 12540
rect 21672 12486 21718 12538
rect 21718 12486 21728 12538
rect 21752 12486 21782 12538
rect 21782 12486 21794 12538
rect 21794 12486 21808 12538
rect 21832 12486 21846 12538
rect 21846 12486 21858 12538
rect 21858 12486 21888 12538
rect 21912 12486 21922 12538
rect 21922 12486 21968 12538
rect 21672 12484 21728 12486
rect 21752 12484 21808 12486
rect 21832 12484 21888 12486
rect 21912 12484 21968 12486
rect 21672 11450 21728 11452
rect 21752 11450 21808 11452
rect 21832 11450 21888 11452
rect 21912 11450 21968 11452
rect 21672 11398 21718 11450
rect 21718 11398 21728 11450
rect 21752 11398 21782 11450
rect 21782 11398 21794 11450
rect 21794 11398 21808 11450
rect 21832 11398 21846 11450
rect 21846 11398 21858 11450
rect 21858 11398 21888 11450
rect 21912 11398 21922 11450
rect 21922 11398 21968 11450
rect 21672 11396 21728 11398
rect 21752 11396 21808 11398
rect 21832 11396 21888 11398
rect 21912 11396 21968 11398
rect 28372 18522 28428 18524
rect 28452 18522 28508 18524
rect 28532 18522 28588 18524
rect 28612 18522 28668 18524
rect 28372 18470 28418 18522
rect 28418 18470 28428 18522
rect 28452 18470 28482 18522
rect 28482 18470 28494 18522
rect 28494 18470 28508 18522
rect 28532 18470 28546 18522
rect 28546 18470 28558 18522
rect 28558 18470 28588 18522
rect 28612 18470 28622 18522
rect 28622 18470 28668 18522
rect 28372 18468 28428 18470
rect 28452 18468 28508 18470
rect 28532 18468 28588 18470
rect 28612 18468 28668 18470
rect 29032 17978 29088 17980
rect 29112 17978 29168 17980
rect 29192 17978 29248 17980
rect 29272 17978 29328 17980
rect 29032 17926 29078 17978
rect 29078 17926 29088 17978
rect 29112 17926 29142 17978
rect 29142 17926 29154 17978
rect 29154 17926 29168 17978
rect 29192 17926 29206 17978
rect 29206 17926 29218 17978
rect 29218 17926 29248 17978
rect 29272 17926 29282 17978
rect 29282 17926 29328 17978
rect 29032 17924 29088 17926
rect 29112 17924 29168 17926
rect 29192 17924 29248 17926
rect 29272 17924 29328 17926
rect 28372 17434 28428 17436
rect 28452 17434 28508 17436
rect 28532 17434 28588 17436
rect 28612 17434 28668 17436
rect 28372 17382 28418 17434
rect 28418 17382 28428 17434
rect 28452 17382 28482 17434
rect 28482 17382 28494 17434
rect 28494 17382 28508 17434
rect 28532 17382 28546 17434
rect 28546 17382 28558 17434
rect 28558 17382 28588 17434
rect 28612 17382 28622 17434
rect 28622 17382 28668 17434
rect 28372 17380 28428 17382
rect 28452 17380 28508 17382
rect 28532 17380 28588 17382
rect 28612 17380 28668 17382
rect 29032 16890 29088 16892
rect 29112 16890 29168 16892
rect 29192 16890 29248 16892
rect 29272 16890 29328 16892
rect 29032 16838 29078 16890
rect 29078 16838 29088 16890
rect 29112 16838 29142 16890
rect 29142 16838 29154 16890
rect 29154 16838 29168 16890
rect 29192 16838 29206 16890
rect 29206 16838 29218 16890
rect 29218 16838 29248 16890
rect 29272 16838 29282 16890
rect 29282 16838 29328 16890
rect 29032 16836 29088 16838
rect 29112 16836 29168 16838
rect 29192 16836 29248 16838
rect 29272 16836 29328 16838
rect 28372 16346 28428 16348
rect 28452 16346 28508 16348
rect 28532 16346 28588 16348
rect 28612 16346 28668 16348
rect 28372 16294 28418 16346
rect 28418 16294 28428 16346
rect 28452 16294 28482 16346
rect 28482 16294 28494 16346
rect 28494 16294 28508 16346
rect 28532 16294 28546 16346
rect 28546 16294 28558 16346
rect 28558 16294 28588 16346
rect 28612 16294 28622 16346
rect 28622 16294 28668 16346
rect 28372 16292 28428 16294
rect 28452 16292 28508 16294
rect 28532 16292 28588 16294
rect 28612 16292 28668 16294
rect 30654 19916 30710 19952
rect 30654 19896 30656 19916
rect 30656 19896 30708 19916
rect 30708 19896 30710 19916
rect 30654 19760 30710 19816
rect 29032 15802 29088 15804
rect 29112 15802 29168 15804
rect 29192 15802 29248 15804
rect 29272 15802 29328 15804
rect 29032 15750 29078 15802
rect 29078 15750 29088 15802
rect 29112 15750 29142 15802
rect 29142 15750 29154 15802
rect 29154 15750 29168 15802
rect 29192 15750 29206 15802
rect 29206 15750 29218 15802
rect 29218 15750 29248 15802
rect 29272 15750 29282 15802
rect 29282 15750 29328 15802
rect 29032 15748 29088 15750
rect 29112 15748 29168 15750
rect 29192 15748 29248 15750
rect 29272 15748 29328 15750
rect 26146 12824 26202 12880
rect 21672 10362 21728 10364
rect 21752 10362 21808 10364
rect 21832 10362 21888 10364
rect 21912 10362 21968 10364
rect 21672 10310 21718 10362
rect 21718 10310 21728 10362
rect 21752 10310 21782 10362
rect 21782 10310 21794 10362
rect 21794 10310 21808 10362
rect 21832 10310 21846 10362
rect 21846 10310 21858 10362
rect 21858 10310 21888 10362
rect 21912 10310 21922 10362
rect 21922 10310 21968 10362
rect 21672 10308 21728 10310
rect 21752 10308 21808 10310
rect 21832 10308 21888 10310
rect 21912 10308 21968 10310
rect 21822 9424 21878 9480
rect 21672 9274 21728 9276
rect 21752 9274 21808 9276
rect 21832 9274 21888 9276
rect 21912 9274 21968 9276
rect 21672 9222 21718 9274
rect 21718 9222 21728 9274
rect 21752 9222 21782 9274
rect 21782 9222 21794 9274
rect 21794 9222 21808 9274
rect 21832 9222 21846 9274
rect 21846 9222 21858 9274
rect 21858 9222 21888 9274
rect 21912 9222 21922 9274
rect 21922 9222 21968 9274
rect 21672 9220 21728 9222
rect 21752 9220 21808 9222
rect 21832 9220 21888 9222
rect 21912 9220 21968 9222
rect 21730 8372 21732 8392
rect 21732 8372 21784 8392
rect 21784 8372 21786 8392
rect 22466 9424 22522 9480
rect 21730 8336 21786 8372
rect 21672 8186 21728 8188
rect 21752 8186 21808 8188
rect 21832 8186 21888 8188
rect 21912 8186 21968 8188
rect 21672 8134 21718 8186
rect 21718 8134 21728 8186
rect 21752 8134 21782 8186
rect 21782 8134 21794 8186
rect 21794 8134 21808 8186
rect 21832 8134 21846 8186
rect 21846 8134 21858 8186
rect 21858 8134 21888 8186
rect 21912 8134 21922 8186
rect 21922 8134 21968 8186
rect 21672 8132 21728 8134
rect 21752 8132 21808 8134
rect 21832 8132 21888 8134
rect 21912 8132 21968 8134
rect 21672 7098 21728 7100
rect 21752 7098 21808 7100
rect 21832 7098 21888 7100
rect 21912 7098 21968 7100
rect 21672 7046 21718 7098
rect 21718 7046 21728 7098
rect 21752 7046 21782 7098
rect 21782 7046 21794 7098
rect 21794 7046 21808 7098
rect 21832 7046 21846 7098
rect 21846 7046 21858 7098
rect 21858 7046 21888 7098
rect 21912 7046 21922 7098
rect 21922 7046 21968 7098
rect 21672 7044 21728 7046
rect 21752 7044 21808 7046
rect 21832 7044 21888 7046
rect 21912 7044 21968 7046
rect 23570 9596 23572 9616
rect 23572 9596 23624 9616
rect 23624 9596 23626 9616
rect 23570 9560 23626 9596
rect 23662 9460 23664 9480
rect 23664 9460 23716 9480
rect 23716 9460 23718 9480
rect 23662 9424 23718 9460
rect 24582 12144 24638 12200
rect 24490 11872 24546 11928
rect 23386 8336 23442 8392
rect 26606 12144 26662 12200
rect 26238 9444 26294 9480
rect 28372 15258 28428 15260
rect 28452 15258 28508 15260
rect 28532 15258 28588 15260
rect 28612 15258 28668 15260
rect 28372 15206 28418 15258
rect 28418 15206 28428 15258
rect 28452 15206 28482 15258
rect 28482 15206 28494 15258
rect 28494 15206 28508 15258
rect 28532 15206 28546 15258
rect 28546 15206 28558 15258
rect 28558 15206 28588 15258
rect 28612 15206 28622 15258
rect 28622 15206 28668 15258
rect 28372 15204 28428 15206
rect 28452 15204 28508 15206
rect 28532 15204 28588 15206
rect 28612 15204 28668 15206
rect 29032 14714 29088 14716
rect 29112 14714 29168 14716
rect 29192 14714 29248 14716
rect 29272 14714 29328 14716
rect 29032 14662 29078 14714
rect 29078 14662 29088 14714
rect 29112 14662 29142 14714
rect 29142 14662 29154 14714
rect 29154 14662 29168 14714
rect 29192 14662 29206 14714
rect 29206 14662 29218 14714
rect 29218 14662 29248 14714
rect 29272 14662 29282 14714
rect 29282 14662 29328 14714
rect 29032 14660 29088 14662
rect 29112 14660 29168 14662
rect 29192 14660 29248 14662
rect 29272 14660 29328 14662
rect 28372 14170 28428 14172
rect 28452 14170 28508 14172
rect 28532 14170 28588 14172
rect 28612 14170 28668 14172
rect 28372 14118 28418 14170
rect 28418 14118 28428 14170
rect 28452 14118 28482 14170
rect 28482 14118 28494 14170
rect 28494 14118 28508 14170
rect 28532 14118 28546 14170
rect 28546 14118 28558 14170
rect 28558 14118 28588 14170
rect 28612 14118 28622 14170
rect 28622 14118 28668 14170
rect 28372 14116 28428 14118
rect 28452 14116 28508 14118
rect 28532 14116 28588 14118
rect 28612 14116 28668 14118
rect 28998 13812 29000 13832
rect 29000 13812 29052 13832
rect 29052 13812 29054 13832
rect 28998 13776 29054 13812
rect 29032 13626 29088 13628
rect 29112 13626 29168 13628
rect 29192 13626 29248 13628
rect 29272 13626 29328 13628
rect 29032 13574 29078 13626
rect 29078 13574 29088 13626
rect 29112 13574 29142 13626
rect 29142 13574 29154 13626
rect 29154 13574 29168 13626
rect 29192 13574 29206 13626
rect 29206 13574 29218 13626
rect 29218 13574 29248 13626
rect 29272 13574 29282 13626
rect 29282 13574 29328 13626
rect 29032 13572 29088 13574
rect 29112 13572 29168 13574
rect 29192 13572 29248 13574
rect 29272 13572 29328 13574
rect 28998 13252 29054 13288
rect 28998 13232 29000 13252
rect 29000 13232 29052 13252
rect 29052 13232 29054 13252
rect 26238 9424 26240 9444
rect 26240 9424 26292 9444
rect 26292 9424 26294 9444
rect 25134 8472 25190 8528
rect 21012 6554 21068 6556
rect 21092 6554 21148 6556
rect 21172 6554 21228 6556
rect 21252 6554 21308 6556
rect 21012 6502 21058 6554
rect 21058 6502 21068 6554
rect 21092 6502 21122 6554
rect 21122 6502 21134 6554
rect 21134 6502 21148 6554
rect 21172 6502 21186 6554
rect 21186 6502 21198 6554
rect 21198 6502 21228 6554
rect 21252 6502 21262 6554
rect 21262 6502 21308 6554
rect 21012 6500 21068 6502
rect 21092 6500 21148 6502
rect 21172 6500 21228 6502
rect 21252 6500 21308 6502
rect 21362 6296 21418 6352
rect 21672 6010 21728 6012
rect 21752 6010 21808 6012
rect 21832 6010 21888 6012
rect 21912 6010 21968 6012
rect 21672 5958 21718 6010
rect 21718 5958 21728 6010
rect 21752 5958 21782 6010
rect 21782 5958 21794 6010
rect 21794 5958 21808 6010
rect 21832 5958 21846 6010
rect 21846 5958 21858 6010
rect 21858 5958 21888 6010
rect 21912 5958 21922 6010
rect 21922 5958 21968 6010
rect 21672 5956 21728 5958
rect 21752 5956 21808 5958
rect 21832 5956 21888 5958
rect 21912 5956 21968 5958
rect 21012 5466 21068 5468
rect 21092 5466 21148 5468
rect 21172 5466 21228 5468
rect 21252 5466 21308 5468
rect 21012 5414 21058 5466
rect 21058 5414 21068 5466
rect 21092 5414 21122 5466
rect 21122 5414 21134 5466
rect 21134 5414 21148 5466
rect 21172 5414 21186 5466
rect 21186 5414 21198 5466
rect 21198 5414 21228 5466
rect 21252 5414 21262 5466
rect 21262 5414 21308 5466
rect 21012 5412 21068 5414
rect 21092 5412 21148 5414
rect 21172 5412 21228 5414
rect 21252 5412 21308 5414
rect 22742 5616 22798 5672
rect 21672 4922 21728 4924
rect 21752 4922 21808 4924
rect 21832 4922 21888 4924
rect 21912 4922 21968 4924
rect 21672 4870 21718 4922
rect 21718 4870 21728 4922
rect 21752 4870 21782 4922
rect 21782 4870 21794 4922
rect 21794 4870 21808 4922
rect 21832 4870 21846 4922
rect 21846 4870 21858 4922
rect 21858 4870 21888 4922
rect 21912 4870 21922 4922
rect 21922 4870 21968 4922
rect 21672 4868 21728 4870
rect 21752 4868 21808 4870
rect 21832 4868 21888 4870
rect 21912 4868 21968 4870
rect 21012 4378 21068 4380
rect 21092 4378 21148 4380
rect 21172 4378 21228 4380
rect 21252 4378 21308 4380
rect 21012 4326 21058 4378
rect 21058 4326 21068 4378
rect 21092 4326 21122 4378
rect 21122 4326 21134 4378
rect 21134 4326 21148 4378
rect 21172 4326 21186 4378
rect 21186 4326 21198 4378
rect 21198 4326 21228 4378
rect 21252 4326 21262 4378
rect 21262 4326 21308 4378
rect 21012 4324 21068 4326
rect 21092 4324 21148 4326
rect 21172 4324 21228 4326
rect 21252 4324 21308 4326
rect 21672 3834 21728 3836
rect 21752 3834 21808 3836
rect 21832 3834 21888 3836
rect 21912 3834 21968 3836
rect 21672 3782 21718 3834
rect 21718 3782 21728 3834
rect 21752 3782 21782 3834
rect 21782 3782 21794 3834
rect 21794 3782 21808 3834
rect 21832 3782 21846 3834
rect 21846 3782 21858 3834
rect 21858 3782 21888 3834
rect 21912 3782 21922 3834
rect 21922 3782 21968 3834
rect 21672 3780 21728 3782
rect 21752 3780 21808 3782
rect 21832 3780 21888 3782
rect 21912 3780 21968 3782
rect 27526 9424 27582 9480
rect 28372 13082 28428 13084
rect 28452 13082 28508 13084
rect 28532 13082 28588 13084
rect 28612 13082 28668 13084
rect 28372 13030 28418 13082
rect 28418 13030 28428 13082
rect 28452 13030 28482 13082
rect 28482 13030 28494 13082
rect 28494 13030 28508 13082
rect 28532 13030 28546 13082
rect 28546 13030 28558 13082
rect 28558 13030 28588 13082
rect 28612 13030 28622 13082
rect 28622 13030 28668 13082
rect 28372 13028 28428 13030
rect 28452 13028 28508 13030
rect 28532 13028 28588 13030
rect 28612 13028 28668 13030
rect 28906 12824 28962 12880
rect 29550 13776 29606 13832
rect 29032 12538 29088 12540
rect 29112 12538 29168 12540
rect 29192 12538 29248 12540
rect 29272 12538 29328 12540
rect 29032 12486 29078 12538
rect 29078 12486 29088 12538
rect 29112 12486 29142 12538
rect 29142 12486 29154 12538
rect 29154 12486 29168 12538
rect 29192 12486 29206 12538
rect 29206 12486 29218 12538
rect 29218 12486 29248 12538
rect 29272 12486 29282 12538
rect 29282 12486 29328 12538
rect 29032 12484 29088 12486
rect 29112 12484 29168 12486
rect 29192 12484 29248 12486
rect 29272 12484 29328 12486
rect 28372 11994 28428 11996
rect 28452 11994 28508 11996
rect 28532 11994 28588 11996
rect 28612 11994 28668 11996
rect 28372 11942 28418 11994
rect 28418 11942 28428 11994
rect 28452 11942 28482 11994
rect 28482 11942 28494 11994
rect 28494 11942 28508 11994
rect 28532 11942 28546 11994
rect 28546 11942 28558 11994
rect 28558 11942 28588 11994
rect 28612 11942 28622 11994
rect 28622 11942 28668 11994
rect 28372 11940 28428 11942
rect 28452 11940 28508 11942
rect 28532 11940 28588 11942
rect 28612 11940 28668 11942
rect 31666 32000 31722 32056
rect 31114 27376 31170 27432
rect 33138 33360 33194 33416
rect 33046 30640 33102 30696
rect 33138 27240 33194 27296
rect 33138 25236 33140 25256
rect 33140 25236 33192 25256
rect 33192 25236 33194 25256
rect 33138 25200 33194 25236
rect 29734 13232 29790 13288
rect 29032 11450 29088 11452
rect 29112 11450 29168 11452
rect 29192 11450 29248 11452
rect 29272 11450 29328 11452
rect 29032 11398 29078 11450
rect 29078 11398 29088 11450
rect 29112 11398 29142 11450
rect 29142 11398 29154 11450
rect 29154 11398 29168 11450
rect 29192 11398 29206 11450
rect 29206 11398 29218 11450
rect 29218 11398 29248 11450
rect 29272 11398 29282 11450
rect 29282 11398 29328 11450
rect 29032 11396 29088 11398
rect 29112 11396 29168 11398
rect 29192 11396 29248 11398
rect 29272 11396 29328 11398
rect 28372 10906 28428 10908
rect 28452 10906 28508 10908
rect 28532 10906 28588 10908
rect 28612 10906 28668 10908
rect 28372 10854 28418 10906
rect 28418 10854 28428 10906
rect 28452 10854 28482 10906
rect 28482 10854 28494 10906
rect 28494 10854 28508 10906
rect 28532 10854 28546 10906
rect 28546 10854 28558 10906
rect 28558 10854 28588 10906
rect 28612 10854 28622 10906
rect 28622 10854 28668 10906
rect 28372 10852 28428 10854
rect 28452 10852 28508 10854
rect 28532 10852 28588 10854
rect 28612 10852 28668 10854
rect 28372 9818 28428 9820
rect 28452 9818 28508 9820
rect 28532 9818 28588 9820
rect 28612 9818 28668 9820
rect 28372 9766 28418 9818
rect 28418 9766 28428 9818
rect 28452 9766 28482 9818
rect 28482 9766 28494 9818
rect 28494 9766 28508 9818
rect 28532 9766 28546 9818
rect 28546 9766 28558 9818
rect 28558 9766 28588 9818
rect 28612 9766 28622 9818
rect 28622 9766 28668 9818
rect 28372 9764 28428 9766
rect 28452 9764 28508 9766
rect 28532 9764 28588 9766
rect 28612 9764 28668 9766
rect 25870 7928 25926 7984
rect 21012 3290 21068 3292
rect 21092 3290 21148 3292
rect 21172 3290 21228 3292
rect 21252 3290 21308 3292
rect 21012 3238 21058 3290
rect 21058 3238 21068 3290
rect 21092 3238 21122 3290
rect 21122 3238 21134 3290
rect 21134 3238 21148 3290
rect 21172 3238 21186 3290
rect 21186 3238 21198 3290
rect 21198 3238 21228 3290
rect 21252 3238 21262 3290
rect 21262 3238 21308 3290
rect 21012 3236 21068 3238
rect 21092 3236 21148 3238
rect 21172 3236 21228 3238
rect 21252 3236 21308 3238
rect 21672 2746 21728 2748
rect 21752 2746 21808 2748
rect 21832 2746 21888 2748
rect 21912 2746 21968 2748
rect 21672 2694 21718 2746
rect 21718 2694 21728 2746
rect 21752 2694 21782 2746
rect 21782 2694 21794 2746
rect 21794 2694 21808 2746
rect 21832 2694 21846 2746
rect 21846 2694 21858 2746
rect 21858 2694 21888 2746
rect 21912 2694 21922 2746
rect 21922 2694 21968 2746
rect 21672 2692 21728 2694
rect 21752 2692 21808 2694
rect 21832 2692 21888 2694
rect 21912 2692 21968 2694
rect 28630 9424 28686 9480
rect 28372 8730 28428 8732
rect 28452 8730 28508 8732
rect 28532 8730 28588 8732
rect 28612 8730 28668 8732
rect 28372 8678 28418 8730
rect 28418 8678 28428 8730
rect 28452 8678 28482 8730
rect 28482 8678 28494 8730
rect 28494 8678 28508 8730
rect 28532 8678 28546 8730
rect 28546 8678 28558 8730
rect 28558 8678 28588 8730
rect 28612 8678 28622 8730
rect 28622 8678 28668 8730
rect 28372 8676 28428 8678
rect 28452 8676 28508 8678
rect 28532 8676 28588 8678
rect 28612 8676 28668 8678
rect 28446 8472 28502 8528
rect 29032 10362 29088 10364
rect 29112 10362 29168 10364
rect 29192 10362 29248 10364
rect 29272 10362 29328 10364
rect 29032 10310 29078 10362
rect 29078 10310 29088 10362
rect 29112 10310 29142 10362
rect 29142 10310 29154 10362
rect 29154 10310 29168 10362
rect 29192 10310 29206 10362
rect 29206 10310 29218 10362
rect 29218 10310 29248 10362
rect 29272 10310 29282 10362
rect 29282 10310 29328 10362
rect 29032 10308 29088 10310
rect 29112 10308 29168 10310
rect 29192 10308 29248 10310
rect 29272 10308 29328 10310
rect 29182 9444 29238 9480
rect 29182 9424 29184 9444
rect 29184 9424 29236 9444
rect 29236 9424 29238 9444
rect 29032 9274 29088 9276
rect 29112 9274 29168 9276
rect 29192 9274 29248 9276
rect 29272 9274 29328 9276
rect 29032 9222 29078 9274
rect 29078 9222 29088 9274
rect 29112 9222 29142 9274
rect 29142 9222 29154 9274
rect 29154 9222 29168 9274
rect 29192 9222 29206 9274
rect 29206 9222 29218 9274
rect 29218 9222 29248 9274
rect 29272 9222 29282 9274
rect 29282 9222 29328 9274
rect 29032 9220 29088 9222
rect 29112 9220 29168 9222
rect 29192 9220 29248 9222
rect 29272 9220 29328 9222
rect 28170 7948 28226 7984
rect 28170 7928 28172 7948
rect 28172 7928 28224 7948
rect 28224 7928 28226 7948
rect 28372 7642 28428 7644
rect 28452 7642 28508 7644
rect 28532 7642 28588 7644
rect 28612 7642 28668 7644
rect 28372 7590 28418 7642
rect 28418 7590 28428 7642
rect 28452 7590 28482 7642
rect 28482 7590 28494 7642
rect 28494 7590 28508 7642
rect 28532 7590 28546 7642
rect 28546 7590 28558 7642
rect 28558 7590 28588 7642
rect 28612 7590 28622 7642
rect 28622 7590 28668 7642
rect 28372 7588 28428 7590
rect 28452 7588 28508 7590
rect 28532 7588 28588 7590
rect 28612 7588 28668 7590
rect 29032 8186 29088 8188
rect 29112 8186 29168 8188
rect 29192 8186 29248 8188
rect 29272 8186 29328 8188
rect 29032 8134 29078 8186
rect 29078 8134 29088 8186
rect 29112 8134 29142 8186
rect 29142 8134 29154 8186
rect 29154 8134 29168 8186
rect 29192 8134 29206 8186
rect 29206 8134 29218 8186
rect 29218 8134 29248 8186
rect 29272 8134 29282 8186
rect 29282 8134 29328 8186
rect 29032 8132 29088 8134
rect 29112 8132 29168 8134
rect 29192 8132 29248 8134
rect 29272 8132 29328 8134
rect 29458 7792 29514 7848
rect 28372 6554 28428 6556
rect 28452 6554 28508 6556
rect 28532 6554 28588 6556
rect 28612 6554 28668 6556
rect 28372 6502 28418 6554
rect 28418 6502 28428 6554
rect 28452 6502 28482 6554
rect 28482 6502 28494 6554
rect 28494 6502 28508 6554
rect 28532 6502 28546 6554
rect 28546 6502 28558 6554
rect 28558 6502 28588 6554
rect 28612 6502 28622 6554
rect 28622 6502 28668 6554
rect 28372 6500 28428 6502
rect 28452 6500 28508 6502
rect 28532 6500 28588 6502
rect 28612 6500 28668 6502
rect 29032 7098 29088 7100
rect 29112 7098 29168 7100
rect 29192 7098 29248 7100
rect 29272 7098 29328 7100
rect 29032 7046 29078 7098
rect 29078 7046 29088 7098
rect 29112 7046 29142 7098
rect 29142 7046 29154 7098
rect 29154 7046 29168 7098
rect 29192 7046 29206 7098
rect 29206 7046 29218 7098
rect 29218 7046 29248 7098
rect 29272 7046 29282 7098
rect 29282 7046 29328 7098
rect 29032 7044 29088 7046
rect 29112 7044 29168 7046
rect 29192 7044 29248 7046
rect 29272 7044 29328 7046
rect 29032 6010 29088 6012
rect 29112 6010 29168 6012
rect 29192 6010 29248 6012
rect 29272 6010 29328 6012
rect 29032 5958 29078 6010
rect 29078 5958 29088 6010
rect 29112 5958 29142 6010
rect 29142 5958 29154 6010
rect 29154 5958 29168 6010
rect 29192 5958 29206 6010
rect 29206 5958 29218 6010
rect 29218 5958 29248 6010
rect 29272 5958 29282 6010
rect 29282 5958 29328 6010
rect 29032 5956 29088 5958
rect 29112 5956 29168 5958
rect 29192 5956 29248 5958
rect 29272 5956 29328 5958
rect 29734 5616 29790 5672
rect 28372 5466 28428 5468
rect 28452 5466 28508 5468
rect 28532 5466 28588 5468
rect 28612 5466 28668 5468
rect 28372 5414 28418 5466
rect 28418 5414 28428 5466
rect 28452 5414 28482 5466
rect 28482 5414 28494 5466
rect 28494 5414 28508 5466
rect 28532 5414 28546 5466
rect 28546 5414 28558 5466
rect 28558 5414 28588 5466
rect 28612 5414 28622 5466
rect 28622 5414 28668 5466
rect 28372 5412 28428 5414
rect 28452 5412 28508 5414
rect 28532 5412 28588 5414
rect 28612 5412 28668 5414
rect 29032 4922 29088 4924
rect 29112 4922 29168 4924
rect 29192 4922 29248 4924
rect 29272 4922 29328 4924
rect 29032 4870 29078 4922
rect 29078 4870 29088 4922
rect 29112 4870 29142 4922
rect 29142 4870 29154 4922
rect 29154 4870 29168 4922
rect 29192 4870 29206 4922
rect 29206 4870 29218 4922
rect 29218 4870 29248 4922
rect 29272 4870 29282 4922
rect 29282 4870 29328 4922
rect 29032 4868 29088 4870
rect 29112 4868 29168 4870
rect 29192 4868 29248 4870
rect 29272 4868 29328 4870
rect 30562 13404 30564 13424
rect 30564 13404 30616 13424
rect 30616 13404 30618 13424
rect 30562 13368 30618 13404
rect 33138 23840 33194 23896
rect 31666 22480 31722 22536
rect 33046 20440 33102 20496
rect 33138 19080 33194 19136
rect 31022 13776 31078 13832
rect 28372 4378 28428 4380
rect 28452 4378 28508 4380
rect 28532 4378 28588 4380
rect 28612 4378 28668 4380
rect 28372 4326 28418 4378
rect 28418 4326 28428 4378
rect 28452 4326 28482 4378
rect 28482 4326 28494 4378
rect 28494 4326 28508 4378
rect 28532 4326 28546 4378
rect 28546 4326 28558 4378
rect 28558 4326 28588 4378
rect 28612 4326 28622 4378
rect 28622 4326 28668 4378
rect 28372 4324 28428 4326
rect 28452 4324 28508 4326
rect 28532 4324 28588 4326
rect 28612 4324 28668 4326
rect 33138 17040 33194 17096
rect 33138 15680 33194 15736
rect 33138 14356 33140 14376
rect 33140 14356 33192 14376
rect 33192 14356 33194 14376
rect 33138 14320 33194 14356
rect 31758 13368 31814 13424
rect 33138 12300 33194 12336
rect 33138 12280 33140 12300
rect 33140 12280 33192 12300
rect 33192 12280 33194 12300
rect 31390 10920 31446 10976
rect 29032 3834 29088 3836
rect 29112 3834 29168 3836
rect 29192 3834 29248 3836
rect 29272 3834 29328 3836
rect 29032 3782 29078 3834
rect 29078 3782 29088 3834
rect 29112 3782 29142 3834
rect 29142 3782 29154 3834
rect 29154 3782 29168 3834
rect 29192 3782 29206 3834
rect 29206 3782 29218 3834
rect 29218 3782 29248 3834
rect 29272 3782 29282 3834
rect 29282 3782 29328 3834
rect 29032 3780 29088 3782
rect 29112 3780 29168 3782
rect 29192 3780 29248 3782
rect 29272 3780 29328 3782
rect 28372 3290 28428 3292
rect 28452 3290 28508 3292
rect 28532 3290 28588 3292
rect 28612 3290 28668 3292
rect 28372 3238 28418 3290
rect 28418 3238 28428 3290
rect 28452 3238 28482 3290
rect 28482 3238 28494 3290
rect 28494 3238 28508 3290
rect 28532 3238 28546 3290
rect 28546 3238 28558 3290
rect 28558 3238 28588 3290
rect 28612 3238 28622 3290
rect 28622 3238 28668 3290
rect 28372 3236 28428 3238
rect 28452 3236 28508 3238
rect 28532 3236 28588 3238
rect 28612 3236 28668 3238
rect 29032 2746 29088 2748
rect 29112 2746 29168 2748
rect 29192 2746 29248 2748
rect 29272 2746 29328 2748
rect 29032 2694 29078 2746
rect 29078 2694 29088 2746
rect 29112 2694 29142 2746
rect 29142 2694 29154 2746
rect 29154 2694 29168 2746
rect 29192 2694 29206 2746
rect 29206 2694 29218 2746
rect 29218 2694 29248 2746
rect 29272 2694 29282 2746
rect 29282 2694 29328 2746
rect 29032 2692 29088 2694
rect 29112 2692 29168 2694
rect 29192 2692 29248 2694
rect 29272 2692 29328 2694
rect 33138 9560 33194 9616
rect 31666 9016 31722 9072
rect 31574 7792 31630 7848
rect 33138 7520 33194 7576
rect 33138 6196 33140 6216
rect 33140 6196 33192 6216
rect 33192 6196 33194 6216
rect 33138 6160 33194 6196
rect 31666 5208 31722 5264
rect 33046 4140 33102 4176
rect 33046 4120 33048 4140
rect 33048 4120 33100 4140
rect 33100 4120 33102 4140
rect 31666 1400 31722 1456
rect 33138 2760 33194 2816
<< metal3 >>
rect 0 34098 800 34128
rect 4521 34098 4587 34101
rect 0 34096 4587 34098
rect 0 34040 4526 34096
rect 4582 34040 4587 34096
rect 0 34038 4587 34040
rect 0 34008 800 34038
rect 4521 34035 4587 34038
rect 33133 33418 33199 33421
rect 34168 33418 34968 33448
rect 33133 33416 34968 33418
rect 33133 33360 33138 33416
rect 33194 33360 34968 33416
rect 33133 33358 34968 33360
rect 33133 33355 33199 33358
rect 34168 33328 34968 33358
rect 6942 32128 7258 32129
rect 0 32058 800 32088
rect 6942 32064 6948 32128
rect 7012 32064 7028 32128
rect 7092 32064 7108 32128
rect 7172 32064 7188 32128
rect 7252 32064 7258 32128
rect 6942 32063 7258 32064
rect 14302 32128 14618 32129
rect 14302 32064 14308 32128
rect 14372 32064 14388 32128
rect 14452 32064 14468 32128
rect 14532 32064 14548 32128
rect 14612 32064 14618 32128
rect 14302 32063 14618 32064
rect 21662 32128 21978 32129
rect 21662 32064 21668 32128
rect 21732 32064 21748 32128
rect 21812 32064 21828 32128
rect 21892 32064 21908 32128
rect 21972 32064 21978 32128
rect 21662 32063 21978 32064
rect 29022 32128 29338 32129
rect 29022 32064 29028 32128
rect 29092 32064 29108 32128
rect 29172 32064 29188 32128
rect 29252 32064 29268 32128
rect 29332 32064 29338 32128
rect 29022 32063 29338 32064
rect 2773 32058 2839 32061
rect 0 32056 2839 32058
rect 0 32000 2778 32056
rect 2834 32000 2839 32056
rect 0 31998 2839 32000
rect 0 31968 800 31998
rect 2773 31995 2839 31998
rect 31661 32058 31727 32061
rect 34168 32058 34968 32088
rect 31661 32056 34968 32058
rect 31661 32000 31666 32056
rect 31722 32000 34968 32056
rect 31661 31998 34968 32000
rect 31661 31995 31727 31998
rect 34168 31968 34968 31998
rect 13302 31860 13308 31924
rect 13372 31922 13378 31924
rect 18781 31922 18847 31925
rect 13372 31920 18847 31922
rect 13372 31864 18786 31920
rect 18842 31864 18847 31920
rect 13372 31862 18847 31864
rect 13372 31860 13378 31862
rect 18781 31859 18847 31862
rect 17718 31724 17724 31788
rect 17788 31786 17794 31788
rect 17861 31786 17927 31789
rect 17788 31784 17927 31786
rect 17788 31728 17866 31784
rect 17922 31728 17927 31784
rect 17788 31726 17927 31728
rect 17788 31724 17794 31726
rect 17861 31723 17927 31726
rect 6282 31584 6598 31585
rect 6282 31520 6288 31584
rect 6352 31520 6368 31584
rect 6432 31520 6448 31584
rect 6512 31520 6528 31584
rect 6592 31520 6598 31584
rect 6282 31519 6598 31520
rect 13642 31584 13958 31585
rect 13642 31520 13648 31584
rect 13712 31520 13728 31584
rect 13792 31520 13808 31584
rect 13872 31520 13888 31584
rect 13952 31520 13958 31584
rect 13642 31519 13958 31520
rect 21002 31584 21318 31585
rect 21002 31520 21008 31584
rect 21072 31520 21088 31584
rect 21152 31520 21168 31584
rect 21232 31520 21248 31584
rect 21312 31520 21318 31584
rect 21002 31519 21318 31520
rect 28362 31584 28678 31585
rect 28362 31520 28368 31584
rect 28432 31520 28448 31584
rect 28512 31520 28528 31584
rect 28592 31520 28608 31584
rect 28672 31520 28678 31584
rect 28362 31519 28678 31520
rect 14549 31378 14615 31381
rect 29637 31378 29703 31381
rect 14549 31376 29703 31378
rect 14549 31320 14554 31376
rect 14610 31320 29642 31376
rect 29698 31320 29703 31376
rect 14549 31318 29703 31320
rect 14549 31315 14615 31318
rect 29637 31315 29703 31318
rect 24485 31106 24551 31109
rect 25221 31106 25287 31109
rect 24485 31104 25287 31106
rect 24485 31048 24490 31104
rect 24546 31048 25226 31104
rect 25282 31048 25287 31104
rect 24485 31046 25287 31048
rect 24485 31043 24551 31046
rect 25221 31043 25287 31046
rect 25589 31106 25655 31109
rect 26601 31106 26667 31109
rect 25589 31104 26667 31106
rect 25589 31048 25594 31104
rect 25650 31048 26606 31104
rect 26662 31048 26667 31104
rect 25589 31046 26667 31048
rect 25589 31043 25655 31046
rect 26601 31043 26667 31046
rect 6942 31040 7258 31041
rect 6942 30976 6948 31040
rect 7012 30976 7028 31040
rect 7092 30976 7108 31040
rect 7172 30976 7188 31040
rect 7252 30976 7258 31040
rect 6942 30975 7258 30976
rect 14302 31040 14618 31041
rect 14302 30976 14308 31040
rect 14372 30976 14388 31040
rect 14452 30976 14468 31040
rect 14532 30976 14548 31040
rect 14612 30976 14618 31040
rect 14302 30975 14618 30976
rect 21662 31040 21978 31041
rect 21662 30976 21668 31040
rect 21732 30976 21748 31040
rect 21812 30976 21828 31040
rect 21892 30976 21908 31040
rect 21972 30976 21978 31040
rect 21662 30975 21978 30976
rect 29022 31040 29338 31041
rect 29022 30976 29028 31040
rect 29092 30976 29108 31040
rect 29172 30976 29188 31040
rect 29252 30976 29268 31040
rect 29332 30976 29338 31040
rect 29022 30975 29338 30976
rect 0 30698 800 30728
rect 1301 30698 1367 30701
rect 0 30696 1367 30698
rect 0 30640 1306 30696
rect 1362 30640 1367 30696
rect 0 30638 1367 30640
rect 0 30608 800 30638
rect 1301 30635 1367 30638
rect 33041 30698 33107 30701
rect 34168 30698 34968 30728
rect 33041 30696 34968 30698
rect 33041 30640 33046 30696
rect 33102 30640 34968 30696
rect 33041 30638 34968 30640
rect 33041 30635 33107 30638
rect 34168 30608 34968 30638
rect 6282 30496 6598 30497
rect 6282 30432 6288 30496
rect 6352 30432 6368 30496
rect 6432 30432 6448 30496
rect 6512 30432 6528 30496
rect 6592 30432 6598 30496
rect 6282 30431 6598 30432
rect 13642 30496 13958 30497
rect 13642 30432 13648 30496
rect 13712 30432 13728 30496
rect 13792 30432 13808 30496
rect 13872 30432 13888 30496
rect 13952 30432 13958 30496
rect 13642 30431 13958 30432
rect 21002 30496 21318 30497
rect 21002 30432 21008 30496
rect 21072 30432 21088 30496
rect 21152 30432 21168 30496
rect 21232 30432 21248 30496
rect 21312 30432 21318 30496
rect 21002 30431 21318 30432
rect 28362 30496 28678 30497
rect 28362 30432 28368 30496
rect 28432 30432 28448 30496
rect 28512 30432 28528 30496
rect 28592 30432 28608 30496
rect 28672 30432 28678 30496
rect 28362 30431 28678 30432
rect 25773 30154 25839 30157
rect 26969 30154 27035 30157
rect 25773 30152 27035 30154
rect 25773 30096 25778 30152
rect 25834 30096 26974 30152
rect 27030 30096 27035 30152
rect 25773 30094 27035 30096
rect 25773 30091 25839 30094
rect 26969 30091 27035 30094
rect 6942 29952 7258 29953
rect 6942 29888 6948 29952
rect 7012 29888 7028 29952
rect 7092 29888 7108 29952
rect 7172 29888 7188 29952
rect 7252 29888 7258 29952
rect 6942 29887 7258 29888
rect 14302 29952 14618 29953
rect 14302 29888 14308 29952
rect 14372 29888 14388 29952
rect 14452 29888 14468 29952
rect 14532 29888 14548 29952
rect 14612 29888 14618 29952
rect 14302 29887 14618 29888
rect 21662 29952 21978 29953
rect 21662 29888 21668 29952
rect 21732 29888 21748 29952
rect 21812 29888 21828 29952
rect 21892 29888 21908 29952
rect 21972 29888 21978 29952
rect 21662 29887 21978 29888
rect 29022 29952 29338 29953
rect 29022 29888 29028 29952
rect 29092 29888 29108 29952
rect 29172 29888 29188 29952
rect 29252 29888 29268 29952
rect 29332 29888 29338 29952
rect 29022 29887 29338 29888
rect 6282 29408 6598 29409
rect 6282 29344 6288 29408
rect 6352 29344 6368 29408
rect 6432 29344 6448 29408
rect 6512 29344 6528 29408
rect 6592 29344 6598 29408
rect 6282 29343 6598 29344
rect 13642 29408 13958 29409
rect 13642 29344 13648 29408
rect 13712 29344 13728 29408
rect 13792 29344 13808 29408
rect 13872 29344 13888 29408
rect 13952 29344 13958 29408
rect 13642 29343 13958 29344
rect 21002 29408 21318 29409
rect 21002 29344 21008 29408
rect 21072 29344 21088 29408
rect 21152 29344 21168 29408
rect 21232 29344 21248 29408
rect 21312 29344 21318 29408
rect 21002 29343 21318 29344
rect 28362 29408 28678 29409
rect 28362 29344 28368 29408
rect 28432 29344 28448 29408
rect 28512 29344 28528 29408
rect 28592 29344 28608 29408
rect 28672 29344 28678 29408
rect 28362 29343 28678 29344
rect 6942 28864 7258 28865
rect 6942 28800 6948 28864
rect 7012 28800 7028 28864
rect 7092 28800 7108 28864
rect 7172 28800 7188 28864
rect 7252 28800 7258 28864
rect 6942 28799 7258 28800
rect 14302 28864 14618 28865
rect 14302 28800 14308 28864
rect 14372 28800 14388 28864
rect 14452 28800 14468 28864
rect 14532 28800 14548 28864
rect 14612 28800 14618 28864
rect 14302 28799 14618 28800
rect 21662 28864 21978 28865
rect 21662 28800 21668 28864
rect 21732 28800 21748 28864
rect 21812 28800 21828 28864
rect 21892 28800 21908 28864
rect 21972 28800 21978 28864
rect 21662 28799 21978 28800
rect 29022 28864 29338 28865
rect 29022 28800 29028 28864
rect 29092 28800 29108 28864
rect 29172 28800 29188 28864
rect 29252 28800 29268 28864
rect 29332 28800 29338 28864
rect 29022 28799 29338 28800
rect 0 28658 800 28688
rect 3509 28658 3575 28661
rect 0 28656 3575 28658
rect 0 28600 3514 28656
rect 3570 28600 3575 28656
rect 0 28598 3575 28600
rect 0 28568 800 28598
rect 3509 28595 3575 28598
rect 26141 28658 26207 28661
rect 28901 28658 28967 28661
rect 26141 28656 28967 28658
rect 26141 28600 26146 28656
rect 26202 28600 28906 28656
rect 28962 28600 28967 28656
rect 26141 28598 28967 28600
rect 26141 28595 26207 28598
rect 28901 28595 28967 28598
rect 30373 28658 30439 28661
rect 34168 28658 34968 28688
rect 30373 28656 34968 28658
rect 30373 28600 30378 28656
rect 30434 28600 34968 28656
rect 30373 28598 34968 28600
rect 30373 28595 30439 28598
rect 34168 28568 34968 28598
rect 6282 28320 6598 28321
rect 6282 28256 6288 28320
rect 6352 28256 6368 28320
rect 6432 28256 6448 28320
rect 6512 28256 6528 28320
rect 6592 28256 6598 28320
rect 6282 28255 6598 28256
rect 13642 28320 13958 28321
rect 13642 28256 13648 28320
rect 13712 28256 13728 28320
rect 13792 28256 13808 28320
rect 13872 28256 13888 28320
rect 13952 28256 13958 28320
rect 13642 28255 13958 28256
rect 21002 28320 21318 28321
rect 21002 28256 21008 28320
rect 21072 28256 21088 28320
rect 21152 28256 21168 28320
rect 21232 28256 21248 28320
rect 21312 28256 21318 28320
rect 21002 28255 21318 28256
rect 28362 28320 28678 28321
rect 28362 28256 28368 28320
rect 28432 28256 28448 28320
rect 28512 28256 28528 28320
rect 28592 28256 28608 28320
rect 28672 28256 28678 28320
rect 28362 28255 28678 28256
rect 16573 28116 16639 28117
rect 16573 28112 16620 28116
rect 16684 28114 16690 28116
rect 29453 28114 29519 28117
rect 30189 28114 30255 28117
rect 16573 28056 16578 28112
rect 16573 28052 16620 28056
rect 16684 28054 16730 28114
rect 29453 28112 30255 28114
rect 29453 28056 29458 28112
rect 29514 28056 30194 28112
rect 30250 28056 30255 28112
rect 29453 28054 30255 28056
rect 16684 28052 16690 28054
rect 16573 28051 16639 28052
rect 29453 28051 29519 28054
rect 30189 28051 30255 28054
rect 29361 27978 29427 27981
rect 30741 27978 30807 27981
rect 29361 27976 30807 27978
rect 29361 27920 29366 27976
rect 29422 27920 30746 27976
rect 30802 27920 30807 27976
rect 29361 27918 30807 27920
rect 29361 27915 29427 27918
rect 30741 27915 30807 27918
rect 6942 27776 7258 27777
rect 6942 27712 6948 27776
rect 7012 27712 7028 27776
rect 7092 27712 7108 27776
rect 7172 27712 7188 27776
rect 7252 27712 7258 27776
rect 6942 27711 7258 27712
rect 14302 27776 14618 27777
rect 14302 27712 14308 27776
rect 14372 27712 14388 27776
rect 14452 27712 14468 27776
rect 14532 27712 14548 27776
rect 14612 27712 14618 27776
rect 14302 27711 14618 27712
rect 21662 27776 21978 27777
rect 21662 27712 21668 27776
rect 21732 27712 21748 27776
rect 21812 27712 21828 27776
rect 21892 27712 21908 27776
rect 21972 27712 21978 27776
rect 21662 27711 21978 27712
rect 29022 27776 29338 27777
rect 29022 27712 29028 27776
rect 29092 27712 29108 27776
rect 29172 27712 29188 27776
rect 29252 27712 29268 27776
rect 29332 27712 29338 27776
rect 29022 27711 29338 27712
rect 11053 27708 11119 27709
rect 11053 27704 11100 27708
rect 11164 27706 11170 27708
rect 11053 27648 11058 27704
rect 11053 27644 11100 27648
rect 11164 27646 11210 27706
rect 11164 27644 11170 27646
rect 11053 27643 11119 27644
rect 6821 27570 6887 27573
rect 9213 27570 9279 27573
rect 6821 27568 9279 27570
rect 6821 27512 6826 27568
rect 6882 27512 9218 27568
rect 9274 27512 9279 27568
rect 6821 27510 9279 27512
rect 6821 27507 6887 27510
rect 9213 27507 9279 27510
rect 29545 27434 29611 27437
rect 30097 27434 30163 27437
rect 31109 27434 31175 27437
rect 29545 27432 31175 27434
rect 29545 27376 29550 27432
rect 29606 27376 30102 27432
rect 30158 27376 31114 27432
rect 31170 27376 31175 27432
rect 29545 27374 31175 27376
rect 29545 27371 29611 27374
rect 30097 27371 30163 27374
rect 31109 27371 31175 27374
rect 0 27298 800 27328
rect 1301 27298 1367 27301
rect 0 27296 1367 27298
rect 0 27240 1306 27296
rect 1362 27240 1367 27296
rect 0 27238 1367 27240
rect 0 27208 800 27238
rect 1301 27235 1367 27238
rect 33133 27298 33199 27301
rect 34168 27298 34968 27328
rect 33133 27296 34968 27298
rect 33133 27240 33138 27296
rect 33194 27240 34968 27296
rect 33133 27238 34968 27240
rect 33133 27235 33199 27238
rect 6282 27232 6598 27233
rect 6282 27168 6288 27232
rect 6352 27168 6368 27232
rect 6432 27168 6448 27232
rect 6512 27168 6528 27232
rect 6592 27168 6598 27232
rect 6282 27167 6598 27168
rect 13642 27232 13958 27233
rect 13642 27168 13648 27232
rect 13712 27168 13728 27232
rect 13792 27168 13808 27232
rect 13872 27168 13888 27232
rect 13952 27168 13958 27232
rect 13642 27167 13958 27168
rect 21002 27232 21318 27233
rect 21002 27168 21008 27232
rect 21072 27168 21088 27232
rect 21152 27168 21168 27232
rect 21232 27168 21248 27232
rect 21312 27168 21318 27232
rect 21002 27167 21318 27168
rect 28362 27232 28678 27233
rect 28362 27168 28368 27232
rect 28432 27168 28448 27232
rect 28512 27168 28528 27232
rect 28592 27168 28608 27232
rect 28672 27168 28678 27232
rect 34168 27208 34968 27238
rect 28362 27167 28678 27168
rect 23565 27026 23631 27029
rect 24393 27026 24459 27029
rect 23565 27024 24459 27026
rect 23565 26968 23570 27024
rect 23626 26968 24398 27024
rect 24454 26968 24459 27024
rect 23565 26966 24459 26968
rect 23565 26963 23631 26966
rect 24393 26963 24459 26966
rect 25773 27026 25839 27029
rect 27521 27026 27587 27029
rect 25773 27024 27587 27026
rect 25773 26968 25778 27024
rect 25834 26968 27526 27024
rect 27582 26968 27587 27024
rect 25773 26966 27587 26968
rect 25773 26963 25839 26966
rect 27521 26963 27587 26966
rect 6942 26688 7258 26689
rect 6942 26624 6948 26688
rect 7012 26624 7028 26688
rect 7092 26624 7108 26688
rect 7172 26624 7188 26688
rect 7252 26624 7258 26688
rect 6942 26623 7258 26624
rect 14302 26688 14618 26689
rect 14302 26624 14308 26688
rect 14372 26624 14388 26688
rect 14452 26624 14468 26688
rect 14532 26624 14548 26688
rect 14612 26624 14618 26688
rect 14302 26623 14618 26624
rect 21662 26688 21978 26689
rect 21662 26624 21668 26688
rect 21732 26624 21748 26688
rect 21812 26624 21828 26688
rect 21892 26624 21908 26688
rect 21972 26624 21978 26688
rect 21662 26623 21978 26624
rect 29022 26688 29338 26689
rect 29022 26624 29028 26688
rect 29092 26624 29108 26688
rect 29172 26624 29188 26688
rect 29252 26624 29268 26688
rect 29332 26624 29338 26688
rect 29022 26623 29338 26624
rect 15101 26346 15167 26349
rect 19149 26346 19215 26349
rect 15101 26344 19215 26346
rect 15101 26288 15106 26344
rect 15162 26288 19154 26344
rect 19210 26288 19215 26344
rect 15101 26286 19215 26288
rect 15101 26283 15167 26286
rect 19149 26283 19215 26286
rect 6282 26144 6598 26145
rect 6282 26080 6288 26144
rect 6352 26080 6368 26144
rect 6432 26080 6448 26144
rect 6512 26080 6528 26144
rect 6592 26080 6598 26144
rect 6282 26079 6598 26080
rect 13642 26144 13958 26145
rect 13642 26080 13648 26144
rect 13712 26080 13728 26144
rect 13792 26080 13808 26144
rect 13872 26080 13888 26144
rect 13952 26080 13958 26144
rect 13642 26079 13958 26080
rect 21002 26144 21318 26145
rect 21002 26080 21008 26144
rect 21072 26080 21088 26144
rect 21152 26080 21168 26144
rect 21232 26080 21248 26144
rect 21312 26080 21318 26144
rect 21002 26079 21318 26080
rect 28362 26144 28678 26145
rect 28362 26080 28368 26144
rect 28432 26080 28448 26144
rect 28512 26080 28528 26144
rect 28592 26080 28608 26144
rect 28672 26080 28678 26144
rect 28362 26079 28678 26080
rect 0 25938 800 25968
rect 3233 25938 3299 25941
rect 0 25936 3299 25938
rect 0 25880 3238 25936
rect 3294 25880 3299 25936
rect 0 25878 3299 25880
rect 0 25848 800 25878
rect 3233 25875 3299 25878
rect 11329 25804 11395 25805
rect 11278 25802 11284 25804
rect 11238 25742 11284 25802
rect 11348 25800 11395 25804
rect 11390 25744 11395 25800
rect 11278 25740 11284 25742
rect 11348 25740 11395 25744
rect 11329 25739 11395 25740
rect 6942 25600 7258 25601
rect 6942 25536 6948 25600
rect 7012 25536 7028 25600
rect 7092 25536 7108 25600
rect 7172 25536 7188 25600
rect 7252 25536 7258 25600
rect 6942 25535 7258 25536
rect 14302 25600 14618 25601
rect 14302 25536 14308 25600
rect 14372 25536 14388 25600
rect 14452 25536 14468 25600
rect 14532 25536 14548 25600
rect 14612 25536 14618 25600
rect 14302 25535 14618 25536
rect 21662 25600 21978 25601
rect 21662 25536 21668 25600
rect 21732 25536 21748 25600
rect 21812 25536 21828 25600
rect 21892 25536 21908 25600
rect 21972 25536 21978 25600
rect 21662 25535 21978 25536
rect 29022 25600 29338 25601
rect 29022 25536 29028 25600
rect 29092 25536 29108 25600
rect 29172 25536 29188 25600
rect 29252 25536 29268 25600
rect 29332 25536 29338 25600
rect 29022 25535 29338 25536
rect 33133 25258 33199 25261
rect 34168 25258 34968 25288
rect 33133 25256 34968 25258
rect 33133 25200 33138 25256
rect 33194 25200 34968 25256
rect 33133 25198 34968 25200
rect 33133 25195 33199 25198
rect 34168 25168 34968 25198
rect 6282 25056 6598 25057
rect 6282 24992 6288 25056
rect 6352 24992 6368 25056
rect 6432 24992 6448 25056
rect 6512 24992 6528 25056
rect 6592 24992 6598 25056
rect 6282 24991 6598 24992
rect 13642 25056 13958 25057
rect 13642 24992 13648 25056
rect 13712 24992 13728 25056
rect 13792 24992 13808 25056
rect 13872 24992 13888 25056
rect 13952 24992 13958 25056
rect 13642 24991 13958 24992
rect 21002 25056 21318 25057
rect 21002 24992 21008 25056
rect 21072 24992 21088 25056
rect 21152 24992 21168 25056
rect 21232 24992 21248 25056
rect 21312 24992 21318 25056
rect 21002 24991 21318 24992
rect 28362 25056 28678 25057
rect 28362 24992 28368 25056
rect 28432 24992 28448 25056
rect 28512 24992 28528 25056
rect 28592 24992 28608 25056
rect 28672 24992 28678 25056
rect 28362 24991 28678 24992
rect 9857 24714 9923 24717
rect 12249 24714 12315 24717
rect 9857 24712 12315 24714
rect 9857 24656 9862 24712
rect 9918 24656 12254 24712
rect 12310 24656 12315 24712
rect 9857 24654 12315 24656
rect 9857 24651 9923 24654
rect 12249 24651 12315 24654
rect 6942 24512 7258 24513
rect 6942 24448 6948 24512
rect 7012 24448 7028 24512
rect 7092 24448 7108 24512
rect 7172 24448 7188 24512
rect 7252 24448 7258 24512
rect 6942 24447 7258 24448
rect 14302 24512 14618 24513
rect 14302 24448 14308 24512
rect 14372 24448 14388 24512
rect 14452 24448 14468 24512
rect 14532 24448 14548 24512
rect 14612 24448 14618 24512
rect 14302 24447 14618 24448
rect 21662 24512 21978 24513
rect 21662 24448 21668 24512
rect 21732 24448 21748 24512
rect 21812 24448 21828 24512
rect 21892 24448 21908 24512
rect 21972 24448 21978 24512
rect 21662 24447 21978 24448
rect 29022 24512 29338 24513
rect 29022 24448 29028 24512
rect 29092 24448 29108 24512
rect 29172 24448 29188 24512
rect 29252 24448 29268 24512
rect 29332 24448 29338 24512
rect 29022 24447 29338 24448
rect 11053 24170 11119 24173
rect 11789 24170 11855 24173
rect 15193 24170 15259 24173
rect 11053 24168 15259 24170
rect 11053 24112 11058 24168
rect 11114 24112 11794 24168
rect 11850 24112 15198 24168
rect 15254 24112 15259 24168
rect 11053 24110 15259 24112
rect 11053 24107 11119 24110
rect 11789 24107 11855 24110
rect 15193 24107 15259 24110
rect 6282 23968 6598 23969
rect 0 23898 800 23928
rect 6282 23904 6288 23968
rect 6352 23904 6368 23968
rect 6432 23904 6448 23968
rect 6512 23904 6528 23968
rect 6592 23904 6598 23968
rect 6282 23903 6598 23904
rect 13642 23968 13958 23969
rect 13642 23904 13648 23968
rect 13712 23904 13728 23968
rect 13792 23904 13808 23968
rect 13872 23904 13888 23968
rect 13952 23904 13958 23968
rect 13642 23903 13958 23904
rect 21002 23968 21318 23969
rect 21002 23904 21008 23968
rect 21072 23904 21088 23968
rect 21152 23904 21168 23968
rect 21232 23904 21248 23968
rect 21312 23904 21318 23968
rect 21002 23903 21318 23904
rect 28362 23968 28678 23969
rect 28362 23904 28368 23968
rect 28432 23904 28448 23968
rect 28512 23904 28528 23968
rect 28592 23904 28608 23968
rect 28672 23904 28678 23968
rect 28362 23903 28678 23904
rect 1301 23898 1367 23901
rect 0 23896 1367 23898
rect 0 23840 1306 23896
rect 1362 23840 1367 23896
rect 0 23838 1367 23840
rect 0 23808 800 23838
rect 1301 23835 1367 23838
rect 33133 23898 33199 23901
rect 34168 23898 34968 23928
rect 33133 23896 34968 23898
rect 33133 23840 33138 23896
rect 33194 23840 34968 23896
rect 33133 23838 34968 23840
rect 33133 23835 33199 23838
rect 34168 23808 34968 23838
rect 11605 23762 11671 23765
rect 13118 23762 13124 23764
rect 11605 23760 13124 23762
rect 11605 23704 11610 23760
rect 11666 23704 13124 23760
rect 11605 23702 13124 23704
rect 11605 23699 11671 23702
rect 13118 23700 13124 23702
rect 13188 23762 13194 23764
rect 16113 23762 16179 23765
rect 13188 23760 16179 23762
rect 13188 23704 16118 23760
rect 16174 23704 16179 23760
rect 13188 23702 16179 23704
rect 13188 23700 13194 23702
rect 16113 23699 16179 23702
rect 25497 23626 25563 23629
rect 26785 23626 26851 23629
rect 25497 23624 26851 23626
rect 25497 23568 25502 23624
rect 25558 23568 26790 23624
rect 26846 23568 26851 23624
rect 25497 23566 26851 23568
rect 25497 23563 25563 23566
rect 26785 23563 26851 23566
rect 6942 23424 7258 23425
rect 6942 23360 6948 23424
rect 7012 23360 7028 23424
rect 7092 23360 7108 23424
rect 7172 23360 7188 23424
rect 7252 23360 7258 23424
rect 6942 23359 7258 23360
rect 14302 23424 14618 23425
rect 14302 23360 14308 23424
rect 14372 23360 14388 23424
rect 14452 23360 14468 23424
rect 14532 23360 14548 23424
rect 14612 23360 14618 23424
rect 14302 23359 14618 23360
rect 21662 23424 21978 23425
rect 21662 23360 21668 23424
rect 21732 23360 21748 23424
rect 21812 23360 21828 23424
rect 21892 23360 21908 23424
rect 21972 23360 21978 23424
rect 21662 23359 21978 23360
rect 29022 23424 29338 23425
rect 29022 23360 29028 23424
rect 29092 23360 29108 23424
rect 29172 23360 29188 23424
rect 29252 23360 29268 23424
rect 29332 23360 29338 23424
rect 29022 23359 29338 23360
rect 24577 23354 24643 23357
rect 26049 23354 26115 23357
rect 27245 23354 27311 23357
rect 24577 23352 27311 23354
rect 24577 23296 24582 23352
rect 24638 23296 26054 23352
rect 26110 23296 27250 23352
rect 27306 23296 27311 23352
rect 24577 23294 27311 23296
rect 24577 23291 24643 23294
rect 26049 23291 26115 23294
rect 27245 23291 27311 23294
rect 9949 23218 10015 23221
rect 14365 23218 14431 23221
rect 9949 23216 14431 23218
rect 9949 23160 9954 23216
rect 10010 23160 14370 23216
rect 14426 23160 14431 23216
rect 9949 23158 14431 23160
rect 9949 23155 10015 23158
rect 14365 23155 14431 23158
rect 13537 23082 13603 23085
rect 18137 23082 18203 23085
rect 13537 23080 18203 23082
rect 13537 23024 13542 23080
rect 13598 23024 18142 23080
rect 18198 23024 18203 23080
rect 13537 23022 18203 23024
rect 13537 23019 13603 23022
rect 18137 23019 18203 23022
rect 6282 22880 6598 22881
rect 6282 22816 6288 22880
rect 6352 22816 6368 22880
rect 6432 22816 6448 22880
rect 6512 22816 6528 22880
rect 6592 22816 6598 22880
rect 6282 22815 6598 22816
rect 13642 22880 13958 22881
rect 13642 22816 13648 22880
rect 13712 22816 13728 22880
rect 13792 22816 13808 22880
rect 13872 22816 13888 22880
rect 13952 22816 13958 22880
rect 13642 22815 13958 22816
rect 21002 22880 21318 22881
rect 21002 22816 21008 22880
rect 21072 22816 21088 22880
rect 21152 22816 21168 22880
rect 21232 22816 21248 22880
rect 21312 22816 21318 22880
rect 21002 22815 21318 22816
rect 28362 22880 28678 22881
rect 28362 22816 28368 22880
rect 28432 22816 28448 22880
rect 28512 22816 28528 22880
rect 28592 22816 28608 22880
rect 28672 22816 28678 22880
rect 28362 22815 28678 22816
rect 21541 22674 21607 22677
rect 26049 22674 26115 22677
rect 21541 22672 26115 22674
rect 21541 22616 21546 22672
rect 21602 22616 26054 22672
rect 26110 22616 26115 22672
rect 21541 22614 26115 22616
rect 21541 22611 21607 22614
rect 26049 22611 26115 22614
rect 0 22538 800 22568
rect 1301 22538 1367 22541
rect 0 22536 1367 22538
rect 0 22480 1306 22536
rect 1362 22480 1367 22536
rect 0 22478 1367 22480
rect 0 22448 800 22478
rect 1301 22475 1367 22478
rect 12157 22538 12223 22541
rect 14457 22538 14523 22541
rect 12157 22536 14523 22538
rect 12157 22480 12162 22536
rect 12218 22480 14462 22536
rect 14518 22480 14523 22536
rect 12157 22478 14523 22480
rect 12157 22475 12223 22478
rect 14457 22475 14523 22478
rect 21633 22538 21699 22541
rect 26693 22538 26759 22541
rect 27429 22538 27495 22541
rect 21633 22536 27495 22538
rect 21633 22480 21638 22536
rect 21694 22480 26698 22536
rect 26754 22480 27434 22536
rect 27490 22480 27495 22536
rect 21633 22478 27495 22480
rect 21633 22475 21699 22478
rect 26693 22475 26759 22478
rect 27429 22475 27495 22478
rect 31661 22538 31727 22541
rect 34168 22538 34968 22568
rect 31661 22536 34968 22538
rect 31661 22480 31666 22536
rect 31722 22480 34968 22536
rect 31661 22478 34968 22480
rect 31661 22475 31727 22478
rect 34168 22448 34968 22478
rect 25313 22402 25379 22405
rect 26969 22402 27035 22405
rect 25313 22400 27035 22402
rect 25313 22344 25318 22400
rect 25374 22344 26974 22400
rect 27030 22344 27035 22400
rect 25313 22342 27035 22344
rect 25313 22339 25379 22342
rect 26969 22339 27035 22342
rect 6942 22336 7258 22337
rect 6942 22272 6948 22336
rect 7012 22272 7028 22336
rect 7092 22272 7108 22336
rect 7172 22272 7188 22336
rect 7252 22272 7258 22336
rect 6942 22271 7258 22272
rect 14302 22336 14618 22337
rect 14302 22272 14308 22336
rect 14372 22272 14388 22336
rect 14452 22272 14468 22336
rect 14532 22272 14548 22336
rect 14612 22272 14618 22336
rect 14302 22271 14618 22272
rect 21662 22336 21978 22337
rect 21662 22272 21668 22336
rect 21732 22272 21748 22336
rect 21812 22272 21828 22336
rect 21892 22272 21908 22336
rect 21972 22272 21978 22336
rect 21662 22271 21978 22272
rect 29022 22336 29338 22337
rect 29022 22272 29028 22336
rect 29092 22272 29108 22336
rect 29172 22272 29188 22336
rect 29252 22272 29268 22336
rect 29332 22272 29338 22336
rect 29022 22271 29338 22272
rect 15101 22266 15167 22269
rect 16389 22266 16455 22269
rect 15101 22264 16455 22266
rect 15101 22208 15106 22264
rect 15162 22208 16394 22264
rect 16450 22208 16455 22264
rect 15101 22206 16455 22208
rect 15101 22203 15167 22206
rect 16389 22203 16455 22206
rect 24669 22130 24735 22133
rect 27337 22130 27403 22133
rect 24669 22128 27403 22130
rect 24669 22072 24674 22128
rect 24730 22072 27342 22128
rect 27398 22072 27403 22128
rect 24669 22070 27403 22072
rect 24669 22067 24735 22070
rect 27337 22067 27403 22070
rect 6282 21792 6598 21793
rect 6282 21728 6288 21792
rect 6352 21728 6368 21792
rect 6432 21728 6448 21792
rect 6512 21728 6528 21792
rect 6592 21728 6598 21792
rect 6282 21727 6598 21728
rect 13642 21792 13958 21793
rect 13642 21728 13648 21792
rect 13712 21728 13728 21792
rect 13792 21728 13808 21792
rect 13872 21728 13888 21792
rect 13952 21728 13958 21792
rect 13642 21727 13958 21728
rect 21002 21792 21318 21793
rect 21002 21728 21008 21792
rect 21072 21728 21088 21792
rect 21152 21728 21168 21792
rect 21232 21728 21248 21792
rect 21312 21728 21318 21792
rect 21002 21727 21318 21728
rect 28362 21792 28678 21793
rect 28362 21728 28368 21792
rect 28432 21728 28448 21792
rect 28512 21728 28528 21792
rect 28592 21728 28608 21792
rect 28672 21728 28678 21792
rect 28362 21727 28678 21728
rect 6942 21248 7258 21249
rect 6942 21184 6948 21248
rect 7012 21184 7028 21248
rect 7092 21184 7108 21248
rect 7172 21184 7188 21248
rect 7252 21184 7258 21248
rect 6942 21183 7258 21184
rect 14302 21248 14618 21249
rect 14302 21184 14308 21248
rect 14372 21184 14388 21248
rect 14452 21184 14468 21248
rect 14532 21184 14548 21248
rect 14612 21184 14618 21248
rect 14302 21183 14618 21184
rect 21662 21248 21978 21249
rect 21662 21184 21668 21248
rect 21732 21184 21748 21248
rect 21812 21184 21828 21248
rect 21892 21184 21908 21248
rect 21972 21184 21978 21248
rect 21662 21183 21978 21184
rect 29022 21248 29338 21249
rect 29022 21184 29028 21248
rect 29092 21184 29108 21248
rect 29172 21184 29188 21248
rect 29252 21184 29268 21248
rect 29332 21184 29338 21248
rect 29022 21183 29338 21184
rect 15285 21178 15351 21181
rect 16665 21178 16731 21181
rect 15285 21176 16731 21178
rect 15285 21120 15290 21176
rect 15346 21120 16670 21176
rect 16726 21120 16731 21176
rect 15285 21118 16731 21120
rect 15285 21115 15351 21118
rect 16665 21115 16731 21118
rect 3325 21042 3391 21045
rect 29729 21042 29795 21045
rect 3325 21040 29795 21042
rect 3325 20984 3330 21040
rect 3386 20984 29734 21040
rect 29790 20984 29795 21040
rect 3325 20982 29795 20984
rect 3325 20979 3391 20982
rect 29729 20979 29795 20982
rect 13813 20906 13879 20909
rect 24526 20906 24532 20908
rect 13813 20904 24532 20906
rect 13813 20848 13818 20904
rect 13874 20848 24532 20904
rect 13813 20846 24532 20848
rect 13813 20843 13879 20846
rect 24526 20844 24532 20846
rect 24596 20844 24602 20908
rect 14733 20772 14799 20773
rect 14733 20770 14780 20772
rect 14688 20768 14780 20770
rect 14688 20712 14738 20768
rect 14688 20710 14780 20712
rect 14733 20708 14780 20710
rect 14844 20708 14850 20772
rect 16021 20770 16087 20773
rect 16430 20770 16436 20772
rect 16021 20768 16436 20770
rect 16021 20712 16026 20768
rect 16082 20712 16436 20768
rect 16021 20710 16436 20712
rect 14733 20707 14799 20708
rect 16021 20707 16087 20710
rect 16430 20708 16436 20710
rect 16500 20708 16506 20772
rect 6282 20704 6598 20705
rect 6282 20640 6288 20704
rect 6352 20640 6368 20704
rect 6432 20640 6448 20704
rect 6512 20640 6528 20704
rect 6592 20640 6598 20704
rect 6282 20639 6598 20640
rect 13642 20704 13958 20705
rect 13642 20640 13648 20704
rect 13712 20640 13728 20704
rect 13792 20640 13808 20704
rect 13872 20640 13888 20704
rect 13952 20640 13958 20704
rect 13642 20639 13958 20640
rect 21002 20704 21318 20705
rect 21002 20640 21008 20704
rect 21072 20640 21088 20704
rect 21152 20640 21168 20704
rect 21232 20640 21248 20704
rect 21312 20640 21318 20704
rect 21002 20639 21318 20640
rect 28362 20704 28678 20705
rect 28362 20640 28368 20704
rect 28432 20640 28448 20704
rect 28512 20640 28528 20704
rect 28592 20640 28608 20704
rect 28672 20640 28678 20704
rect 28362 20639 28678 20640
rect 0 20498 800 20528
rect 3049 20498 3115 20501
rect 0 20496 3115 20498
rect 0 20440 3054 20496
rect 3110 20440 3115 20496
rect 0 20438 3115 20440
rect 0 20408 800 20438
rect 3049 20435 3115 20438
rect 9673 20498 9739 20501
rect 11278 20498 11284 20500
rect 9673 20496 11284 20498
rect 9673 20440 9678 20496
rect 9734 20440 11284 20496
rect 9673 20438 11284 20440
rect 9673 20435 9739 20438
rect 11278 20436 11284 20438
rect 11348 20436 11354 20500
rect 20897 20498 20963 20501
rect 28073 20498 28139 20501
rect 20897 20496 28139 20498
rect 20897 20440 20902 20496
rect 20958 20440 28078 20496
rect 28134 20440 28139 20496
rect 20897 20438 28139 20440
rect 20897 20435 20963 20438
rect 28073 20435 28139 20438
rect 33041 20498 33107 20501
rect 34168 20498 34968 20528
rect 33041 20496 34968 20498
rect 33041 20440 33046 20496
rect 33102 20440 34968 20496
rect 33041 20438 34968 20440
rect 33041 20435 33107 20438
rect 34168 20408 34968 20438
rect 20437 20362 20503 20365
rect 24393 20362 24459 20365
rect 20437 20360 24459 20362
rect 20437 20304 20442 20360
rect 20498 20304 24398 20360
rect 24454 20304 24459 20360
rect 20437 20302 24459 20304
rect 20437 20299 20503 20302
rect 24393 20299 24459 20302
rect 6942 20160 7258 20161
rect 6942 20096 6948 20160
rect 7012 20096 7028 20160
rect 7092 20096 7108 20160
rect 7172 20096 7188 20160
rect 7252 20096 7258 20160
rect 6942 20095 7258 20096
rect 14302 20160 14618 20161
rect 14302 20096 14308 20160
rect 14372 20096 14388 20160
rect 14452 20096 14468 20160
rect 14532 20096 14548 20160
rect 14612 20096 14618 20160
rect 14302 20095 14618 20096
rect 21662 20160 21978 20161
rect 21662 20096 21668 20160
rect 21732 20096 21748 20160
rect 21812 20096 21828 20160
rect 21892 20096 21908 20160
rect 21972 20096 21978 20160
rect 21662 20095 21978 20096
rect 29022 20160 29338 20161
rect 29022 20096 29028 20160
rect 29092 20096 29108 20160
rect 29172 20096 29188 20160
rect 29252 20096 29268 20160
rect 29332 20096 29338 20160
rect 29022 20095 29338 20096
rect 11605 19954 11671 19957
rect 15193 19954 15259 19957
rect 11605 19952 15259 19954
rect 11605 19896 11610 19952
rect 11666 19896 15198 19952
rect 15254 19896 15259 19952
rect 11605 19894 15259 19896
rect 11605 19891 11671 19894
rect 15193 19891 15259 19894
rect 15326 19892 15332 19956
rect 15396 19954 15402 19956
rect 15653 19954 15719 19957
rect 15396 19952 15719 19954
rect 15396 19896 15658 19952
rect 15714 19896 15719 19952
rect 15396 19894 15719 19896
rect 15396 19892 15402 19894
rect 15653 19891 15719 19894
rect 15929 19954 15995 19957
rect 18597 19954 18663 19957
rect 30649 19954 30715 19957
rect 15929 19952 30715 19954
rect 15929 19896 15934 19952
rect 15990 19896 18602 19952
rect 18658 19896 30654 19952
rect 30710 19896 30715 19952
rect 15929 19894 30715 19896
rect 15929 19891 15995 19894
rect 18597 19891 18663 19894
rect 30649 19891 30715 19894
rect 12985 19818 13051 19821
rect 17585 19818 17651 19821
rect 12985 19816 17651 19818
rect 12985 19760 12990 19816
rect 13046 19760 17590 19816
rect 17646 19760 17651 19816
rect 12985 19758 17651 19760
rect 12985 19755 13051 19758
rect 17585 19755 17651 19758
rect 18873 19818 18939 19821
rect 30649 19818 30715 19821
rect 18873 19816 30715 19818
rect 18873 19760 18878 19816
rect 18934 19760 30654 19816
rect 30710 19760 30715 19816
rect 18873 19758 30715 19760
rect 18873 19755 18939 19758
rect 30649 19755 30715 19758
rect 23749 19682 23815 19685
rect 25313 19682 25379 19685
rect 23749 19680 25379 19682
rect 23749 19624 23754 19680
rect 23810 19624 25318 19680
rect 25374 19624 25379 19680
rect 23749 19622 25379 19624
rect 23749 19619 23815 19622
rect 25313 19619 25379 19622
rect 6282 19616 6598 19617
rect 6282 19552 6288 19616
rect 6352 19552 6368 19616
rect 6432 19552 6448 19616
rect 6512 19552 6528 19616
rect 6592 19552 6598 19616
rect 6282 19551 6598 19552
rect 13642 19616 13958 19617
rect 13642 19552 13648 19616
rect 13712 19552 13728 19616
rect 13792 19552 13808 19616
rect 13872 19552 13888 19616
rect 13952 19552 13958 19616
rect 13642 19551 13958 19552
rect 21002 19616 21318 19617
rect 21002 19552 21008 19616
rect 21072 19552 21088 19616
rect 21152 19552 21168 19616
rect 21232 19552 21248 19616
rect 21312 19552 21318 19616
rect 21002 19551 21318 19552
rect 28362 19616 28678 19617
rect 28362 19552 28368 19616
rect 28432 19552 28448 19616
rect 28512 19552 28528 19616
rect 28592 19552 28608 19616
rect 28672 19552 28678 19616
rect 28362 19551 28678 19552
rect 12934 19348 12940 19412
rect 13004 19410 13010 19412
rect 13077 19410 13143 19413
rect 13004 19408 13143 19410
rect 13004 19352 13082 19408
rect 13138 19352 13143 19408
rect 13004 19350 13143 19352
rect 13004 19348 13010 19350
rect 13077 19347 13143 19350
rect 13537 19410 13603 19413
rect 14733 19410 14799 19413
rect 13537 19408 14799 19410
rect 13537 19352 13542 19408
rect 13598 19352 14738 19408
rect 14794 19352 14799 19408
rect 13537 19350 14799 19352
rect 13537 19347 13603 19350
rect 14733 19347 14799 19350
rect 9857 19274 9923 19277
rect 12198 19274 12204 19276
rect 9857 19272 12204 19274
rect 9857 19216 9862 19272
rect 9918 19216 12204 19272
rect 9857 19214 12204 19216
rect 9857 19211 9923 19214
rect 12198 19212 12204 19214
rect 12268 19274 12274 19276
rect 14549 19274 14615 19277
rect 12268 19272 14615 19274
rect 12268 19216 14554 19272
rect 14610 19216 14615 19272
rect 12268 19214 14615 19216
rect 12268 19212 12274 19214
rect 14549 19211 14615 19214
rect 14733 19274 14799 19277
rect 14733 19272 14842 19274
rect 14733 19216 14738 19272
rect 14794 19216 14842 19272
rect 14733 19211 14842 19216
rect 0 19138 800 19168
rect 1301 19138 1367 19141
rect 0 19136 1367 19138
rect 0 19080 1306 19136
rect 1362 19080 1367 19136
rect 0 19078 1367 19080
rect 0 19048 800 19078
rect 1301 19075 1367 19078
rect 6942 19072 7258 19073
rect 6942 19008 6948 19072
rect 7012 19008 7028 19072
rect 7092 19008 7108 19072
rect 7172 19008 7188 19072
rect 7252 19008 7258 19072
rect 6942 19007 7258 19008
rect 14302 19072 14618 19073
rect 14302 19008 14308 19072
rect 14372 19008 14388 19072
rect 14452 19008 14468 19072
rect 14532 19008 14548 19072
rect 14612 19008 14618 19072
rect 14302 19007 14618 19008
rect 14365 18866 14431 18869
rect 14782 18866 14842 19211
rect 33133 19138 33199 19141
rect 34168 19138 34968 19168
rect 33133 19136 34968 19138
rect 33133 19080 33138 19136
rect 33194 19080 34968 19136
rect 33133 19078 34968 19080
rect 33133 19075 33199 19078
rect 21662 19072 21978 19073
rect 21662 19008 21668 19072
rect 21732 19008 21748 19072
rect 21812 19008 21828 19072
rect 21892 19008 21908 19072
rect 21972 19008 21978 19072
rect 21662 19007 21978 19008
rect 29022 19072 29338 19073
rect 29022 19008 29028 19072
rect 29092 19008 29108 19072
rect 29172 19008 29188 19072
rect 29252 19008 29268 19072
rect 29332 19008 29338 19072
rect 34168 19048 34968 19078
rect 29022 19007 29338 19008
rect 14365 18864 14842 18866
rect 14365 18808 14370 18864
rect 14426 18808 14842 18864
rect 14365 18806 14842 18808
rect 21357 18866 21423 18869
rect 26877 18866 26943 18869
rect 21357 18864 26943 18866
rect 21357 18808 21362 18864
rect 21418 18808 26882 18864
rect 26938 18808 26943 18864
rect 21357 18806 26943 18808
rect 14365 18803 14431 18806
rect 21357 18803 21423 18806
rect 26877 18803 26943 18806
rect 21357 18730 21423 18733
rect 28809 18730 28875 18733
rect 21357 18728 28875 18730
rect 21357 18672 21362 18728
rect 21418 18672 28814 18728
rect 28870 18672 28875 18728
rect 21357 18670 28875 18672
rect 21357 18667 21423 18670
rect 28809 18667 28875 18670
rect 6282 18528 6598 18529
rect 6282 18464 6288 18528
rect 6352 18464 6368 18528
rect 6432 18464 6448 18528
rect 6512 18464 6528 18528
rect 6592 18464 6598 18528
rect 6282 18463 6598 18464
rect 13642 18528 13958 18529
rect 13642 18464 13648 18528
rect 13712 18464 13728 18528
rect 13792 18464 13808 18528
rect 13872 18464 13888 18528
rect 13952 18464 13958 18528
rect 13642 18463 13958 18464
rect 21002 18528 21318 18529
rect 21002 18464 21008 18528
rect 21072 18464 21088 18528
rect 21152 18464 21168 18528
rect 21232 18464 21248 18528
rect 21312 18464 21318 18528
rect 21002 18463 21318 18464
rect 28362 18528 28678 18529
rect 28362 18464 28368 18528
rect 28432 18464 28448 18528
rect 28512 18464 28528 18528
rect 28592 18464 28608 18528
rect 28672 18464 28678 18528
rect 28362 18463 28678 18464
rect 19609 18458 19675 18461
rect 20805 18458 20871 18461
rect 19609 18456 20871 18458
rect 19609 18400 19614 18456
rect 19670 18400 20810 18456
rect 20866 18400 20871 18456
rect 19609 18398 20871 18400
rect 19609 18395 19675 18398
rect 20805 18395 20871 18398
rect 15101 18322 15167 18325
rect 15837 18322 15903 18325
rect 15101 18320 15903 18322
rect 15101 18264 15106 18320
rect 15162 18264 15842 18320
rect 15898 18264 15903 18320
rect 15101 18262 15903 18264
rect 15101 18259 15167 18262
rect 15837 18259 15903 18262
rect 19517 18322 19583 18325
rect 20437 18322 20503 18325
rect 19517 18320 20503 18322
rect 19517 18264 19522 18320
rect 19578 18264 20442 18320
rect 20498 18264 20503 18320
rect 19517 18262 20503 18264
rect 19517 18259 19583 18262
rect 20437 18259 20503 18262
rect 14365 18186 14431 18189
rect 15745 18186 15811 18189
rect 14365 18184 15811 18186
rect 14365 18128 14370 18184
rect 14426 18128 15750 18184
rect 15806 18128 15811 18184
rect 14365 18126 15811 18128
rect 14365 18123 14431 18126
rect 15745 18123 15811 18126
rect 19793 18186 19859 18189
rect 20621 18186 20687 18189
rect 19793 18184 20687 18186
rect 19793 18128 19798 18184
rect 19854 18128 20626 18184
rect 20682 18128 20687 18184
rect 19793 18126 20687 18128
rect 19793 18123 19859 18126
rect 20621 18123 20687 18126
rect 16849 18050 16915 18053
rect 17401 18050 17467 18053
rect 19057 18050 19123 18053
rect 16849 18048 19123 18050
rect 16849 17992 16854 18048
rect 16910 17992 17406 18048
rect 17462 17992 19062 18048
rect 19118 17992 19123 18048
rect 16849 17990 19123 17992
rect 16849 17987 16915 17990
rect 17401 17987 17467 17990
rect 19057 17987 19123 17990
rect 6942 17984 7258 17985
rect 6942 17920 6948 17984
rect 7012 17920 7028 17984
rect 7092 17920 7108 17984
rect 7172 17920 7188 17984
rect 7252 17920 7258 17984
rect 6942 17919 7258 17920
rect 14302 17984 14618 17985
rect 14302 17920 14308 17984
rect 14372 17920 14388 17984
rect 14452 17920 14468 17984
rect 14532 17920 14548 17984
rect 14612 17920 14618 17984
rect 14302 17919 14618 17920
rect 21662 17984 21978 17985
rect 21662 17920 21668 17984
rect 21732 17920 21748 17984
rect 21812 17920 21828 17984
rect 21892 17920 21908 17984
rect 21972 17920 21978 17984
rect 21662 17919 21978 17920
rect 29022 17984 29338 17985
rect 29022 17920 29028 17984
rect 29092 17920 29108 17984
rect 29172 17920 29188 17984
rect 29252 17920 29268 17984
rect 29332 17920 29338 17984
rect 29022 17919 29338 17920
rect 16481 17914 16547 17917
rect 18965 17914 19031 17917
rect 16481 17912 19031 17914
rect 16481 17856 16486 17912
rect 16542 17856 18970 17912
rect 19026 17856 19031 17912
rect 16481 17854 19031 17856
rect 16481 17851 16547 17854
rect 18965 17851 19031 17854
rect 0 17778 800 17808
rect 4061 17778 4127 17781
rect 0 17776 4127 17778
rect 0 17720 4066 17776
rect 4122 17720 4127 17776
rect 0 17718 4127 17720
rect 0 17688 800 17718
rect 4061 17715 4127 17718
rect 13997 17778 14063 17781
rect 18873 17778 18939 17781
rect 13997 17776 18939 17778
rect 13997 17720 14002 17776
rect 14058 17720 18878 17776
rect 18934 17720 18939 17776
rect 13997 17718 18939 17720
rect 13997 17715 14106 17718
rect 18873 17715 18939 17718
rect 6282 17440 6598 17441
rect 6282 17376 6288 17440
rect 6352 17376 6368 17440
rect 6432 17376 6448 17440
rect 6512 17376 6528 17440
rect 6592 17376 6598 17440
rect 6282 17375 6598 17376
rect 13642 17440 13958 17441
rect 13642 17376 13648 17440
rect 13712 17376 13728 17440
rect 13792 17376 13808 17440
rect 13872 17376 13888 17440
rect 13952 17376 13958 17440
rect 13642 17375 13958 17376
rect 14046 17373 14106 17715
rect 21002 17440 21318 17441
rect 21002 17376 21008 17440
rect 21072 17376 21088 17440
rect 21152 17376 21168 17440
rect 21232 17376 21248 17440
rect 21312 17376 21318 17440
rect 21002 17375 21318 17376
rect 28362 17440 28678 17441
rect 28362 17376 28368 17440
rect 28432 17376 28448 17440
rect 28512 17376 28528 17440
rect 28592 17376 28608 17440
rect 28672 17376 28678 17440
rect 28362 17375 28678 17376
rect 14046 17368 14155 17373
rect 14046 17312 14094 17368
rect 14150 17312 14155 17368
rect 14046 17310 14155 17312
rect 14089 17307 14155 17310
rect 14549 17370 14615 17373
rect 15009 17370 15075 17373
rect 14549 17368 15075 17370
rect 14549 17312 14554 17368
rect 14610 17312 15014 17368
rect 15070 17312 15075 17368
rect 14549 17310 15075 17312
rect 14549 17307 14615 17310
rect 15009 17307 15075 17310
rect 13077 17234 13143 17237
rect 15285 17234 15351 17237
rect 17769 17234 17835 17237
rect 13077 17232 17835 17234
rect 13077 17176 13082 17232
rect 13138 17176 15290 17232
rect 15346 17176 17774 17232
rect 17830 17176 17835 17232
rect 13077 17174 17835 17176
rect 13077 17171 13143 17174
rect 15285 17171 15351 17174
rect 17769 17171 17835 17174
rect 13353 17098 13419 17101
rect 16481 17098 16547 17101
rect 13353 17096 16547 17098
rect 13353 17040 13358 17096
rect 13414 17040 16486 17096
rect 16542 17040 16547 17096
rect 13353 17038 16547 17040
rect 13353 17035 13419 17038
rect 16481 17035 16547 17038
rect 17033 17098 17099 17101
rect 18321 17098 18387 17101
rect 17033 17096 18387 17098
rect 17033 17040 17038 17096
rect 17094 17040 18326 17096
rect 18382 17040 18387 17096
rect 17033 17038 18387 17040
rect 17033 17035 17099 17038
rect 18321 17035 18387 17038
rect 33133 17098 33199 17101
rect 34168 17098 34968 17128
rect 33133 17096 34968 17098
rect 33133 17040 33138 17096
rect 33194 17040 34968 17096
rect 33133 17038 34968 17040
rect 33133 17035 33199 17038
rect 34168 17008 34968 17038
rect 6942 16896 7258 16897
rect 6942 16832 6948 16896
rect 7012 16832 7028 16896
rect 7092 16832 7108 16896
rect 7172 16832 7188 16896
rect 7252 16832 7258 16896
rect 6942 16831 7258 16832
rect 14302 16896 14618 16897
rect 14302 16832 14308 16896
rect 14372 16832 14388 16896
rect 14452 16832 14468 16896
rect 14532 16832 14548 16896
rect 14612 16832 14618 16896
rect 14302 16831 14618 16832
rect 21662 16896 21978 16897
rect 21662 16832 21668 16896
rect 21732 16832 21748 16896
rect 21812 16832 21828 16896
rect 21892 16832 21908 16896
rect 21972 16832 21978 16896
rect 21662 16831 21978 16832
rect 29022 16896 29338 16897
rect 29022 16832 29028 16896
rect 29092 16832 29108 16896
rect 29172 16832 29188 16896
rect 29252 16832 29268 16896
rect 29332 16832 29338 16896
rect 29022 16831 29338 16832
rect 10961 16690 11027 16693
rect 15653 16690 15719 16693
rect 10961 16688 15719 16690
rect 10961 16632 10966 16688
rect 11022 16632 15658 16688
rect 15714 16632 15719 16688
rect 10961 16630 15719 16632
rect 10961 16627 11027 16630
rect 15653 16627 15719 16630
rect 10409 16554 10475 16557
rect 11094 16554 11100 16556
rect 10409 16552 11100 16554
rect 10409 16496 10414 16552
rect 10470 16496 11100 16552
rect 10409 16494 11100 16496
rect 10409 16491 10475 16494
rect 11094 16492 11100 16494
rect 11164 16492 11170 16556
rect 12525 16554 12591 16557
rect 16614 16554 16620 16556
rect 12525 16552 16620 16554
rect 12525 16496 12530 16552
rect 12586 16496 16620 16552
rect 12525 16494 16620 16496
rect 12525 16491 12591 16494
rect 16614 16492 16620 16494
rect 16684 16492 16690 16556
rect 6282 16352 6598 16353
rect 6282 16288 6288 16352
rect 6352 16288 6368 16352
rect 6432 16288 6448 16352
rect 6512 16288 6528 16352
rect 6592 16288 6598 16352
rect 6282 16287 6598 16288
rect 13642 16352 13958 16353
rect 13642 16288 13648 16352
rect 13712 16288 13728 16352
rect 13792 16288 13808 16352
rect 13872 16288 13888 16352
rect 13952 16288 13958 16352
rect 13642 16287 13958 16288
rect 21002 16352 21318 16353
rect 21002 16288 21008 16352
rect 21072 16288 21088 16352
rect 21152 16288 21168 16352
rect 21232 16288 21248 16352
rect 21312 16288 21318 16352
rect 21002 16287 21318 16288
rect 28362 16352 28678 16353
rect 28362 16288 28368 16352
rect 28432 16288 28448 16352
rect 28512 16288 28528 16352
rect 28592 16288 28608 16352
rect 28672 16288 28678 16352
rect 28362 16287 28678 16288
rect 14089 16146 14155 16149
rect 15469 16146 15535 16149
rect 14089 16144 15535 16146
rect 14089 16088 14094 16144
rect 14150 16088 15474 16144
rect 15530 16088 15535 16144
rect 14089 16086 15535 16088
rect 14089 16083 14155 16086
rect 15469 16083 15535 16086
rect 6942 15808 7258 15809
rect 0 15738 800 15768
rect 6942 15744 6948 15808
rect 7012 15744 7028 15808
rect 7092 15744 7108 15808
rect 7172 15744 7188 15808
rect 7252 15744 7258 15808
rect 6942 15743 7258 15744
rect 14302 15808 14618 15809
rect 14302 15744 14308 15808
rect 14372 15744 14388 15808
rect 14452 15744 14468 15808
rect 14532 15744 14548 15808
rect 14612 15744 14618 15808
rect 14302 15743 14618 15744
rect 21662 15808 21978 15809
rect 21662 15744 21668 15808
rect 21732 15744 21748 15808
rect 21812 15744 21828 15808
rect 21892 15744 21908 15808
rect 21972 15744 21978 15808
rect 21662 15743 21978 15744
rect 29022 15808 29338 15809
rect 29022 15744 29028 15808
rect 29092 15744 29108 15808
rect 29172 15744 29188 15808
rect 29252 15744 29268 15808
rect 29332 15744 29338 15808
rect 29022 15743 29338 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 33133 15738 33199 15741
rect 34168 15738 34968 15768
rect 33133 15736 34968 15738
rect 33133 15680 33138 15736
rect 33194 15680 34968 15736
rect 33133 15678 34968 15680
rect 33133 15675 33199 15678
rect 34168 15648 34968 15678
rect 6282 15264 6598 15265
rect 6282 15200 6288 15264
rect 6352 15200 6368 15264
rect 6432 15200 6448 15264
rect 6512 15200 6528 15264
rect 6592 15200 6598 15264
rect 6282 15199 6598 15200
rect 13642 15264 13958 15265
rect 13642 15200 13648 15264
rect 13712 15200 13728 15264
rect 13792 15200 13808 15264
rect 13872 15200 13888 15264
rect 13952 15200 13958 15264
rect 13642 15199 13958 15200
rect 21002 15264 21318 15265
rect 21002 15200 21008 15264
rect 21072 15200 21088 15264
rect 21152 15200 21168 15264
rect 21232 15200 21248 15264
rect 21312 15200 21318 15264
rect 21002 15199 21318 15200
rect 28362 15264 28678 15265
rect 28362 15200 28368 15264
rect 28432 15200 28448 15264
rect 28512 15200 28528 15264
rect 28592 15200 28608 15264
rect 28672 15200 28678 15264
rect 28362 15199 28678 15200
rect 15377 15196 15443 15197
rect 15326 15132 15332 15196
rect 15396 15194 15443 15196
rect 15396 15192 15488 15194
rect 15438 15136 15488 15192
rect 15396 15134 15488 15136
rect 15396 15132 15443 15134
rect 15377 15131 15443 15132
rect 11789 15058 11855 15061
rect 13353 15058 13419 15061
rect 11789 15056 13419 15058
rect 11789 15000 11794 15056
rect 11850 15000 13358 15056
rect 13414 15000 13419 15056
rect 11789 14998 13419 15000
rect 11789 14995 11855 14998
rect 13353 14995 13419 14998
rect 11513 14922 11579 14925
rect 14089 14922 14155 14925
rect 11513 14920 14155 14922
rect 11513 14864 11518 14920
rect 11574 14864 14094 14920
rect 14150 14864 14155 14920
rect 11513 14862 14155 14864
rect 11513 14859 11579 14862
rect 14089 14859 14155 14862
rect 12801 14786 12867 14789
rect 13353 14786 13419 14789
rect 12801 14784 13419 14786
rect 12801 14728 12806 14784
rect 12862 14728 13358 14784
rect 13414 14728 13419 14784
rect 12801 14726 13419 14728
rect 12801 14723 12867 14726
rect 13353 14723 13419 14726
rect 6942 14720 7258 14721
rect 6942 14656 6948 14720
rect 7012 14656 7028 14720
rect 7092 14656 7108 14720
rect 7172 14656 7188 14720
rect 7252 14656 7258 14720
rect 6942 14655 7258 14656
rect 14302 14720 14618 14721
rect 14302 14656 14308 14720
rect 14372 14656 14388 14720
rect 14452 14656 14468 14720
rect 14532 14656 14548 14720
rect 14612 14656 14618 14720
rect 14302 14655 14618 14656
rect 21662 14720 21978 14721
rect 21662 14656 21668 14720
rect 21732 14656 21748 14720
rect 21812 14656 21828 14720
rect 21892 14656 21908 14720
rect 21972 14656 21978 14720
rect 21662 14655 21978 14656
rect 29022 14720 29338 14721
rect 29022 14656 29028 14720
rect 29092 14656 29108 14720
rect 29172 14656 29188 14720
rect 29252 14656 29268 14720
rect 29332 14656 29338 14720
rect 29022 14655 29338 14656
rect 0 14378 800 14408
rect 1301 14378 1367 14381
rect 0 14376 1367 14378
rect 0 14320 1306 14376
rect 1362 14320 1367 14376
rect 0 14318 1367 14320
rect 0 14288 800 14318
rect 1301 14315 1367 14318
rect 7741 14378 7807 14381
rect 16665 14378 16731 14381
rect 7741 14376 16731 14378
rect 7741 14320 7746 14376
rect 7802 14320 16670 14376
rect 16726 14320 16731 14376
rect 7741 14318 16731 14320
rect 7741 14315 7807 14318
rect 16665 14315 16731 14318
rect 33133 14378 33199 14381
rect 34168 14378 34968 14408
rect 33133 14376 34968 14378
rect 33133 14320 33138 14376
rect 33194 14320 34968 14376
rect 33133 14318 34968 14320
rect 33133 14315 33199 14318
rect 34168 14288 34968 14318
rect 12249 14244 12315 14245
rect 12198 14180 12204 14244
rect 12268 14242 12315 14244
rect 20069 14242 20135 14245
rect 12268 14240 13554 14242
rect 12310 14184 13554 14240
rect 12268 14182 13554 14184
rect 12268 14180 12315 14182
rect 12249 14179 12315 14180
rect 6282 14176 6598 14177
rect 6282 14112 6288 14176
rect 6352 14112 6368 14176
rect 6432 14112 6448 14176
rect 6512 14112 6528 14176
rect 6592 14112 6598 14176
rect 6282 14111 6598 14112
rect 13494 13970 13554 14182
rect 19290 14240 20135 14242
rect 19290 14184 20074 14240
rect 20130 14184 20135 14240
rect 19290 14182 20135 14184
rect 13642 14176 13958 14177
rect 13642 14112 13648 14176
rect 13712 14112 13728 14176
rect 13792 14112 13808 14176
rect 13872 14112 13888 14176
rect 13952 14112 13958 14176
rect 13642 14111 13958 14112
rect 19290 13970 19350 14182
rect 20069 14179 20135 14182
rect 21002 14176 21318 14177
rect 21002 14112 21008 14176
rect 21072 14112 21088 14176
rect 21152 14112 21168 14176
rect 21232 14112 21248 14176
rect 21312 14112 21318 14176
rect 21002 14111 21318 14112
rect 28362 14176 28678 14177
rect 28362 14112 28368 14176
rect 28432 14112 28448 14176
rect 28512 14112 28528 14176
rect 28592 14112 28608 14176
rect 28672 14112 28678 14176
rect 28362 14111 28678 14112
rect 13494 13910 19350 13970
rect 28993 13834 29059 13837
rect 29545 13834 29611 13837
rect 31017 13834 31083 13837
rect 28993 13832 31083 13834
rect 28993 13776 28998 13832
rect 29054 13776 29550 13832
rect 29606 13776 31022 13832
rect 31078 13776 31083 13832
rect 28993 13774 31083 13776
rect 28993 13771 29059 13774
rect 29545 13771 29611 13774
rect 31017 13771 31083 13774
rect 16430 13636 16436 13700
rect 16500 13698 16506 13700
rect 17125 13698 17191 13701
rect 16500 13696 17191 13698
rect 16500 13640 17130 13696
rect 17186 13640 17191 13696
rect 16500 13638 17191 13640
rect 16500 13636 16506 13638
rect 17125 13635 17191 13638
rect 6942 13632 7258 13633
rect 6942 13568 6948 13632
rect 7012 13568 7028 13632
rect 7092 13568 7108 13632
rect 7172 13568 7188 13632
rect 7252 13568 7258 13632
rect 6942 13567 7258 13568
rect 14302 13632 14618 13633
rect 14302 13568 14308 13632
rect 14372 13568 14388 13632
rect 14452 13568 14468 13632
rect 14532 13568 14548 13632
rect 14612 13568 14618 13632
rect 14302 13567 14618 13568
rect 21662 13632 21978 13633
rect 21662 13568 21668 13632
rect 21732 13568 21748 13632
rect 21812 13568 21828 13632
rect 21892 13568 21908 13632
rect 21972 13568 21978 13632
rect 21662 13567 21978 13568
rect 29022 13632 29338 13633
rect 29022 13568 29028 13632
rect 29092 13568 29108 13632
rect 29172 13568 29188 13632
rect 29252 13568 29268 13632
rect 29332 13568 29338 13632
rect 29022 13567 29338 13568
rect 30557 13426 30623 13429
rect 31753 13426 31819 13429
rect 30557 13424 31819 13426
rect 30557 13368 30562 13424
rect 30618 13368 31758 13424
rect 31814 13368 31819 13424
rect 30557 13366 31819 13368
rect 30557 13363 30623 13366
rect 31753 13363 31819 13366
rect 28993 13290 29059 13293
rect 29729 13290 29795 13293
rect 28993 13288 29795 13290
rect 28993 13232 28998 13288
rect 29054 13232 29734 13288
rect 29790 13232 29795 13288
rect 28993 13230 29795 13232
rect 28993 13227 29059 13230
rect 29729 13227 29795 13230
rect 6282 13088 6598 13089
rect 0 13018 800 13048
rect 6282 13024 6288 13088
rect 6352 13024 6368 13088
rect 6432 13024 6448 13088
rect 6512 13024 6528 13088
rect 6592 13024 6598 13088
rect 6282 13023 6598 13024
rect 13642 13088 13958 13089
rect 13642 13024 13648 13088
rect 13712 13024 13728 13088
rect 13792 13024 13808 13088
rect 13872 13024 13888 13088
rect 13952 13024 13958 13088
rect 13642 13023 13958 13024
rect 21002 13088 21318 13089
rect 21002 13024 21008 13088
rect 21072 13024 21088 13088
rect 21152 13024 21168 13088
rect 21232 13024 21248 13088
rect 21312 13024 21318 13088
rect 21002 13023 21318 13024
rect 28362 13088 28678 13089
rect 28362 13024 28368 13088
rect 28432 13024 28448 13088
rect 28512 13024 28528 13088
rect 28592 13024 28608 13088
rect 28672 13024 28678 13088
rect 28362 13023 28678 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 26141 12882 26207 12885
rect 28901 12882 28967 12885
rect 26141 12880 28967 12882
rect 26141 12824 26146 12880
rect 26202 12824 28906 12880
rect 28962 12824 28967 12880
rect 26141 12822 28967 12824
rect 26141 12819 26207 12822
rect 28901 12819 28967 12822
rect 6942 12544 7258 12545
rect 6942 12480 6948 12544
rect 7012 12480 7028 12544
rect 7092 12480 7108 12544
rect 7172 12480 7188 12544
rect 7252 12480 7258 12544
rect 6942 12479 7258 12480
rect 14302 12544 14618 12545
rect 14302 12480 14308 12544
rect 14372 12480 14388 12544
rect 14452 12480 14468 12544
rect 14532 12480 14548 12544
rect 14612 12480 14618 12544
rect 14302 12479 14618 12480
rect 21662 12544 21978 12545
rect 21662 12480 21668 12544
rect 21732 12480 21748 12544
rect 21812 12480 21828 12544
rect 21892 12480 21908 12544
rect 21972 12480 21978 12544
rect 21662 12479 21978 12480
rect 29022 12544 29338 12545
rect 29022 12480 29028 12544
rect 29092 12480 29108 12544
rect 29172 12480 29188 12544
rect 29252 12480 29268 12544
rect 29332 12480 29338 12544
rect 29022 12479 29338 12480
rect 8109 12474 8175 12477
rect 11053 12474 11119 12477
rect 8109 12472 11119 12474
rect 8109 12416 8114 12472
rect 8170 12416 11058 12472
rect 11114 12416 11119 12472
rect 8109 12414 11119 12416
rect 8109 12411 8175 12414
rect 11053 12411 11119 12414
rect 6913 12338 6979 12341
rect 11145 12338 11211 12341
rect 6913 12336 11211 12338
rect 6913 12280 6918 12336
rect 6974 12280 11150 12336
rect 11206 12280 11211 12336
rect 6913 12278 11211 12280
rect 6913 12275 6979 12278
rect 11145 12275 11211 12278
rect 33133 12338 33199 12341
rect 34168 12338 34968 12368
rect 33133 12336 34968 12338
rect 33133 12280 33138 12336
rect 33194 12280 34968 12336
rect 33133 12278 34968 12280
rect 33133 12275 33199 12278
rect 34168 12248 34968 12278
rect 24577 12202 24643 12205
rect 26601 12202 26667 12205
rect 24577 12200 26667 12202
rect 24577 12144 24582 12200
rect 24638 12144 26606 12200
rect 26662 12144 26667 12200
rect 24577 12142 26667 12144
rect 24577 12139 24643 12142
rect 26601 12139 26667 12142
rect 6282 12000 6598 12001
rect 6282 11936 6288 12000
rect 6352 11936 6368 12000
rect 6432 11936 6448 12000
rect 6512 11936 6528 12000
rect 6592 11936 6598 12000
rect 6282 11935 6598 11936
rect 13642 12000 13958 12001
rect 13642 11936 13648 12000
rect 13712 11936 13728 12000
rect 13792 11936 13808 12000
rect 13872 11936 13888 12000
rect 13952 11936 13958 12000
rect 13642 11935 13958 11936
rect 21002 12000 21318 12001
rect 21002 11936 21008 12000
rect 21072 11936 21088 12000
rect 21152 11936 21168 12000
rect 21232 11936 21248 12000
rect 21312 11936 21318 12000
rect 21002 11935 21318 11936
rect 28362 12000 28678 12001
rect 28362 11936 28368 12000
rect 28432 11936 28448 12000
rect 28512 11936 28528 12000
rect 28592 11936 28608 12000
rect 28672 11936 28678 12000
rect 28362 11935 28678 11936
rect 24485 11932 24551 11933
rect 24485 11930 24532 11932
rect 24440 11928 24532 11930
rect 24440 11872 24490 11928
rect 24440 11870 24532 11872
rect 24485 11868 24532 11870
rect 24596 11868 24602 11932
rect 24485 11867 24551 11868
rect 6942 11456 7258 11457
rect 6942 11392 6948 11456
rect 7012 11392 7028 11456
rect 7092 11392 7108 11456
rect 7172 11392 7188 11456
rect 7252 11392 7258 11456
rect 6942 11391 7258 11392
rect 14302 11456 14618 11457
rect 14302 11392 14308 11456
rect 14372 11392 14388 11456
rect 14452 11392 14468 11456
rect 14532 11392 14548 11456
rect 14612 11392 14618 11456
rect 14302 11391 14618 11392
rect 21662 11456 21978 11457
rect 21662 11392 21668 11456
rect 21732 11392 21748 11456
rect 21812 11392 21828 11456
rect 21892 11392 21908 11456
rect 21972 11392 21978 11456
rect 21662 11391 21978 11392
rect 29022 11456 29338 11457
rect 29022 11392 29028 11456
rect 29092 11392 29108 11456
rect 29172 11392 29188 11456
rect 29252 11392 29268 11456
rect 29332 11392 29338 11456
rect 29022 11391 29338 11392
rect 13997 11250 14063 11253
rect 14774 11250 14780 11252
rect 13997 11248 14780 11250
rect 13997 11192 14002 11248
rect 14058 11192 14780 11248
rect 13997 11190 14780 11192
rect 13997 11187 14063 11190
rect 14774 11188 14780 11190
rect 14844 11188 14850 11252
rect 0 10978 800 11008
rect 3233 10978 3299 10981
rect 0 10976 3299 10978
rect 0 10920 3238 10976
rect 3294 10920 3299 10976
rect 0 10918 3299 10920
rect 0 10888 800 10918
rect 3233 10915 3299 10918
rect 31385 10978 31451 10981
rect 34168 10978 34968 11008
rect 31385 10976 34968 10978
rect 31385 10920 31390 10976
rect 31446 10920 34968 10976
rect 31385 10918 34968 10920
rect 31385 10915 31451 10918
rect 6282 10912 6598 10913
rect 6282 10848 6288 10912
rect 6352 10848 6368 10912
rect 6432 10848 6448 10912
rect 6512 10848 6528 10912
rect 6592 10848 6598 10912
rect 6282 10847 6598 10848
rect 13642 10912 13958 10913
rect 13642 10848 13648 10912
rect 13712 10848 13728 10912
rect 13792 10848 13808 10912
rect 13872 10848 13888 10912
rect 13952 10848 13958 10912
rect 13642 10847 13958 10848
rect 21002 10912 21318 10913
rect 21002 10848 21008 10912
rect 21072 10848 21088 10912
rect 21152 10848 21168 10912
rect 21232 10848 21248 10912
rect 21312 10848 21318 10912
rect 21002 10847 21318 10848
rect 28362 10912 28678 10913
rect 28362 10848 28368 10912
rect 28432 10848 28448 10912
rect 28512 10848 28528 10912
rect 28592 10848 28608 10912
rect 28672 10848 28678 10912
rect 34168 10888 34968 10918
rect 28362 10847 28678 10848
rect 6942 10368 7258 10369
rect 6942 10304 6948 10368
rect 7012 10304 7028 10368
rect 7092 10304 7108 10368
rect 7172 10304 7188 10368
rect 7252 10304 7258 10368
rect 6942 10303 7258 10304
rect 14302 10368 14618 10369
rect 14302 10304 14308 10368
rect 14372 10304 14388 10368
rect 14452 10304 14468 10368
rect 14532 10304 14548 10368
rect 14612 10304 14618 10368
rect 14302 10303 14618 10304
rect 21662 10368 21978 10369
rect 21662 10304 21668 10368
rect 21732 10304 21748 10368
rect 21812 10304 21828 10368
rect 21892 10304 21908 10368
rect 21972 10304 21978 10368
rect 21662 10303 21978 10304
rect 29022 10368 29338 10369
rect 29022 10304 29028 10368
rect 29092 10304 29108 10368
rect 29172 10304 29188 10368
rect 29252 10304 29268 10368
rect 29332 10304 29338 10368
rect 29022 10303 29338 10304
rect 6282 9824 6598 9825
rect 6282 9760 6288 9824
rect 6352 9760 6368 9824
rect 6432 9760 6448 9824
rect 6512 9760 6528 9824
rect 6592 9760 6598 9824
rect 6282 9759 6598 9760
rect 13642 9824 13958 9825
rect 13642 9760 13648 9824
rect 13712 9760 13728 9824
rect 13792 9760 13808 9824
rect 13872 9760 13888 9824
rect 13952 9760 13958 9824
rect 13642 9759 13958 9760
rect 21002 9824 21318 9825
rect 21002 9760 21008 9824
rect 21072 9760 21088 9824
rect 21152 9760 21168 9824
rect 21232 9760 21248 9824
rect 21312 9760 21318 9824
rect 21002 9759 21318 9760
rect 28362 9824 28678 9825
rect 28362 9760 28368 9824
rect 28432 9760 28448 9824
rect 28512 9760 28528 9824
rect 28592 9760 28608 9824
rect 28672 9760 28678 9824
rect 28362 9759 28678 9760
rect 0 9618 800 9648
rect 3049 9618 3115 9621
rect 0 9616 3115 9618
rect 0 9560 3054 9616
rect 3110 9560 3115 9616
rect 0 9558 3115 9560
rect 0 9528 800 9558
rect 3049 9555 3115 9558
rect 20253 9618 20319 9621
rect 23565 9618 23631 9621
rect 20253 9616 23631 9618
rect 20253 9560 20258 9616
rect 20314 9560 23570 9616
rect 23626 9560 23631 9616
rect 20253 9558 23631 9560
rect 20253 9555 20319 9558
rect 23565 9555 23631 9558
rect 33133 9618 33199 9621
rect 34168 9618 34968 9648
rect 33133 9616 34968 9618
rect 33133 9560 33138 9616
rect 33194 9560 34968 9616
rect 33133 9558 34968 9560
rect 33133 9555 33199 9558
rect 34168 9528 34968 9558
rect 21817 9482 21883 9485
rect 22461 9482 22527 9485
rect 23657 9482 23723 9485
rect 21817 9480 23723 9482
rect 21817 9424 21822 9480
rect 21878 9424 22466 9480
rect 22522 9424 23662 9480
rect 23718 9424 23723 9480
rect 21817 9422 23723 9424
rect 21817 9419 21883 9422
rect 22461 9419 22527 9422
rect 23657 9419 23723 9422
rect 26233 9482 26299 9485
rect 27521 9482 27587 9485
rect 28625 9482 28691 9485
rect 29177 9482 29243 9485
rect 26233 9480 29243 9482
rect 26233 9424 26238 9480
rect 26294 9424 27526 9480
rect 27582 9424 28630 9480
rect 28686 9424 29182 9480
rect 29238 9424 29243 9480
rect 26233 9422 29243 9424
rect 26233 9419 26299 9422
rect 27521 9419 27587 9422
rect 28625 9419 28691 9422
rect 29177 9419 29243 9422
rect 6942 9280 7258 9281
rect 6942 9216 6948 9280
rect 7012 9216 7028 9280
rect 7092 9216 7108 9280
rect 7172 9216 7188 9280
rect 7252 9216 7258 9280
rect 6942 9215 7258 9216
rect 14302 9280 14618 9281
rect 14302 9216 14308 9280
rect 14372 9216 14388 9280
rect 14452 9216 14468 9280
rect 14532 9216 14548 9280
rect 14612 9216 14618 9280
rect 14302 9215 14618 9216
rect 21662 9280 21978 9281
rect 21662 9216 21668 9280
rect 21732 9216 21748 9280
rect 21812 9216 21828 9280
rect 21892 9216 21908 9280
rect 21972 9216 21978 9280
rect 21662 9215 21978 9216
rect 29022 9280 29338 9281
rect 29022 9216 29028 9280
rect 29092 9216 29108 9280
rect 29172 9216 29188 9280
rect 29252 9216 29268 9280
rect 29332 9216 29338 9280
rect 29022 9215 29338 9216
rect 10869 9074 10935 9077
rect 31661 9074 31727 9077
rect 10869 9072 31727 9074
rect 10869 9016 10874 9072
rect 10930 9016 31666 9072
rect 31722 9016 31727 9072
rect 10869 9014 31727 9016
rect 10869 9011 10935 9014
rect 31661 9011 31727 9014
rect 6282 8736 6598 8737
rect 6282 8672 6288 8736
rect 6352 8672 6368 8736
rect 6432 8672 6448 8736
rect 6512 8672 6528 8736
rect 6592 8672 6598 8736
rect 6282 8671 6598 8672
rect 13642 8736 13958 8737
rect 13642 8672 13648 8736
rect 13712 8672 13728 8736
rect 13792 8672 13808 8736
rect 13872 8672 13888 8736
rect 13952 8672 13958 8736
rect 13642 8671 13958 8672
rect 21002 8736 21318 8737
rect 21002 8672 21008 8736
rect 21072 8672 21088 8736
rect 21152 8672 21168 8736
rect 21232 8672 21248 8736
rect 21312 8672 21318 8736
rect 21002 8671 21318 8672
rect 28362 8736 28678 8737
rect 28362 8672 28368 8736
rect 28432 8672 28448 8736
rect 28512 8672 28528 8736
rect 28592 8672 28608 8736
rect 28672 8672 28678 8736
rect 28362 8671 28678 8672
rect 25129 8530 25195 8533
rect 28441 8530 28507 8533
rect 25129 8528 28507 8530
rect 25129 8472 25134 8528
rect 25190 8472 28446 8528
rect 28502 8472 28507 8528
rect 25129 8470 28507 8472
rect 25129 8467 25195 8470
rect 28441 8467 28507 8470
rect 21725 8394 21791 8397
rect 23381 8394 23447 8397
rect 21725 8392 23447 8394
rect 21725 8336 21730 8392
rect 21786 8336 23386 8392
rect 23442 8336 23447 8392
rect 21725 8334 23447 8336
rect 21725 8331 21791 8334
rect 23381 8331 23447 8334
rect 13118 8196 13124 8260
rect 13188 8258 13194 8260
rect 13261 8258 13327 8261
rect 13188 8256 13327 8258
rect 13188 8200 13266 8256
rect 13322 8200 13327 8256
rect 13188 8198 13327 8200
rect 13188 8196 13194 8198
rect 13261 8195 13327 8198
rect 6942 8192 7258 8193
rect 6942 8128 6948 8192
rect 7012 8128 7028 8192
rect 7092 8128 7108 8192
rect 7172 8128 7188 8192
rect 7252 8128 7258 8192
rect 6942 8127 7258 8128
rect 14302 8192 14618 8193
rect 14302 8128 14308 8192
rect 14372 8128 14388 8192
rect 14452 8128 14468 8192
rect 14532 8128 14548 8192
rect 14612 8128 14618 8192
rect 14302 8127 14618 8128
rect 21662 8192 21978 8193
rect 21662 8128 21668 8192
rect 21732 8128 21748 8192
rect 21812 8128 21828 8192
rect 21892 8128 21908 8192
rect 21972 8128 21978 8192
rect 21662 8127 21978 8128
rect 29022 8192 29338 8193
rect 29022 8128 29028 8192
rect 29092 8128 29108 8192
rect 29172 8128 29188 8192
rect 29252 8128 29268 8192
rect 29332 8128 29338 8192
rect 29022 8127 29338 8128
rect 25865 7986 25931 7989
rect 28165 7986 28231 7989
rect 25865 7984 28231 7986
rect 25865 7928 25870 7984
rect 25926 7928 28170 7984
rect 28226 7928 28231 7984
rect 25865 7926 28231 7928
rect 25865 7923 25931 7926
rect 28165 7923 28231 7926
rect 29453 7850 29519 7853
rect 31569 7850 31635 7853
rect 29453 7848 31635 7850
rect 29453 7792 29458 7848
rect 29514 7792 31574 7848
rect 31630 7792 31635 7848
rect 29453 7790 31635 7792
rect 29453 7787 29519 7790
rect 31569 7787 31635 7790
rect 6282 7648 6598 7649
rect 0 7578 800 7608
rect 6282 7584 6288 7648
rect 6352 7584 6368 7648
rect 6432 7584 6448 7648
rect 6512 7584 6528 7648
rect 6592 7584 6598 7648
rect 6282 7583 6598 7584
rect 13642 7648 13958 7649
rect 13642 7584 13648 7648
rect 13712 7584 13728 7648
rect 13792 7584 13808 7648
rect 13872 7584 13888 7648
rect 13952 7584 13958 7648
rect 13642 7583 13958 7584
rect 21002 7648 21318 7649
rect 21002 7584 21008 7648
rect 21072 7584 21088 7648
rect 21152 7584 21168 7648
rect 21232 7584 21248 7648
rect 21312 7584 21318 7648
rect 21002 7583 21318 7584
rect 28362 7648 28678 7649
rect 28362 7584 28368 7648
rect 28432 7584 28448 7648
rect 28512 7584 28528 7648
rect 28592 7584 28608 7648
rect 28672 7584 28678 7648
rect 28362 7583 28678 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 33133 7578 33199 7581
rect 34168 7578 34968 7608
rect 33133 7576 34968 7578
rect 33133 7520 33138 7576
rect 33194 7520 34968 7576
rect 33133 7518 34968 7520
rect 33133 7515 33199 7518
rect 34168 7488 34968 7518
rect 6942 7104 7258 7105
rect 6942 7040 6948 7104
rect 7012 7040 7028 7104
rect 7092 7040 7108 7104
rect 7172 7040 7188 7104
rect 7252 7040 7258 7104
rect 6942 7039 7258 7040
rect 14302 7104 14618 7105
rect 14302 7040 14308 7104
rect 14372 7040 14388 7104
rect 14452 7040 14468 7104
rect 14532 7040 14548 7104
rect 14612 7040 14618 7104
rect 14302 7039 14618 7040
rect 21662 7104 21978 7105
rect 21662 7040 21668 7104
rect 21732 7040 21748 7104
rect 21812 7040 21828 7104
rect 21892 7040 21908 7104
rect 21972 7040 21978 7104
rect 21662 7039 21978 7040
rect 29022 7104 29338 7105
rect 29022 7040 29028 7104
rect 29092 7040 29108 7104
rect 29172 7040 29188 7104
rect 29252 7040 29268 7104
rect 29332 7040 29338 7104
rect 29022 7039 29338 7040
rect 12985 6898 13051 6901
rect 13302 6898 13308 6900
rect 12985 6896 13308 6898
rect 12985 6840 12990 6896
rect 13046 6840 13308 6896
rect 12985 6838 13308 6840
rect 12985 6835 13051 6838
rect 13302 6836 13308 6838
rect 13372 6836 13378 6900
rect 17718 6836 17724 6900
rect 17788 6898 17794 6900
rect 18597 6898 18663 6901
rect 17788 6896 18663 6898
rect 17788 6840 18602 6896
rect 18658 6840 18663 6896
rect 17788 6838 18663 6840
rect 17788 6836 17794 6838
rect 18597 6835 18663 6838
rect 6282 6560 6598 6561
rect 6282 6496 6288 6560
rect 6352 6496 6368 6560
rect 6432 6496 6448 6560
rect 6512 6496 6528 6560
rect 6592 6496 6598 6560
rect 6282 6495 6598 6496
rect 13642 6560 13958 6561
rect 13642 6496 13648 6560
rect 13712 6496 13728 6560
rect 13792 6496 13808 6560
rect 13872 6496 13888 6560
rect 13952 6496 13958 6560
rect 13642 6495 13958 6496
rect 21002 6560 21318 6561
rect 21002 6496 21008 6560
rect 21072 6496 21088 6560
rect 21152 6496 21168 6560
rect 21232 6496 21248 6560
rect 21312 6496 21318 6560
rect 21002 6495 21318 6496
rect 28362 6560 28678 6561
rect 28362 6496 28368 6560
rect 28432 6496 28448 6560
rect 28512 6496 28528 6560
rect 28592 6496 28608 6560
rect 28672 6496 28678 6560
rect 28362 6495 28678 6496
rect 15285 6354 15351 6357
rect 21357 6354 21423 6357
rect 15285 6352 21423 6354
rect 15285 6296 15290 6352
rect 15346 6296 21362 6352
rect 21418 6296 21423 6352
rect 15285 6294 21423 6296
rect 15285 6291 15351 6294
rect 21357 6291 21423 6294
rect 0 6218 800 6248
rect 1301 6218 1367 6221
rect 0 6216 1367 6218
rect 0 6160 1306 6216
rect 1362 6160 1367 6216
rect 0 6158 1367 6160
rect 0 6128 800 6158
rect 1301 6155 1367 6158
rect 33133 6218 33199 6221
rect 34168 6218 34968 6248
rect 33133 6216 34968 6218
rect 33133 6160 33138 6216
rect 33194 6160 34968 6216
rect 33133 6158 34968 6160
rect 33133 6155 33199 6158
rect 34168 6128 34968 6158
rect 6942 6016 7258 6017
rect 6942 5952 6948 6016
rect 7012 5952 7028 6016
rect 7092 5952 7108 6016
rect 7172 5952 7188 6016
rect 7252 5952 7258 6016
rect 6942 5951 7258 5952
rect 14302 6016 14618 6017
rect 14302 5952 14308 6016
rect 14372 5952 14388 6016
rect 14452 5952 14468 6016
rect 14532 5952 14548 6016
rect 14612 5952 14618 6016
rect 14302 5951 14618 5952
rect 21662 6016 21978 6017
rect 21662 5952 21668 6016
rect 21732 5952 21748 6016
rect 21812 5952 21828 6016
rect 21892 5952 21908 6016
rect 21972 5952 21978 6016
rect 21662 5951 21978 5952
rect 29022 6016 29338 6017
rect 29022 5952 29028 6016
rect 29092 5952 29108 6016
rect 29172 5952 29188 6016
rect 29252 5952 29268 6016
rect 29332 5952 29338 6016
rect 29022 5951 29338 5952
rect 22737 5674 22803 5677
rect 29729 5674 29795 5677
rect 22737 5672 29795 5674
rect 22737 5616 22742 5672
rect 22798 5616 29734 5672
rect 29790 5616 29795 5672
rect 22737 5614 29795 5616
rect 22737 5611 22803 5614
rect 29729 5611 29795 5614
rect 12985 5540 13051 5541
rect 12934 5476 12940 5540
rect 13004 5538 13051 5540
rect 13004 5536 13096 5538
rect 13046 5480 13096 5536
rect 13004 5478 13096 5480
rect 13004 5476 13051 5478
rect 12985 5475 13051 5476
rect 6282 5472 6598 5473
rect 6282 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6598 5472
rect 6282 5407 6598 5408
rect 13642 5472 13958 5473
rect 13642 5408 13648 5472
rect 13712 5408 13728 5472
rect 13792 5408 13808 5472
rect 13872 5408 13888 5472
rect 13952 5408 13958 5472
rect 13642 5407 13958 5408
rect 21002 5472 21318 5473
rect 21002 5408 21008 5472
rect 21072 5408 21088 5472
rect 21152 5408 21168 5472
rect 21232 5408 21248 5472
rect 21312 5408 21318 5472
rect 21002 5407 21318 5408
rect 28362 5472 28678 5473
rect 28362 5408 28368 5472
rect 28432 5408 28448 5472
rect 28512 5408 28528 5472
rect 28592 5408 28608 5472
rect 28672 5408 28678 5472
rect 28362 5407 28678 5408
rect 15745 5266 15811 5269
rect 18045 5266 18111 5269
rect 15745 5264 18111 5266
rect 15745 5208 15750 5264
rect 15806 5208 18050 5264
rect 18106 5208 18111 5264
rect 15745 5206 18111 5208
rect 15745 5203 15811 5206
rect 18045 5203 18111 5206
rect 19241 5266 19307 5269
rect 31661 5266 31727 5269
rect 19241 5264 31727 5266
rect 19241 5208 19246 5264
rect 19302 5208 31666 5264
rect 31722 5208 31727 5264
rect 19241 5206 31727 5208
rect 19241 5203 19307 5206
rect 31661 5203 31727 5206
rect 18597 5130 18663 5133
rect 20713 5130 20779 5133
rect 18597 5128 20779 5130
rect 18597 5072 18602 5128
rect 18658 5072 20718 5128
rect 20774 5072 20779 5128
rect 18597 5070 20779 5072
rect 18597 5067 18663 5070
rect 20713 5067 20779 5070
rect 6942 4928 7258 4929
rect 0 4858 800 4888
rect 6942 4864 6948 4928
rect 7012 4864 7028 4928
rect 7092 4864 7108 4928
rect 7172 4864 7188 4928
rect 7252 4864 7258 4928
rect 6942 4863 7258 4864
rect 14302 4928 14618 4929
rect 14302 4864 14308 4928
rect 14372 4864 14388 4928
rect 14452 4864 14468 4928
rect 14532 4864 14548 4928
rect 14612 4864 14618 4928
rect 14302 4863 14618 4864
rect 21662 4928 21978 4929
rect 21662 4864 21668 4928
rect 21732 4864 21748 4928
rect 21812 4864 21828 4928
rect 21892 4864 21908 4928
rect 21972 4864 21978 4928
rect 21662 4863 21978 4864
rect 29022 4928 29338 4929
rect 29022 4864 29028 4928
rect 29092 4864 29108 4928
rect 29172 4864 29188 4928
rect 29252 4864 29268 4928
rect 29332 4864 29338 4928
rect 29022 4863 29338 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 6282 4384 6598 4385
rect 6282 4320 6288 4384
rect 6352 4320 6368 4384
rect 6432 4320 6448 4384
rect 6512 4320 6528 4384
rect 6592 4320 6598 4384
rect 6282 4319 6598 4320
rect 13642 4384 13958 4385
rect 13642 4320 13648 4384
rect 13712 4320 13728 4384
rect 13792 4320 13808 4384
rect 13872 4320 13888 4384
rect 13952 4320 13958 4384
rect 13642 4319 13958 4320
rect 21002 4384 21318 4385
rect 21002 4320 21008 4384
rect 21072 4320 21088 4384
rect 21152 4320 21168 4384
rect 21232 4320 21248 4384
rect 21312 4320 21318 4384
rect 21002 4319 21318 4320
rect 28362 4384 28678 4385
rect 28362 4320 28368 4384
rect 28432 4320 28448 4384
rect 28512 4320 28528 4384
rect 28592 4320 28608 4384
rect 28672 4320 28678 4384
rect 28362 4319 28678 4320
rect 33041 4178 33107 4181
rect 34168 4178 34968 4208
rect 33041 4176 34968 4178
rect 33041 4120 33046 4176
rect 33102 4120 34968 4176
rect 33041 4118 34968 4120
rect 33041 4115 33107 4118
rect 34168 4088 34968 4118
rect 6942 3840 7258 3841
rect 6942 3776 6948 3840
rect 7012 3776 7028 3840
rect 7092 3776 7108 3840
rect 7172 3776 7188 3840
rect 7252 3776 7258 3840
rect 6942 3775 7258 3776
rect 14302 3840 14618 3841
rect 14302 3776 14308 3840
rect 14372 3776 14388 3840
rect 14452 3776 14468 3840
rect 14532 3776 14548 3840
rect 14612 3776 14618 3840
rect 14302 3775 14618 3776
rect 21662 3840 21978 3841
rect 21662 3776 21668 3840
rect 21732 3776 21748 3840
rect 21812 3776 21828 3840
rect 21892 3776 21908 3840
rect 21972 3776 21978 3840
rect 21662 3775 21978 3776
rect 29022 3840 29338 3841
rect 29022 3776 29028 3840
rect 29092 3776 29108 3840
rect 29172 3776 29188 3840
rect 29252 3776 29268 3840
rect 29332 3776 29338 3840
rect 29022 3775 29338 3776
rect 6282 3296 6598 3297
rect 6282 3232 6288 3296
rect 6352 3232 6368 3296
rect 6432 3232 6448 3296
rect 6512 3232 6528 3296
rect 6592 3232 6598 3296
rect 6282 3231 6598 3232
rect 13642 3296 13958 3297
rect 13642 3232 13648 3296
rect 13712 3232 13728 3296
rect 13792 3232 13808 3296
rect 13872 3232 13888 3296
rect 13952 3232 13958 3296
rect 13642 3231 13958 3232
rect 21002 3296 21318 3297
rect 21002 3232 21008 3296
rect 21072 3232 21088 3296
rect 21152 3232 21168 3296
rect 21232 3232 21248 3296
rect 21312 3232 21318 3296
rect 21002 3231 21318 3232
rect 28362 3296 28678 3297
rect 28362 3232 28368 3296
rect 28432 3232 28448 3296
rect 28512 3232 28528 3296
rect 28592 3232 28608 3296
rect 28672 3232 28678 3296
rect 28362 3231 28678 3232
rect 0 2818 800 2848
rect 3601 2818 3667 2821
rect 0 2816 3667 2818
rect 0 2760 3606 2816
rect 3662 2760 3667 2816
rect 0 2758 3667 2760
rect 0 2728 800 2758
rect 3601 2755 3667 2758
rect 33133 2818 33199 2821
rect 34168 2818 34968 2848
rect 33133 2816 34968 2818
rect 33133 2760 33138 2816
rect 33194 2760 34968 2816
rect 33133 2758 34968 2760
rect 33133 2755 33199 2758
rect 6942 2752 7258 2753
rect 6942 2688 6948 2752
rect 7012 2688 7028 2752
rect 7092 2688 7108 2752
rect 7172 2688 7188 2752
rect 7252 2688 7258 2752
rect 6942 2687 7258 2688
rect 14302 2752 14618 2753
rect 14302 2688 14308 2752
rect 14372 2688 14388 2752
rect 14452 2688 14468 2752
rect 14532 2688 14548 2752
rect 14612 2688 14618 2752
rect 14302 2687 14618 2688
rect 21662 2752 21978 2753
rect 21662 2688 21668 2752
rect 21732 2688 21748 2752
rect 21812 2688 21828 2752
rect 21892 2688 21908 2752
rect 21972 2688 21978 2752
rect 21662 2687 21978 2688
rect 29022 2752 29338 2753
rect 29022 2688 29028 2752
rect 29092 2688 29108 2752
rect 29172 2688 29188 2752
rect 29252 2688 29268 2752
rect 29332 2688 29338 2752
rect 34168 2728 34968 2758
rect 29022 2687 29338 2688
rect 0 1458 800 1488
rect 3049 1458 3115 1461
rect 0 1456 3115 1458
rect 0 1400 3054 1456
rect 3110 1400 3115 1456
rect 0 1398 3115 1400
rect 0 1368 800 1398
rect 3049 1395 3115 1398
rect 31661 1458 31727 1461
rect 34168 1458 34968 1488
rect 31661 1456 34968 1458
rect 31661 1400 31666 1456
rect 31722 1400 34968 1456
rect 31661 1398 34968 1400
rect 31661 1395 31727 1398
rect 34168 1368 34968 1398
<< via3 >>
rect 6948 32124 7012 32128
rect 6948 32068 6952 32124
rect 6952 32068 7008 32124
rect 7008 32068 7012 32124
rect 6948 32064 7012 32068
rect 7028 32124 7092 32128
rect 7028 32068 7032 32124
rect 7032 32068 7088 32124
rect 7088 32068 7092 32124
rect 7028 32064 7092 32068
rect 7108 32124 7172 32128
rect 7108 32068 7112 32124
rect 7112 32068 7168 32124
rect 7168 32068 7172 32124
rect 7108 32064 7172 32068
rect 7188 32124 7252 32128
rect 7188 32068 7192 32124
rect 7192 32068 7248 32124
rect 7248 32068 7252 32124
rect 7188 32064 7252 32068
rect 14308 32124 14372 32128
rect 14308 32068 14312 32124
rect 14312 32068 14368 32124
rect 14368 32068 14372 32124
rect 14308 32064 14372 32068
rect 14388 32124 14452 32128
rect 14388 32068 14392 32124
rect 14392 32068 14448 32124
rect 14448 32068 14452 32124
rect 14388 32064 14452 32068
rect 14468 32124 14532 32128
rect 14468 32068 14472 32124
rect 14472 32068 14528 32124
rect 14528 32068 14532 32124
rect 14468 32064 14532 32068
rect 14548 32124 14612 32128
rect 14548 32068 14552 32124
rect 14552 32068 14608 32124
rect 14608 32068 14612 32124
rect 14548 32064 14612 32068
rect 21668 32124 21732 32128
rect 21668 32068 21672 32124
rect 21672 32068 21728 32124
rect 21728 32068 21732 32124
rect 21668 32064 21732 32068
rect 21748 32124 21812 32128
rect 21748 32068 21752 32124
rect 21752 32068 21808 32124
rect 21808 32068 21812 32124
rect 21748 32064 21812 32068
rect 21828 32124 21892 32128
rect 21828 32068 21832 32124
rect 21832 32068 21888 32124
rect 21888 32068 21892 32124
rect 21828 32064 21892 32068
rect 21908 32124 21972 32128
rect 21908 32068 21912 32124
rect 21912 32068 21968 32124
rect 21968 32068 21972 32124
rect 21908 32064 21972 32068
rect 29028 32124 29092 32128
rect 29028 32068 29032 32124
rect 29032 32068 29088 32124
rect 29088 32068 29092 32124
rect 29028 32064 29092 32068
rect 29108 32124 29172 32128
rect 29108 32068 29112 32124
rect 29112 32068 29168 32124
rect 29168 32068 29172 32124
rect 29108 32064 29172 32068
rect 29188 32124 29252 32128
rect 29188 32068 29192 32124
rect 29192 32068 29248 32124
rect 29248 32068 29252 32124
rect 29188 32064 29252 32068
rect 29268 32124 29332 32128
rect 29268 32068 29272 32124
rect 29272 32068 29328 32124
rect 29328 32068 29332 32124
rect 29268 32064 29332 32068
rect 13308 31860 13372 31924
rect 17724 31724 17788 31788
rect 6288 31580 6352 31584
rect 6288 31524 6292 31580
rect 6292 31524 6348 31580
rect 6348 31524 6352 31580
rect 6288 31520 6352 31524
rect 6368 31580 6432 31584
rect 6368 31524 6372 31580
rect 6372 31524 6428 31580
rect 6428 31524 6432 31580
rect 6368 31520 6432 31524
rect 6448 31580 6512 31584
rect 6448 31524 6452 31580
rect 6452 31524 6508 31580
rect 6508 31524 6512 31580
rect 6448 31520 6512 31524
rect 6528 31580 6592 31584
rect 6528 31524 6532 31580
rect 6532 31524 6588 31580
rect 6588 31524 6592 31580
rect 6528 31520 6592 31524
rect 13648 31580 13712 31584
rect 13648 31524 13652 31580
rect 13652 31524 13708 31580
rect 13708 31524 13712 31580
rect 13648 31520 13712 31524
rect 13728 31580 13792 31584
rect 13728 31524 13732 31580
rect 13732 31524 13788 31580
rect 13788 31524 13792 31580
rect 13728 31520 13792 31524
rect 13808 31580 13872 31584
rect 13808 31524 13812 31580
rect 13812 31524 13868 31580
rect 13868 31524 13872 31580
rect 13808 31520 13872 31524
rect 13888 31580 13952 31584
rect 13888 31524 13892 31580
rect 13892 31524 13948 31580
rect 13948 31524 13952 31580
rect 13888 31520 13952 31524
rect 21008 31580 21072 31584
rect 21008 31524 21012 31580
rect 21012 31524 21068 31580
rect 21068 31524 21072 31580
rect 21008 31520 21072 31524
rect 21088 31580 21152 31584
rect 21088 31524 21092 31580
rect 21092 31524 21148 31580
rect 21148 31524 21152 31580
rect 21088 31520 21152 31524
rect 21168 31580 21232 31584
rect 21168 31524 21172 31580
rect 21172 31524 21228 31580
rect 21228 31524 21232 31580
rect 21168 31520 21232 31524
rect 21248 31580 21312 31584
rect 21248 31524 21252 31580
rect 21252 31524 21308 31580
rect 21308 31524 21312 31580
rect 21248 31520 21312 31524
rect 28368 31580 28432 31584
rect 28368 31524 28372 31580
rect 28372 31524 28428 31580
rect 28428 31524 28432 31580
rect 28368 31520 28432 31524
rect 28448 31580 28512 31584
rect 28448 31524 28452 31580
rect 28452 31524 28508 31580
rect 28508 31524 28512 31580
rect 28448 31520 28512 31524
rect 28528 31580 28592 31584
rect 28528 31524 28532 31580
rect 28532 31524 28588 31580
rect 28588 31524 28592 31580
rect 28528 31520 28592 31524
rect 28608 31580 28672 31584
rect 28608 31524 28612 31580
rect 28612 31524 28668 31580
rect 28668 31524 28672 31580
rect 28608 31520 28672 31524
rect 6948 31036 7012 31040
rect 6948 30980 6952 31036
rect 6952 30980 7008 31036
rect 7008 30980 7012 31036
rect 6948 30976 7012 30980
rect 7028 31036 7092 31040
rect 7028 30980 7032 31036
rect 7032 30980 7088 31036
rect 7088 30980 7092 31036
rect 7028 30976 7092 30980
rect 7108 31036 7172 31040
rect 7108 30980 7112 31036
rect 7112 30980 7168 31036
rect 7168 30980 7172 31036
rect 7108 30976 7172 30980
rect 7188 31036 7252 31040
rect 7188 30980 7192 31036
rect 7192 30980 7248 31036
rect 7248 30980 7252 31036
rect 7188 30976 7252 30980
rect 14308 31036 14372 31040
rect 14308 30980 14312 31036
rect 14312 30980 14368 31036
rect 14368 30980 14372 31036
rect 14308 30976 14372 30980
rect 14388 31036 14452 31040
rect 14388 30980 14392 31036
rect 14392 30980 14448 31036
rect 14448 30980 14452 31036
rect 14388 30976 14452 30980
rect 14468 31036 14532 31040
rect 14468 30980 14472 31036
rect 14472 30980 14528 31036
rect 14528 30980 14532 31036
rect 14468 30976 14532 30980
rect 14548 31036 14612 31040
rect 14548 30980 14552 31036
rect 14552 30980 14608 31036
rect 14608 30980 14612 31036
rect 14548 30976 14612 30980
rect 21668 31036 21732 31040
rect 21668 30980 21672 31036
rect 21672 30980 21728 31036
rect 21728 30980 21732 31036
rect 21668 30976 21732 30980
rect 21748 31036 21812 31040
rect 21748 30980 21752 31036
rect 21752 30980 21808 31036
rect 21808 30980 21812 31036
rect 21748 30976 21812 30980
rect 21828 31036 21892 31040
rect 21828 30980 21832 31036
rect 21832 30980 21888 31036
rect 21888 30980 21892 31036
rect 21828 30976 21892 30980
rect 21908 31036 21972 31040
rect 21908 30980 21912 31036
rect 21912 30980 21968 31036
rect 21968 30980 21972 31036
rect 21908 30976 21972 30980
rect 29028 31036 29092 31040
rect 29028 30980 29032 31036
rect 29032 30980 29088 31036
rect 29088 30980 29092 31036
rect 29028 30976 29092 30980
rect 29108 31036 29172 31040
rect 29108 30980 29112 31036
rect 29112 30980 29168 31036
rect 29168 30980 29172 31036
rect 29108 30976 29172 30980
rect 29188 31036 29252 31040
rect 29188 30980 29192 31036
rect 29192 30980 29248 31036
rect 29248 30980 29252 31036
rect 29188 30976 29252 30980
rect 29268 31036 29332 31040
rect 29268 30980 29272 31036
rect 29272 30980 29328 31036
rect 29328 30980 29332 31036
rect 29268 30976 29332 30980
rect 6288 30492 6352 30496
rect 6288 30436 6292 30492
rect 6292 30436 6348 30492
rect 6348 30436 6352 30492
rect 6288 30432 6352 30436
rect 6368 30492 6432 30496
rect 6368 30436 6372 30492
rect 6372 30436 6428 30492
rect 6428 30436 6432 30492
rect 6368 30432 6432 30436
rect 6448 30492 6512 30496
rect 6448 30436 6452 30492
rect 6452 30436 6508 30492
rect 6508 30436 6512 30492
rect 6448 30432 6512 30436
rect 6528 30492 6592 30496
rect 6528 30436 6532 30492
rect 6532 30436 6588 30492
rect 6588 30436 6592 30492
rect 6528 30432 6592 30436
rect 13648 30492 13712 30496
rect 13648 30436 13652 30492
rect 13652 30436 13708 30492
rect 13708 30436 13712 30492
rect 13648 30432 13712 30436
rect 13728 30492 13792 30496
rect 13728 30436 13732 30492
rect 13732 30436 13788 30492
rect 13788 30436 13792 30492
rect 13728 30432 13792 30436
rect 13808 30492 13872 30496
rect 13808 30436 13812 30492
rect 13812 30436 13868 30492
rect 13868 30436 13872 30492
rect 13808 30432 13872 30436
rect 13888 30492 13952 30496
rect 13888 30436 13892 30492
rect 13892 30436 13948 30492
rect 13948 30436 13952 30492
rect 13888 30432 13952 30436
rect 21008 30492 21072 30496
rect 21008 30436 21012 30492
rect 21012 30436 21068 30492
rect 21068 30436 21072 30492
rect 21008 30432 21072 30436
rect 21088 30492 21152 30496
rect 21088 30436 21092 30492
rect 21092 30436 21148 30492
rect 21148 30436 21152 30492
rect 21088 30432 21152 30436
rect 21168 30492 21232 30496
rect 21168 30436 21172 30492
rect 21172 30436 21228 30492
rect 21228 30436 21232 30492
rect 21168 30432 21232 30436
rect 21248 30492 21312 30496
rect 21248 30436 21252 30492
rect 21252 30436 21308 30492
rect 21308 30436 21312 30492
rect 21248 30432 21312 30436
rect 28368 30492 28432 30496
rect 28368 30436 28372 30492
rect 28372 30436 28428 30492
rect 28428 30436 28432 30492
rect 28368 30432 28432 30436
rect 28448 30492 28512 30496
rect 28448 30436 28452 30492
rect 28452 30436 28508 30492
rect 28508 30436 28512 30492
rect 28448 30432 28512 30436
rect 28528 30492 28592 30496
rect 28528 30436 28532 30492
rect 28532 30436 28588 30492
rect 28588 30436 28592 30492
rect 28528 30432 28592 30436
rect 28608 30492 28672 30496
rect 28608 30436 28612 30492
rect 28612 30436 28668 30492
rect 28668 30436 28672 30492
rect 28608 30432 28672 30436
rect 6948 29948 7012 29952
rect 6948 29892 6952 29948
rect 6952 29892 7008 29948
rect 7008 29892 7012 29948
rect 6948 29888 7012 29892
rect 7028 29948 7092 29952
rect 7028 29892 7032 29948
rect 7032 29892 7088 29948
rect 7088 29892 7092 29948
rect 7028 29888 7092 29892
rect 7108 29948 7172 29952
rect 7108 29892 7112 29948
rect 7112 29892 7168 29948
rect 7168 29892 7172 29948
rect 7108 29888 7172 29892
rect 7188 29948 7252 29952
rect 7188 29892 7192 29948
rect 7192 29892 7248 29948
rect 7248 29892 7252 29948
rect 7188 29888 7252 29892
rect 14308 29948 14372 29952
rect 14308 29892 14312 29948
rect 14312 29892 14368 29948
rect 14368 29892 14372 29948
rect 14308 29888 14372 29892
rect 14388 29948 14452 29952
rect 14388 29892 14392 29948
rect 14392 29892 14448 29948
rect 14448 29892 14452 29948
rect 14388 29888 14452 29892
rect 14468 29948 14532 29952
rect 14468 29892 14472 29948
rect 14472 29892 14528 29948
rect 14528 29892 14532 29948
rect 14468 29888 14532 29892
rect 14548 29948 14612 29952
rect 14548 29892 14552 29948
rect 14552 29892 14608 29948
rect 14608 29892 14612 29948
rect 14548 29888 14612 29892
rect 21668 29948 21732 29952
rect 21668 29892 21672 29948
rect 21672 29892 21728 29948
rect 21728 29892 21732 29948
rect 21668 29888 21732 29892
rect 21748 29948 21812 29952
rect 21748 29892 21752 29948
rect 21752 29892 21808 29948
rect 21808 29892 21812 29948
rect 21748 29888 21812 29892
rect 21828 29948 21892 29952
rect 21828 29892 21832 29948
rect 21832 29892 21888 29948
rect 21888 29892 21892 29948
rect 21828 29888 21892 29892
rect 21908 29948 21972 29952
rect 21908 29892 21912 29948
rect 21912 29892 21968 29948
rect 21968 29892 21972 29948
rect 21908 29888 21972 29892
rect 29028 29948 29092 29952
rect 29028 29892 29032 29948
rect 29032 29892 29088 29948
rect 29088 29892 29092 29948
rect 29028 29888 29092 29892
rect 29108 29948 29172 29952
rect 29108 29892 29112 29948
rect 29112 29892 29168 29948
rect 29168 29892 29172 29948
rect 29108 29888 29172 29892
rect 29188 29948 29252 29952
rect 29188 29892 29192 29948
rect 29192 29892 29248 29948
rect 29248 29892 29252 29948
rect 29188 29888 29252 29892
rect 29268 29948 29332 29952
rect 29268 29892 29272 29948
rect 29272 29892 29328 29948
rect 29328 29892 29332 29948
rect 29268 29888 29332 29892
rect 6288 29404 6352 29408
rect 6288 29348 6292 29404
rect 6292 29348 6348 29404
rect 6348 29348 6352 29404
rect 6288 29344 6352 29348
rect 6368 29404 6432 29408
rect 6368 29348 6372 29404
rect 6372 29348 6428 29404
rect 6428 29348 6432 29404
rect 6368 29344 6432 29348
rect 6448 29404 6512 29408
rect 6448 29348 6452 29404
rect 6452 29348 6508 29404
rect 6508 29348 6512 29404
rect 6448 29344 6512 29348
rect 6528 29404 6592 29408
rect 6528 29348 6532 29404
rect 6532 29348 6588 29404
rect 6588 29348 6592 29404
rect 6528 29344 6592 29348
rect 13648 29404 13712 29408
rect 13648 29348 13652 29404
rect 13652 29348 13708 29404
rect 13708 29348 13712 29404
rect 13648 29344 13712 29348
rect 13728 29404 13792 29408
rect 13728 29348 13732 29404
rect 13732 29348 13788 29404
rect 13788 29348 13792 29404
rect 13728 29344 13792 29348
rect 13808 29404 13872 29408
rect 13808 29348 13812 29404
rect 13812 29348 13868 29404
rect 13868 29348 13872 29404
rect 13808 29344 13872 29348
rect 13888 29404 13952 29408
rect 13888 29348 13892 29404
rect 13892 29348 13948 29404
rect 13948 29348 13952 29404
rect 13888 29344 13952 29348
rect 21008 29404 21072 29408
rect 21008 29348 21012 29404
rect 21012 29348 21068 29404
rect 21068 29348 21072 29404
rect 21008 29344 21072 29348
rect 21088 29404 21152 29408
rect 21088 29348 21092 29404
rect 21092 29348 21148 29404
rect 21148 29348 21152 29404
rect 21088 29344 21152 29348
rect 21168 29404 21232 29408
rect 21168 29348 21172 29404
rect 21172 29348 21228 29404
rect 21228 29348 21232 29404
rect 21168 29344 21232 29348
rect 21248 29404 21312 29408
rect 21248 29348 21252 29404
rect 21252 29348 21308 29404
rect 21308 29348 21312 29404
rect 21248 29344 21312 29348
rect 28368 29404 28432 29408
rect 28368 29348 28372 29404
rect 28372 29348 28428 29404
rect 28428 29348 28432 29404
rect 28368 29344 28432 29348
rect 28448 29404 28512 29408
rect 28448 29348 28452 29404
rect 28452 29348 28508 29404
rect 28508 29348 28512 29404
rect 28448 29344 28512 29348
rect 28528 29404 28592 29408
rect 28528 29348 28532 29404
rect 28532 29348 28588 29404
rect 28588 29348 28592 29404
rect 28528 29344 28592 29348
rect 28608 29404 28672 29408
rect 28608 29348 28612 29404
rect 28612 29348 28668 29404
rect 28668 29348 28672 29404
rect 28608 29344 28672 29348
rect 6948 28860 7012 28864
rect 6948 28804 6952 28860
rect 6952 28804 7008 28860
rect 7008 28804 7012 28860
rect 6948 28800 7012 28804
rect 7028 28860 7092 28864
rect 7028 28804 7032 28860
rect 7032 28804 7088 28860
rect 7088 28804 7092 28860
rect 7028 28800 7092 28804
rect 7108 28860 7172 28864
rect 7108 28804 7112 28860
rect 7112 28804 7168 28860
rect 7168 28804 7172 28860
rect 7108 28800 7172 28804
rect 7188 28860 7252 28864
rect 7188 28804 7192 28860
rect 7192 28804 7248 28860
rect 7248 28804 7252 28860
rect 7188 28800 7252 28804
rect 14308 28860 14372 28864
rect 14308 28804 14312 28860
rect 14312 28804 14368 28860
rect 14368 28804 14372 28860
rect 14308 28800 14372 28804
rect 14388 28860 14452 28864
rect 14388 28804 14392 28860
rect 14392 28804 14448 28860
rect 14448 28804 14452 28860
rect 14388 28800 14452 28804
rect 14468 28860 14532 28864
rect 14468 28804 14472 28860
rect 14472 28804 14528 28860
rect 14528 28804 14532 28860
rect 14468 28800 14532 28804
rect 14548 28860 14612 28864
rect 14548 28804 14552 28860
rect 14552 28804 14608 28860
rect 14608 28804 14612 28860
rect 14548 28800 14612 28804
rect 21668 28860 21732 28864
rect 21668 28804 21672 28860
rect 21672 28804 21728 28860
rect 21728 28804 21732 28860
rect 21668 28800 21732 28804
rect 21748 28860 21812 28864
rect 21748 28804 21752 28860
rect 21752 28804 21808 28860
rect 21808 28804 21812 28860
rect 21748 28800 21812 28804
rect 21828 28860 21892 28864
rect 21828 28804 21832 28860
rect 21832 28804 21888 28860
rect 21888 28804 21892 28860
rect 21828 28800 21892 28804
rect 21908 28860 21972 28864
rect 21908 28804 21912 28860
rect 21912 28804 21968 28860
rect 21968 28804 21972 28860
rect 21908 28800 21972 28804
rect 29028 28860 29092 28864
rect 29028 28804 29032 28860
rect 29032 28804 29088 28860
rect 29088 28804 29092 28860
rect 29028 28800 29092 28804
rect 29108 28860 29172 28864
rect 29108 28804 29112 28860
rect 29112 28804 29168 28860
rect 29168 28804 29172 28860
rect 29108 28800 29172 28804
rect 29188 28860 29252 28864
rect 29188 28804 29192 28860
rect 29192 28804 29248 28860
rect 29248 28804 29252 28860
rect 29188 28800 29252 28804
rect 29268 28860 29332 28864
rect 29268 28804 29272 28860
rect 29272 28804 29328 28860
rect 29328 28804 29332 28860
rect 29268 28800 29332 28804
rect 6288 28316 6352 28320
rect 6288 28260 6292 28316
rect 6292 28260 6348 28316
rect 6348 28260 6352 28316
rect 6288 28256 6352 28260
rect 6368 28316 6432 28320
rect 6368 28260 6372 28316
rect 6372 28260 6428 28316
rect 6428 28260 6432 28316
rect 6368 28256 6432 28260
rect 6448 28316 6512 28320
rect 6448 28260 6452 28316
rect 6452 28260 6508 28316
rect 6508 28260 6512 28316
rect 6448 28256 6512 28260
rect 6528 28316 6592 28320
rect 6528 28260 6532 28316
rect 6532 28260 6588 28316
rect 6588 28260 6592 28316
rect 6528 28256 6592 28260
rect 13648 28316 13712 28320
rect 13648 28260 13652 28316
rect 13652 28260 13708 28316
rect 13708 28260 13712 28316
rect 13648 28256 13712 28260
rect 13728 28316 13792 28320
rect 13728 28260 13732 28316
rect 13732 28260 13788 28316
rect 13788 28260 13792 28316
rect 13728 28256 13792 28260
rect 13808 28316 13872 28320
rect 13808 28260 13812 28316
rect 13812 28260 13868 28316
rect 13868 28260 13872 28316
rect 13808 28256 13872 28260
rect 13888 28316 13952 28320
rect 13888 28260 13892 28316
rect 13892 28260 13948 28316
rect 13948 28260 13952 28316
rect 13888 28256 13952 28260
rect 21008 28316 21072 28320
rect 21008 28260 21012 28316
rect 21012 28260 21068 28316
rect 21068 28260 21072 28316
rect 21008 28256 21072 28260
rect 21088 28316 21152 28320
rect 21088 28260 21092 28316
rect 21092 28260 21148 28316
rect 21148 28260 21152 28316
rect 21088 28256 21152 28260
rect 21168 28316 21232 28320
rect 21168 28260 21172 28316
rect 21172 28260 21228 28316
rect 21228 28260 21232 28316
rect 21168 28256 21232 28260
rect 21248 28316 21312 28320
rect 21248 28260 21252 28316
rect 21252 28260 21308 28316
rect 21308 28260 21312 28316
rect 21248 28256 21312 28260
rect 28368 28316 28432 28320
rect 28368 28260 28372 28316
rect 28372 28260 28428 28316
rect 28428 28260 28432 28316
rect 28368 28256 28432 28260
rect 28448 28316 28512 28320
rect 28448 28260 28452 28316
rect 28452 28260 28508 28316
rect 28508 28260 28512 28316
rect 28448 28256 28512 28260
rect 28528 28316 28592 28320
rect 28528 28260 28532 28316
rect 28532 28260 28588 28316
rect 28588 28260 28592 28316
rect 28528 28256 28592 28260
rect 28608 28316 28672 28320
rect 28608 28260 28612 28316
rect 28612 28260 28668 28316
rect 28668 28260 28672 28316
rect 28608 28256 28672 28260
rect 16620 28112 16684 28116
rect 16620 28056 16634 28112
rect 16634 28056 16684 28112
rect 16620 28052 16684 28056
rect 6948 27772 7012 27776
rect 6948 27716 6952 27772
rect 6952 27716 7008 27772
rect 7008 27716 7012 27772
rect 6948 27712 7012 27716
rect 7028 27772 7092 27776
rect 7028 27716 7032 27772
rect 7032 27716 7088 27772
rect 7088 27716 7092 27772
rect 7028 27712 7092 27716
rect 7108 27772 7172 27776
rect 7108 27716 7112 27772
rect 7112 27716 7168 27772
rect 7168 27716 7172 27772
rect 7108 27712 7172 27716
rect 7188 27772 7252 27776
rect 7188 27716 7192 27772
rect 7192 27716 7248 27772
rect 7248 27716 7252 27772
rect 7188 27712 7252 27716
rect 14308 27772 14372 27776
rect 14308 27716 14312 27772
rect 14312 27716 14368 27772
rect 14368 27716 14372 27772
rect 14308 27712 14372 27716
rect 14388 27772 14452 27776
rect 14388 27716 14392 27772
rect 14392 27716 14448 27772
rect 14448 27716 14452 27772
rect 14388 27712 14452 27716
rect 14468 27772 14532 27776
rect 14468 27716 14472 27772
rect 14472 27716 14528 27772
rect 14528 27716 14532 27772
rect 14468 27712 14532 27716
rect 14548 27772 14612 27776
rect 14548 27716 14552 27772
rect 14552 27716 14608 27772
rect 14608 27716 14612 27772
rect 14548 27712 14612 27716
rect 21668 27772 21732 27776
rect 21668 27716 21672 27772
rect 21672 27716 21728 27772
rect 21728 27716 21732 27772
rect 21668 27712 21732 27716
rect 21748 27772 21812 27776
rect 21748 27716 21752 27772
rect 21752 27716 21808 27772
rect 21808 27716 21812 27772
rect 21748 27712 21812 27716
rect 21828 27772 21892 27776
rect 21828 27716 21832 27772
rect 21832 27716 21888 27772
rect 21888 27716 21892 27772
rect 21828 27712 21892 27716
rect 21908 27772 21972 27776
rect 21908 27716 21912 27772
rect 21912 27716 21968 27772
rect 21968 27716 21972 27772
rect 21908 27712 21972 27716
rect 29028 27772 29092 27776
rect 29028 27716 29032 27772
rect 29032 27716 29088 27772
rect 29088 27716 29092 27772
rect 29028 27712 29092 27716
rect 29108 27772 29172 27776
rect 29108 27716 29112 27772
rect 29112 27716 29168 27772
rect 29168 27716 29172 27772
rect 29108 27712 29172 27716
rect 29188 27772 29252 27776
rect 29188 27716 29192 27772
rect 29192 27716 29248 27772
rect 29248 27716 29252 27772
rect 29188 27712 29252 27716
rect 29268 27772 29332 27776
rect 29268 27716 29272 27772
rect 29272 27716 29328 27772
rect 29328 27716 29332 27772
rect 29268 27712 29332 27716
rect 11100 27704 11164 27708
rect 11100 27648 11114 27704
rect 11114 27648 11164 27704
rect 11100 27644 11164 27648
rect 6288 27228 6352 27232
rect 6288 27172 6292 27228
rect 6292 27172 6348 27228
rect 6348 27172 6352 27228
rect 6288 27168 6352 27172
rect 6368 27228 6432 27232
rect 6368 27172 6372 27228
rect 6372 27172 6428 27228
rect 6428 27172 6432 27228
rect 6368 27168 6432 27172
rect 6448 27228 6512 27232
rect 6448 27172 6452 27228
rect 6452 27172 6508 27228
rect 6508 27172 6512 27228
rect 6448 27168 6512 27172
rect 6528 27228 6592 27232
rect 6528 27172 6532 27228
rect 6532 27172 6588 27228
rect 6588 27172 6592 27228
rect 6528 27168 6592 27172
rect 13648 27228 13712 27232
rect 13648 27172 13652 27228
rect 13652 27172 13708 27228
rect 13708 27172 13712 27228
rect 13648 27168 13712 27172
rect 13728 27228 13792 27232
rect 13728 27172 13732 27228
rect 13732 27172 13788 27228
rect 13788 27172 13792 27228
rect 13728 27168 13792 27172
rect 13808 27228 13872 27232
rect 13808 27172 13812 27228
rect 13812 27172 13868 27228
rect 13868 27172 13872 27228
rect 13808 27168 13872 27172
rect 13888 27228 13952 27232
rect 13888 27172 13892 27228
rect 13892 27172 13948 27228
rect 13948 27172 13952 27228
rect 13888 27168 13952 27172
rect 21008 27228 21072 27232
rect 21008 27172 21012 27228
rect 21012 27172 21068 27228
rect 21068 27172 21072 27228
rect 21008 27168 21072 27172
rect 21088 27228 21152 27232
rect 21088 27172 21092 27228
rect 21092 27172 21148 27228
rect 21148 27172 21152 27228
rect 21088 27168 21152 27172
rect 21168 27228 21232 27232
rect 21168 27172 21172 27228
rect 21172 27172 21228 27228
rect 21228 27172 21232 27228
rect 21168 27168 21232 27172
rect 21248 27228 21312 27232
rect 21248 27172 21252 27228
rect 21252 27172 21308 27228
rect 21308 27172 21312 27228
rect 21248 27168 21312 27172
rect 28368 27228 28432 27232
rect 28368 27172 28372 27228
rect 28372 27172 28428 27228
rect 28428 27172 28432 27228
rect 28368 27168 28432 27172
rect 28448 27228 28512 27232
rect 28448 27172 28452 27228
rect 28452 27172 28508 27228
rect 28508 27172 28512 27228
rect 28448 27168 28512 27172
rect 28528 27228 28592 27232
rect 28528 27172 28532 27228
rect 28532 27172 28588 27228
rect 28588 27172 28592 27228
rect 28528 27168 28592 27172
rect 28608 27228 28672 27232
rect 28608 27172 28612 27228
rect 28612 27172 28668 27228
rect 28668 27172 28672 27228
rect 28608 27168 28672 27172
rect 6948 26684 7012 26688
rect 6948 26628 6952 26684
rect 6952 26628 7008 26684
rect 7008 26628 7012 26684
rect 6948 26624 7012 26628
rect 7028 26684 7092 26688
rect 7028 26628 7032 26684
rect 7032 26628 7088 26684
rect 7088 26628 7092 26684
rect 7028 26624 7092 26628
rect 7108 26684 7172 26688
rect 7108 26628 7112 26684
rect 7112 26628 7168 26684
rect 7168 26628 7172 26684
rect 7108 26624 7172 26628
rect 7188 26684 7252 26688
rect 7188 26628 7192 26684
rect 7192 26628 7248 26684
rect 7248 26628 7252 26684
rect 7188 26624 7252 26628
rect 14308 26684 14372 26688
rect 14308 26628 14312 26684
rect 14312 26628 14368 26684
rect 14368 26628 14372 26684
rect 14308 26624 14372 26628
rect 14388 26684 14452 26688
rect 14388 26628 14392 26684
rect 14392 26628 14448 26684
rect 14448 26628 14452 26684
rect 14388 26624 14452 26628
rect 14468 26684 14532 26688
rect 14468 26628 14472 26684
rect 14472 26628 14528 26684
rect 14528 26628 14532 26684
rect 14468 26624 14532 26628
rect 14548 26684 14612 26688
rect 14548 26628 14552 26684
rect 14552 26628 14608 26684
rect 14608 26628 14612 26684
rect 14548 26624 14612 26628
rect 21668 26684 21732 26688
rect 21668 26628 21672 26684
rect 21672 26628 21728 26684
rect 21728 26628 21732 26684
rect 21668 26624 21732 26628
rect 21748 26684 21812 26688
rect 21748 26628 21752 26684
rect 21752 26628 21808 26684
rect 21808 26628 21812 26684
rect 21748 26624 21812 26628
rect 21828 26684 21892 26688
rect 21828 26628 21832 26684
rect 21832 26628 21888 26684
rect 21888 26628 21892 26684
rect 21828 26624 21892 26628
rect 21908 26684 21972 26688
rect 21908 26628 21912 26684
rect 21912 26628 21968 26684
rect 21968 26628 21972 26684
rect 21908 26624 21972 26628
rect 29028 26684 29092 26688
rect 29028 26628 29032 26684
rect 29032 26628 29088 26684
rect 29088 26628 29092 26684
rect 29028 26624 29092 26628
rect 29108 26684 29172 26688
rect 29108 26628 29112 26684
rect 29112 26628 29168 26684
rect 29168 26628 29172 26684
rect 29108 26624 29172 26628
rect 29188 26684 29252 26688
rect 29188 26628 29192 26684
rect 29192 26628 29248 26684
rect 29248 26628 29252 26684
rect 29188 26624 29252 26628
rect 29268 26684 29332 26688
rect 29268 26628 29272 26684
rect 29272 26628 29328 26684
rect 29328 26628 29332 26684
rect 29268 26624 29332 26628
rect 6288 26140 6352 26144
rect 6288 26084 6292 26140
rect 6292 26084 6348 26140
rect 6348 26084 6352 26140
rect 6288 26080 6352 26084
rect 6368 26140 6432 26144
rect 6368 26084 6372 26140
rect 6372 26084 6428 26140
rect 6428 26084 6432 26140
rect 6368 26080 6432 26084
rect 6448 26140 6512 26144
rect 6448 26084 6452 26140
rect 6452 26084 6508 26140
rect 6508 26084 6512 26140
rect 6448 26080 6512 26084
rect 6528 26140 6592 26144
rect 6528 26084 6532 26140
rect 6532 26084 6588 26140
rect 6588 26084 6592 26140
rect 6528 26080 6592 26084
rect 13648 26140 13712 26144
rect 13648 26084 13652 26140
rect 13652 26084 13708 26140
rect 13708 26084 13712 26140
rect 13648 26080 13712 26084
rect 13728 26140 13792 26144
rect 13728 26084 13732 26140
rect 13732 26084 13788 26140
rect 13788 26084 13792 26140
rect 13728 26080 13792 26084
rect 13808 26140 13872 26144
rect 13808 26084 13812 26140
rect 13812 26084 13868 26140
rect 13868 26084 13872 26140
rect 13808 26080 13872 26084
rect 13888 26140 13952 26144
rect 13888 26084 13892 26140
rect 13892 26084 13948 26140
rect 13948 26084 13952 26140
rect 13888 26080 13952 26084
rect 21008 26140 21072 26144
rect 21008 26084 21012 26140
rect 21012 26084 21068 26140
rect 21068 26084 21072 26140
rect 21008 26080 21072 26084
rect 21088 26140 21152 26144
rect 21088 26084 21092 26140
rect 21092 26084 21148 26140
rect 21148 26084 21152 26140
rect 21088 26080 21152 26084
rect 21168 26140 21232 26144
rect 21168 26084 21172 26140
rect 21172 26084 21228 26140
rect 21228 26084 21232 26140
rect 21168 26080 21232 26084
rect 21248 26140 21312 26144
rect 21248 26084 21252 26140
rect 21252 26084 21308 26140
rect 21308 26084 21312 26140
rect 21248 26080 21312 26084
rect 28368 26140 28432 26144
rect 28368 26084 28372 26140
rect 28372 26084 28428 26140
rect 28428 26084 28432 26140
rect 28368 26080 28432 26084
rect 28448 26140 28512 26144
rect 28448 26084 28452 26140
rect 28452 26084 28508 26140
rect 28508 26084 28512 26140
rect 28448 26080 28512 26084
rect 28528 26140 28592 26144
rect 28528 26084 28532 26140
rect 28532 26084 28588 26140
rect 28588 26084 28592 26140
rect 28528 26080 28592 26084
rect 28608 26140 28672 26144
rect 28608 26084 28612 26140
rect 28612 26084 28668 26140
rect 28668 26084 28672 26140
rect 28608 26080 28672 26084
rect 11284 25800 11348 25804
rect 11284 25744 11334 25800
rect 11334 25744 11348 25800
rect 11284 25740 11348 25744
rect 6948 25596 7012 25600
rect 6948 25540 6952 25596
rect 6952 25540 7008 25596
rect 7008 25540 7012 25596
rect 6948 25536 7012 25540
rect 7028 25596 7092 25600
rect 7028 25540 7032 25596
rect 7032 25540 7088 25596
rect 7088 25540 7092 25596
rect 7028 25536 7092 25540
rect 7108 25596 7172 25600
rect 7108 25540 7112 25596
rect 7112 25540 7168 25596
rect 7168 25540 7172 25596
rect 7108 25536 7172 25540
rect 7188 25596 7252 25600
rect 7188 25540 7192 25596
rect 7192 25540 7248 25596
rect 7248 25540 7252 25596
rect 7188 25536 7252 25540
rect 14308 25596 14372 25600
rect 14308 25540 14312 25596
rect 14312 25540 14368 25596
rect 14368 25540 14372 25596
rect 14308 25536 14372 25540
rect 14388 25596 14452 25600
rect 14388 25540 14392 25596
rect 14392 25540 14448 25596
rect 14448 25540 14452 25596
rect 14388 25536 14452 25540
rect 14468 25596 14532 25600
rect 14468 25540 14472 25596
rect 14472 25540 14528 25596
rect 14528 25540 14532 25596
rect 14468 25536 14532 25540
rect 14548 25596 14612 25600
rect 14548 25540 14552 25596
rect 14552 25540 14608 25596
rect 14608 25540 14612 25596
rect 14548 25536 14612 25540
rect 21668 25596 21732 25600
rect 21668 25540 21672 25596
rect 21672 25540 21728 25596
rect 21728 25540 21732 25596
rect 21668 25536 21732 25540
rect 21748 25596 21812 25600
rect 21748 25540 21752 25596
rect 21752 25540 21808 25596
rect 21808 25540 21812 25596
rect 21748 25536 21812 25540
rect 21828 25596 21892 25600
rect 21828 25540 21832 25596
rect 21832 25540 21888 25596
rect 21888 25540 21892 25596
rect 21828 25536 21892 25540
rect 21908 25596 21972 25600
rect 21908 25540 21912 25596
rect 21912 25540 21968 25596
rect 21968 25540 21972 25596
rect 21908 25536 21972 25540
rect 29028 25596 29092 25600
rect 29028 25540 29032 25596
rect 29032 25540 29088 25596
rect 29088 25540 29092 25596
rect 29028 25536 29092 25540
rect 29108 25596 29172 25600
rect 29108 25540 29112 25596
rect 29112 25540 29168 25596
rect 29168 25540 29172 25596
rect 29108 25536 29172 25540
rect 29188 25596 29252 25600
rect 29188 25540 29192 25596
rect 29192 25540 29248 25596
rect 29248 25540 29252 25596
rect 29188 25536 29252 25540
rect 29268 25596 29332 25600
rect 29268 25540 29272 25596
rect 29272 25540 29328 25596
rect 29328 25540 29332 25596
rect 29268 25536 29332 25540
rect 6288 25052 6352 25056
rect 6288 24996 6292 25052
rect 6292 24996 6348 25052
rect 6348 24996 6352 25052
rect 6288 24992 6352 24996
rect 6368 25052 6432 25056
rect 6368 24996 6372 25052
rect 6372 24996 6428 25052
rect 6428 24996 6432 25052
rect 6368 24992 6432 24996
rect 6448 25052 6512 25056
rect 6448 24996 6452 25052
rect 6452 24996 6508 25052
rect 6508 24996 6512 25052
rect 6448 24992 6512 24996
rect 6528 25052 6592 25056
rect 6528 24996 6532 25052
rect 6532 24996 6588 25052
rect 6588 24996 6592 25052
rect 6528 24992 6592 24996
rect 13648 25052 13712 25056
rect 13648 24996 13652 25052
rect 13652 24996 13708 25052
rect 13708 24996 13712 25052
rect 13648 24992 13712 24996
rect 13728 25052 13792 25056
rect 13728 24996 13732 25052
rect 13732 24996 13788 25052
rect 13788 24996 13792 25052
rect 13728 24992 13792 24996
rect 13808 25052 13872 25056
rect 13808 24996 13812 25052
rect 13812 24996 13868 25052
rect 13868 24996 13872 25052
rect 13808 24992 13872 24996
rect 13888 25052 13952 25056
rect 13888 24996 13892 25052
rect 13892 24996 13948 25052
rect 13948 24996 13952 25052
rect 13888 24992 13952 24996
rect 21008 25052 21072 25056
rect 21008 24996 21012 25052
rect 21012 24996 21068 25052
rect 21068 24996 21072 25052
rect 21008 24992 21072 24996
rect 21088 25052 21152 25056
rect 21088 24996 21092 25052
rect 21092 24996 21148 25052
rect 21148 24996 21152 25052
rect 21088 24992 21152 24996
rect 21168 25052 21232 25056
rect 21168 24996 21172 25052
rect 21172 24996 21228 25052
rect 21228 24996 21232 25052
rect 21168 24992 21232 24996
rect 21248 25052 21312 25056
rect 21248 24996 21252 25052
rect 21252 24996 21308 25052
rect 21308 24996 21312 25052
rect 21248 24992 21312 24996
rect 28368 25052 28432 25056
rect 28368 24996 28372 25052
rect 28372 24996 28428 25052
rect 28428 24996 28432 25052
rect 28368 24992 28432 24996
rect 28448 25052 28512 25056
rect 28448 24996 28452 25052
rect 28452 24996 28508 25052
rect 28508 24996 28512 25052
rect 28448 24992 28512 24996
rect 28528 25052 28592 25056
rect 28528 24996 28532 25052
rect 28532 24996 28588 25052
rect 28588 24996 28592 25052
rect 28528 24992 28592 24996
rect 28608 25052 28672 25056
rect 28608 24996 28612 25052
rect 28612 24996 28668 25052
rect 28668 24996 28672 25052
rect 28608 24992 28672 24996
rect 6948 24508 7012 24512
rect 6948 24452 6952 24508
rect 6952 24452 7008 24508
rect 7008 24452 7012 24508
rect 6948 24448 7012 24452
rect 7028 24508 7092 24512
rect 7028 24452 7032 24508
rect 7032 24452 7088 24508
rect 7088 24452 7092 24508
rect 7028 24448 7092 24452
rect 7108 24508 7172 24512
rect 7108 24452 7112 24508
rect 7112 24452 7168 24508
rect 7168 24452 7172 24508
rect 7108 24448 7172 24452
rect 7188 24508 7252 24512
rect 7188 24452 7192 24508
rect 7192 24452 7248 24508
rect 7248 24452 7252 24508
rect 7188 24448 7252 24452
rect 14308 24508 14372 24512
rect 14308 24452 14312 24508
rect 14312 24452 14368 24508
rect 14368 24452 14372 24508
rect 14308 24448 14372 24452
rect 14388 24508 14452 24512
rect 14388 24452 14392 24508
rect 14392 24452 14448 24508
rect 14448 24452 14452 24508
rect 14388 24448 14452 24452
rect 14468 24508 14532 24512
rect 14468 24452 14472 24508
rect 14472 24452 14528 24508
rect 14528 24452 14532 24508
rect 14468 24448 14532 24452
rect 14548 24508 14612 24512
rect 14548 24452 14552 24508
rect 14552 24452 14608 24508
rect 14608 24452 14612 24508
rect 14548 24448 14612 24452
rect 21668 24508 21732 24512
rect 21668 24452 21672 24508
rect 21672 24452 21728 24508
rect 21728 24452 21732 24508
rect 21668 24448 21732 24452
rect 21748 24508 21812 24512
rect 21748 24452 21752 24508
rect 21752 24452 21808 24508
rect 21808 24452 21812 24508
rect 21748 24448 21812 24452
rect 21828 24508 21892 24512
rect 21828 24452 21832 24508
rect 21832 24452 21888 24508
rect 21888 24452 21892 24508
rect 21828 24448 21892 24452
rect 21908 24508 21972 24512
rect 21908 24452 21912 24508
rect 21912 24452 21968 24508
rect 21968 24452 21972 24508
rect 21908 24448 21972 24452
rect 29028 24508 29092 24512
rect 29028 24452 29032 24508
rect 29032 24452 29088 24508
rect 29088 24452 29092 24508
rect 29028 24448 29092 24452
rect 29108 24508 29172 24512
rect 29108 24452 29112 24508
rect 29112 24452 29168 24508
rect 29168 24452 29172 24508
rect 29108 24448 29172 24452
rect 29188 24508 29252 24512
rect 29188 24452 29192 24508
rect 29192 24452 29248 24508
rect 29248 24452 29252 24508
rect 29188 24448 29252 24452
rect 29268 24508 29332 24512
rect 29268 24452 29272 24508
rect 29272 24452 29328 24508
rect 29328 24452 29332 24508
rect 29268 24448 29332 24452
rect 6288 23964 6352 23968
rect 6288 23908 6292 23964
rect 6292 23908 6348 23964
rect 6348 23908 6352 23964
rect 6288 23904 6352 23908
rect 6368 23964 6432 23968
rect 6368 23908 6372 23964
rect 6372 23908 6428 23964
rect 6428 23908 6432 23964
rect 6368 23904 6432 23908
rect 6448 23964 6512 23968
rect 6448 23908 6452 23964
rect 6452 23908 6508 23964
rect 6508 23908 6512 23964
rect 6448 23904 6512 23908
rect 6528 23964 6592 23968
rect 6528 23908 6532 23964
rect 6532 23908 6588 23964
rect 6588 23908 6592 23964
rect 6528 23904 6592 23908
rect 13648 23964 13712 23968
rect 13648 23908 13652 23964
rect 13652 23908 13708 23964
rect 13708 23908 13712 23964
rect 13648 23904 13712 23908
rect 13728 23964 13792 23968
rect 13728 23908 13732 23964
rect 13732 23908 13788 23964
rect 13788 23908 13792 23964
rect 13728 23904 13792 23908
rect 13808 23964 13872 23968
rect 13808 23908 13812 23964
rect 13812 23908 13868 23964
rect 13868 23908 13872 23964
rect 13808 23904 13872 23908
rect 13888 23964 13952 23968
rect 13888 23908 13892 23964
rect 13892 23908 13948 23964
rect 13948 23908 13952 23964
rect 13888 23904 13952 23908
rect 21008 23964 21072 23968
rect 21008 23908 21012 23964
rect 21012 23908 21068 23964
rect 21068 23908 21072 23964
rect 21008 23904 21072 23908
rect 21088 23964 21152 23968
rect 21088 23908 21092 23964
rect 21092 23908 21148 23964
rect 21148 23908 21152 23964
rect 21088 23904 21152 23908
rect 21168 23964 21232 23968
rect 21168 23908 21172 23964
rect 21172 23908 21228 23964
rect 21228 23908 21232 23964
rect 21168 23904 21232 23908
rect 21248 23964 21312 23968
rect 21248 23908 21252 23964
rect 21252 23908 21308 23964
rect 21308 23908 21312 23964
rect 21248 23904 21312 23908
rect 28368 23964 28432 23968
rect 28368 23908 28372 23964
rect 28372 23908 28428 23964
rect 28428 23908 28432 23964
rect 28368 23904 28432 23908
rect 28448 23964 28512 23968
rect 28448 23908 28452 23964
rect 28452 23908 28508 23964
rect 28508 23908 28512 23964
rect 28448 23904 28512 23908
rect 28528 23964 28592 23968
rect 28528 23908 28532 23964
rect 28532 23908 28588 23964
rect 28588 23908 28592 23964
rect 28528 23904 28592 23908
rect 28608 23964 28672 23968
rect 28608 23908 28612 23964
rect 28612 23908 28668 23964
rect 28668 23908 28672 23964
rect 28608 23904 28672 23908
rect 13124 23700 13188 23764
rect 6948 23420 7012 23424
rect 6948 23364 6952 23420
rect 6952 23364 7008 23420
rect 7008 23364 7012 23420
rect 6948 23360 7012 23364
rect 7028 23420 7092 23424
rect 7028 23364 7032 23420
rect 7032 23364 7088 23420
rect 7088 23364 7092 23420
rect 7028 23360 7092 23364
rect 7108 23420 7172 23424
rect 7108 23364 7112 23420
rect 7112 23364 7168 23420
rect 7168 23364 7172 23420
rect 7108 23360 7172 23364
rect 7188 23420 7252 23424
rect 7188 23364 7192 23420
rect 7192 23364 7248 23420
rect 7248 23364 7252 23420
rect 7188 23360 7252 23364
rect 14308 23420 14372 23424
rect 14308 23364 14312 23420
rect 14312 23364 14368 23420
rect 14368 23364 14372 23420
rect 14308 23360 14372 23364
rect 14388 23420 14452 23424
rect 14388 23364 14392 23420
rect 14392 23364 14448 23420
rect 14448 23364 14452 23420
rect 14388 23360 14452 23364
rect 14468 23420 14532 23424
rect 14468 23364 14472 23420
rect 14472 23364 14528 23420
rect 14528 23364 14532 23420
rect 14468 23360 14532 23364
rect 14548 23420 14612 23424
rect 14548 23364 14552 23420
rect 14552 23364 14608 23420
rect 14608 23364 14612 23420
rect 14548 23360 14612 23364
rect 21668 23420 21732 23424
rect 21668 23364 21672 23420
rect 21672 23364 21728 23420
rect 21728 23364 21732 23420
rect 21668 23360 21732 23364
rect 21748 23420 21812 23424
rect 21748 23364 21752 23420
rect 21752 23364 21808 23420
rect 21808 23364 21812 23420
rect 21748 23360 21812 23364
rect 21828 23420 21892 23424
rect 21828 23364 21832 23420
rect 21832 23364 21888 23420
rect 21888 23364 21892 23420
rect 21828 23360 21892 23364
rect 21908 23420 21972 23424
rect 21908 23364 21912 23420
rect 21912 23364 21968 23420
rect 21968 23364 21972 23420
rect 21908 23360 21972 23364
rect 29028 23420 29092 23424
rect 29028 23364 29032 23420
rect 29032 23364 29088 23420
rect 29088 23364 29092 23420
rect 29028 23360 29092 23364
rect 29108 23420 29172 23424
rect 29108 23364 29112 23420
rect 29112 23364 29168 23420
rect 29168 23364 29172 23420
rect 29108 23360 29172 23364
rect 29188 23420 29252 23424
rect 29188 23364 29192 23420
rect 29192 23364 29248 23420
rect 29248 23364 29252 23420
rect 29188 23360 29252 23364
rect 29268 23420 29332 23424
rect 29268 23364 29272 23420
rect 29272 23364 29328 23420
rect 29328 23364 29332 23420
rect 29268 23360 29332 23364
rect 6288 22876 6352 22880
rect 6288 22820 6292 22876
rect 6292 22820 6348 22876
rect 6348 22820 6352 22876
rect 6288 22816 6352 22820
rect 6368 22876 6432 22880
rect 6368 22820 6372 22876
rect 6372 22820 6428 22876
rect 6428 22820 6432 22876
rect 6368 22816 6432 22820
rect 6448 22876 6512 22880
rect 6448 22820 6452 22876
rect 6452 22820 6508 22876
rect 6508 22820 6512 22876
rect 6448 22816 6512 22820
rect 6528 22876 6592 22880
rect 6528 22820 6532 22876
rect 6532 22820 6588 22876
rect 6588 22820 6592 22876
rect 6528 22816 6592 22820
rect 13648 22876 13712 22880
rect 13648 22820 13652 22876
rect 13652 22820 13708 22876
rect 13708 22820 13712 22876
rect 13648 22816 13712 22820
rect 13728 22876 13792 22880
rect 13728 22820 13732 22876
rect 13732 22820 13788 22876
rect 13788 22820 13792 22876
rect 13728 22816 13792 22820
rect 13808 22876 13872 22880
rect 13808 22820 13812 22876
rect 13812 22820 13868 22876
rect 13868 22820 13872 22876
rect 13808 22816 13872 22820
rect 13888 22876 13952 22880
rect 13888 22820 13892 22876
rect 13892 22820 13948 22876
rect 13948 22820 13952 22876
rect 13888 22816 13952 22820
rect 21008 22876 21072 22880
rect 21008 22820 21012 22876
rect 21012 22820 21068 22876
rect 21068 22820 21072 22876
rect 21008 22816 21072 22820
rect 21088 22876 21152 22880
rect 21088 22820 21092 22876
rect 21092 22820 21148 22876
rect 21148 22820 21152 22876
rect 21088 22816 21152 22820
rect 21168 22876 21232 22880
rect 21168 22820 21172 22876
rect 21172 22820 21228 22876
rect 21228 22820 21232 22876
rect 21168 22816 21232 22820
rect 21248 22876 21312 22880
rect 21248 22820 21252 22876
rect 21252 22820 21308 22876
rect 21308 22820 21312 22876
rect 21248 22816 21312 22820
rect 28368 22876 28432 22880
rect 28368 22820 28372 22876
rect 28372 22820 28428 22876
rect 28428 22820 28432 22876
rect 28368 22816 28432 22820
rect 28448 22876 28512 22880
rect 28448 22820 28452 22876
rect 28452 22820 28508 22876
rect 28508 22820 28512 22876
rect 28448 22816 28512 22820
rect 28528 22876 28592 22880
rect 28528 22820 28532 22876
rect 28532 22820 28588 22876
rect 28588 22820 28592 22876
rect 28528 22816 28592 22820
rect 28608 22876 28672 22880
rect 28608 22820 28612 22876
rect 28612 22820 28668 22876
rect 28668 22820 28672 22876
rect 28608 22816 28672 22820
rect 6948 22332 7012 22336
rect 6948 22276 6952 22332
rect 6952 22276 7008 22332
rect 7008 22276 7012 22332
rect 6948 22272 7012 22276
rect 7028 22332 7092 22336
rect 7028 22276 7032 22332
rect 7032 22276 7088 22332
rect 7088 22276 7092 22332
rect 7028 22272 7092 22276
rect 7108 22332 7172 22336
rect 7108 22276 7112 22332
rect 7112 22276 7168 22332
rect 7168 22276 7172 22332
rect 7108 22272 7172 22276
rect 7188 22332 7252 22336
rect 7188 22276 7192 22332
rect 7192 22276 7248 22332
rect 7248 22276 7252 22332
rect 7188 22272 7252 22276
rect 14308 22332 14372 22336
rect 14308 22276 14312 22332
rect 14312 22276 14368 22332
rect 14368 22276 14372 22332
rect 14308 22272 14372 22276
rect 14388 22332 14452 22336
rect 14388 22276 14392 22332
rect 14392 22276 14448 22332
rect 14448 22276 14452 22332
rect 14388 22272 14452 22276
rect 14468 22332 14532 22336
rect 14468 22276 14472 22332
rect 14472 22276 14528 22332
rect 14528 22276 14532 22332
rect 14468 22272 14532 22276
rect 14548 22332 14612 22336
rect 14548 22276 14552 22332
rect 14552 22276 14608 22332
rect 14608 22276 14612 22332
rect 14548 22272 14612 22276
rect 21668 22332 21732 22336
rect 21668 22276 21672 22332
rect 21672 22276 21728 22332
rect 21728 22276 21732 22332
rect 21668 22272 21732 22276
rect 21748 22332 21812 22336
rect 21748 22276 21752 22332
rect 21752 22276 21808 22332
rect 21808 22276 21812 22332
rect 21748 22272 21812 22276
rect 21828 22332 21892 22336
rect 21828 22276 21832 22332
rect 21832 22276 21888 22332
rect 21888 22276 21892 22332
rect 21828 22272 21892 22276
rect 21908 22332 21972 22336
rect 21908 22276 21912 22332
rect 21912 22276 21968 22332
rect 21968 22276 21972 22332
rect 21908 22272 21972 22276
rect 29028 22332 29092 22336
rect 29028 22276 29032 22332
rect 29032 22276 29088 22332
rect 29088 22276 29092 22332
rect 29028 22272 29092 22276
rect 29108 22332 29172 22336
rect 29108 22276 29112 22332
rect 29112 22276 29168 22332
rect 29168 22276 29172 22332
rect 29108 22272 29172 22276
rect 29188 22332 29252 22336
rect 29188 22276 29192 22332
rect 29192 22276 29248 22332
rect 29248 22276 29252 22332
rect 29188 22272 29252 22276
rect 29268 22332 29332 22336
rect 29268 22276 29272 22332
rect 29272 22276 29328 22332
rect 29328 22276 29332 22332
rect 29268 22272 29332 22276
rect 6288 21788 6352 21792
rect 6288 21732 6292 21788
rect 6292 21732 6348 21788
rect 6348 21732 6352 21788
rect 6288 21728 6352 21732
rect 6368 21788 6432 21792
rect 6368 21732 6372 21788
rect 6372 21732 6428 21788
rect 6428 21732 6432 21788
rect 6368 21728 6432 21732
rect 6448 21788 6512 21792
rect 6448 21732 6452 21788
rect 6452 21732 6508 21788
rect 6508 21732 6512 21788
rect 6448 21728 6512 21732
rect 6528 21788 6592 21792
rect 6528 21732 6532 21788
rect 6532 21732 6588 21788
rect 6588 21732 6592 21788
rect 6528 21728 6592 21732
rect 13648 21788 13712 21792
rect 13648 21732 13652 21788
rect 13652 21732 13708 21788
rect 13708 21732 13712 21788
rect 13648 21728 13712 21732
rect 13728 21788 13792 21792
rect 13728 21732 13732 21788
rect 13732 21732 13788 21788
rect 13788 21732 13792 21788
rect 13728 21728 13792 21732
rect 13808 21788 13872 21792
rect 13808 21732 13812 21788
rect 13812 21732 13868 21788
rect 13868 21732 13872 21788
rect 13808 21728 13872 21732
rect 13888 21788 13952 21792
rect 13888 21732 13892 21788
rect 13892 21732 13948 21788
rect 13948 21732 13952 21788
rect 13888 21728 13952 21732
rect 21008 21788 21072 21792
rect 21008 21732 21012 21788
rect 21012 21732 21068 21788
rect 21068 21732 21072 21788
rect 21008 21728 21072 21732
rect 21088 21788 21152 21792
rect 21088 21732 21092 21788
rect 21092 21732 21148 21788
rect 21148 21732 21152 21788
rect 21088 21728 21152 21732
rect 21168 21788 21232 21792
rect 21168 21732 21172 21788
rect 21172 21732 21228 21788
rect 21228 21732 21232 21788
rect 21168 21728 21232 21732
rect 21248 21788 21312 21792
rect 21248 21732 21252 21788
rect 21252 21732 21308 21788
rect 21308 21732 21312 21788
rect 21248 21728 21312 21732
rect 28368 21788 28432 21792
rect 28368 21732 28372 21788
rect 28372 21732 28428 21788
rect 28428 21732 28432 21788
rect 28368 21728 28432 21732
rect 28448 21788 28512 21792
rect 28448 21732 28452 21788
rect 28452 21732 28508 21788
rect 28508 21732 28512 21788
rect 28448 21728 28512 21732
rect 28528 21788 28592 21792
rect 28528 21732 28532 21788
rect 28532 21732 28588 21788
rect 28588 21732 28592 21788
rect 28528 21728 28592 21732
rect 28608 21788 28672 21792
rect 28608 21732 28612 21788
rect 28612 21732 28668 21788
rect 28668 21732 28672 21788
rect 28608 21728 28672 21732
rect 6948 21244 7012 21248
rect 6948 21188 6952 21244
rect 6952 21188 7008 21244
rect 7008 21188 7012 21244
rect 6948 21184 7012 21188
rect 7028 21244 7092 21248
rect 7028 21188 7032 21244
rect 7032 21188 7088 21244
rect 7088 21188 7092 21244
rect 7028 21184 7092 21188
rect 7108 21244 7172 21248
rect 7108 21188 7112 21244
rect 7112 21188 7168 21244
rect 7168 21188 7172 21244
rect 7108 21184 7172 21188
rect 7188 21244 7252 21248
rect 7188 21188 7192 21244
rect 7192 21188 7248 21244
rect 7248 21188 7252 21244
rect 7188 21184 7252 21188
rect 14308 21244 14372 21248
rect 14308 21188 14312 21244
rect 14312 21188 14368 21244
rect 14368 21188 14372 21244
rect 14308 21184 14372 21188
rect 14388 21244 14452 21248
rect 14388 21188 14392 21244
rect 14392 21188 14448 21244
rect 14448 21188 14452 21244
rect 14388 21184 14452 21188
rect 14468 21244 14532 21248
rect 14468 21188 14472 21244
rect 14472 21188 14528 21244
rect 14528 21188 14532 21244
rect 14468 21184 14532 21188
rect 14548 21244 14612 21248
rect 14548 21188 14552 21244
rect 14552 21188 14608 21244
rect 14608 21188 14612 21244
rect 14548 21184 14612 21188
rect 21668 21244 21732 21248
rect 21668 21188 21672 21244
rect 21672 21188 21728 21244
rect 21728 21188 21732 21244
rect 21668 21184 21732 21188
rect 21748 21244 21812 21248
rect 21748 21188 21752 21244
rect 21752 21188 21808 21244
rect 21808 21188 21812 21244
rect 21748 21184 21812 21188
rect 21828 21244 21892 21248
rect 21828 21188 21832 21244
rect 21832 21188 21888 21244
rect 21888 21188 21892 21244
rect 21828 21184 21892 21188
rect 21908 21244 21972 21248
rect 21908 21188 21912 21244
rect 21912 21188 21968 21244
rect 21968 21188 21972 21244
rect 21908 21184 21972 21188
rect 29028 21244 29092 21248
rect 29028 21188 29032 21244
rect 29032 21188 29088 21244
rect 29088 21188 29092 21244
rect 29028 21184 29092 21188
rect 29108 21244 29172 21248
rect 29108 21188 29112 21244
rect 29112 21188 29168 21244
rect 29168 21188 29172 21244
rect 29108 21184 29172 21188
rect 29188 21244 29252 21248
rect 29188 21188 29192 21244
rect 29192 21188 29248 21244
rect 29248 21188 29252 21244
rect 29188 21184 29252 21188
rect 29268 21244 29332 21248
rect 29268 21188 29272 21244
rect 29272 21188 29328 21244
rect 29328 21188 29332 21244
rect 29268 21184 29332 21188
rect 24532 20844 24596 20908
rect 14780 20768 14844 20772
rect 14780 20712 14794 20768
rect 14794 20712 14844 20768
rect 14780 20708 14844 20712
rect 16436 20708 16500 20772
rect 6288 20700 6352 20704
rect 6288 20644 6292 20700
rect 6292 20644 6348 20700
rect 6348 20644 6352 20700
rect 6288 20640 6352 20644
rect 6368 20700 6432 20704
rect 6368 20644 6372 20700
rect 6372 20644 6428 20700
rect 6428 20644 6432 20700
rect 6368 20640 6432 20644
rect 6448 20700 6512 20704
rect 6448 20644 6452 20700
rect 6452 20644 6508 20700
rect 6508 20644 6512 20700
rect 6448 20640 6512 20644
rect 6528 20700 6592 20704
rect 6528 20644 6532 20700
rect 6532 20644 6588 20700
rect 6588 20644 6592 20700
rect 6528 20640 6592 20644
rect 13648 20700 13712 20704
rect 13648 20644 13652 20700
rect 13652 20644 13708 20700
rect 13708 20644 13712 20700
rect 13648 20640 13712 20644
rect 13728 20700 13792 20704
rect 13728 20644 13732 20700
rect 13732 20644 13788 20700
rect 13788 20644 13792 20700
rect 13728 20640 13792 20644
rect 13808 20700 13872 20704
rect 13808 20644 13812 20700
rect 13812 20644 13868 20700
rect 13868 20644 13872 20700
rect 13808 20640 13872 20644
rect 13888 20700 13952 20704
rect 13888 20644 13892 20700
rect 13892 20644 13948 20700
rect 13948 20644 13952 20700
rect 13888 20640 13952 20644
rect 21008 20700 21072 20704
rect 21008 20644 21012 20700
rect 21012 20644 21068 20700
rect 21068 20644 21072 20700
rect 21008 20640 21072 20644
rect 21088 20700 21152 20704
rect 21088 20644 21092 20700
rect 21092 20644 21148 20700
rect 21148 20644 21152 20700
rect 21088 20640 21152 20644
rect 21168 20700 21232 20704
rect 21168 20644 21172 20700
rect 21172 20644 21228 20700
rect 21228 20644 21232 20700
rect 21168 20640 21232 20644
rect 21248 20700 21312 20704
rect 21248 20644 21252 20700
rect 21252 20644 21308 20700
rect 21308 20644 21312 20700
rect 21248 20640 21312 20644
rect 28368 20700 28432 20704
rect 28368 20644 28372 20700
rect 28372 20644 28428 20700
rect 28428 20644 28432 20700
rect 28368 20640 28432 20644
rect 28448 20700 28512 20704
rect 28448 20644 28452 20700
rect 28452 20644 28508 20700
rect 28508 20644 28512 20700
rect 28448 20640 28512 20644
rect 28528 20700 28592 20704
rect 28528 20644 28532 20700
rect 28532 20644 28588 20700
rect 28588 20644 28592 20700
rect 28528 20640 28592 20644
rect 28608 20700 28672 20704
rect 28608 20644 28612 20700
rect 28612 20644 28668 20700
rect 28668 20644 28672 20700
rect 28608 20640 28672 20644
rect 11284 20436 11348 20500
rect 6948 20156 7012 20160
rect 6948 20100 6952 20156
rect 6952 20100 7008 20156
rect 7008 20100 7012 20156
rect 6948 20096 7012 20100
rect 7028 20156 7092 20160
rect 7028 20100 7032 20156
rect 7032 20100 7088 20156
rect 7088 20100 7092 20156
rect 7028 20096 7092 20100
rect 7108 20156 7172 20160
rect 7108 20100 7112 20156
rect 7112 20100 7168 20156
rect 7168 20100 7172 20156
rect 7108 20096 7172 20100
rect 7188 20156 7252 20160
rect 7188 20100 7192 20156
rect 7192 20100 7248 20156
rect 7248 20100 7252 20156
rect 7188 20096 7252 20100
rect 14308 20156 14372 20160
rect 14308 20100 14312 20156
rect 14312 20100 14368 20156
rect 14368 20100 14372 20156
rect 14308 20096 14372 20100
rect 14388 20156 14452 20160
rect 14388 20100 14392 20156
rect 14392 20100 14448 20156
rect 14448 20100 14452 20156
rect 14388 20096 14452 20100
rect 14468 20156 14532 20160
rect 14468 20100 14472 20156
rect 14472 20100 14528 20156
rect 14528 20100 14532 20156
rect 14468 20096 14532 20100
rect 14548 20156 14612 20160
rect 14548 20100 14552 20156
rect 14552 20100 14608 20156
rect 14608 20100 14612 20156
rect 14548 20096 14612 20100
rect 21668 20156 21732 20160
rect 21668 20100 21672 20156
rect 21672 20100 21728 20156
rect 21728 20100 21732 20156
rect 21668 20096 21732 20100
rect 21748 20156 21812 20160
rect 21748 20100 21752 20156
rect 21752 20100 21808 20156
rect 21808 20100 21812 20156
rect 21748 20096 21812 20100
rect 21828 20156 21892 20160
rect 21828 20100 21832 20156
rect 21832 20100 21888 20156
rect 21888 20100 21892 20156
rect 21828 20096 21892 20100
rect 21908 20156 21972 20160
rect 21908 20100 21912 20156
rect 21912 20100 21968 20156
rect 21968 20100 21972 20156
rect 21908 20096 21972 20100
rect 29028 20156 29092 20160
rect 29028 20100 29032 20156
rect 29032 20100 29088 20156
rect 29088 20100 29092 20156
rect 29028 20096 29092 20100
rect 29108 20156 29172 20160
rect 29108 20100 29112 20156
rect 29112 20100 29168 20156
rect 29168 20100 29172 20156
rect 29108 20096 29172 20100
rect 29188 20156 29252 20160
rect 29188 20100 29192 20156
rect 29192 20100 29248 20156
rect 29248 20100 29252 20156
rect 29188 20096 29252 20100
rect 29268 20156 29332 20160
rect 29268 20100 29272 20156
rect 29272 20100 29328 20156
rect 29328 20100 29332 20156
rect 29268 20096 29332 20100
rect 15332 19892 15396 19956
rect 6288 19612 6352 19616
rect 6288 19556 6292 19612
rect 6292 19556 6348 19612
rect 6348 19556 6352 19612
rect 6288 19552 6352 19556
rect 6368 19612 6432 19616
rect 6368 19556 6372 19612
rect 6372 19556 6428 19612
rect 6428 19556 6432 19612
rect 6368 19552 6432 19556
rect 6448 19612 6512 19616
rect 6448 19556 6452 19612
rect 6452 19556 6508 19612
rect 6508 19556 6512 19612
rect 6448 19552 6512 19556
rect 6528 19612 6592 19616
rect 6528 19556 6532 19612
rect 6532 19556 6588 19612
rect 6588 19556 6592 19612
rect 6528 19552 6592 19556
rect 13648 19612 13712 19616
rect 13648 19556 13652 19612
rect 13652 19556 13708 19612
rect 13708 19556 13712 19612
rect 13648 19552 13712 19556
rect 13728 19612 13792 19616
rect 13728 19556 13732 19612
rect 13732 19556 13788 19612
rect 13788 19556 13792 19612
rect 13728 19552 13792 19556
rect 13808 19612 13872 19616
rect 13808 19556 13812 19612
rect 13812 19556 13868 19612
rect 13868 19556 13872 19612
rect 13808 19552 13872 19556
rect 13888 19612 13952 19616
rect 13888 19556 13892 19612
rect 13892 19556 13948 19612
rect 13948 19556 13952 19612
rect 13888 19552 13952 19556
rect 21008 19612 21072 19616
rect 21008 19556 21012 19612
rect 21012 19556 21068 19612
rect 21068 19556 21072 19612
rect 21008 19552 21072 19556
rect 21088 19612 21152 19616
rect 21088 19556 21092 19612
rect 21092 19556 21148 19612
rect 21148 19556 21152 19612
rect 21088 19552 21152 19556
rect 21168 19612 21232 19616
rect 21168 19556 21172 19612
rect 21172 19556 21228 19612
rect 21228 19556 21232 19612
rect 21168 19552 21232 19556
rect 21248 19612 21312 19616
rect 21248 19556 21252 19612
rect 21252 19556 21308 19612
rect 21308 19556 21312 19612
rect 21248 19552 21312 19556
rect 28368 19612 28432 19616
rect 28368 19556 28372 19612
rect 28372 19556 28428 19612
rect 28428 19556 28432 19612
rect 28368 19552 28432 19556
rect 28448 19612 28512 19616
rect 28448 19556 28452 19612
rect 28452 19556 28508 19612
rect 28508 19556 28512 19612
rect 28448 19552 28512 19556
rect 28528 19612 28592 19616
rect 28528 19556 28532 19612
rect 28532 19556 28588 19612
rect 28588 19556 28592 19612
rect 28528 19552 28592 19556
rect 28608 19612 28672 19616
rect 28608 19556 28612 19612
rect 28612 19556 28668 19612
rect 28668 19556 28672 19612
rect 28608 19552 28672 19556
rect 12940 19348 13004 19412
rect 12204 19212 12268 19276
rect 6948 19068 7012 19072
rect 6948 19012 6952 19068
rect 6952 19012 7008 19068
rect 7008 19012 7012 19068
rect 6948 19008 7012 19012
rect 7028 19068 7092 19072
rect 7028 19012 7032 19068
rect 7032 19012 7088 19068
rect 7088 19012 7092 19068
rect 7028 19008 7092 19012
rect 7108 19068 7172 19072
rect 7108 19012 7112 19068
rect 7112 19012 7168 19068
rect 7168 19012 7172 19068
rect 7108 19008 7172 19012
rect 7188 19068 7252 19072
rect 7188 19012 7192 19068
rect 7192 19012 7248 19068
rect 7248 19012 7252 19068
rect 7188 19008 7252 19012
rect 14308 19068 14372 19072
rect 14308 19012 14312 19068
rect 14312 19012 14368 19068
rect 14368 19012 14372 19068
rect 14308 19008 14372 19012
rect 14388 19068 14452 19072
rect 14388 19012 14392 19068
rect 14392 19012 14448 19068
rect 14448 19012 14452 19068
rect 14388 19008 14452 19012
rect 14468 19068 14532 19072
rect 14468 19012 14472 19068
rect 14472 19012 14528 19068
rect 14528 19012 14532 19068
rect 14468 19008 14532 19012
rect 14548 19068 14612 19072
rect 14548 19012 14552 19068
rect 14552 19012 14608 19068
rect 14608 19012 14612 19068
rect 14548 19008 14612 19012
rect 21668 19068 21732 19072
rect 21668 19012 21672 19068
rect 21672 19012 21728 19068
rect 21728 19012 21732 19068
rect 21668 19008 21732 19012
rect 21748 19068 21812 19072
rect 21748 19012 21752 19068
rect 21752 19012 21808 19068
rect 21808 19012 21812 19068
rect 21748 19008 21812 19012
rect 21828 19068 21892 19072
rect 21828 19012 21832 19068
rect 21832 19012 21888 19068
rect 21888 19012 21892 19068
rect 21828 19008 21892 19012
rect 21908 19068 21972 19072
rect 21908 19012 21912 19068
rect 21912 19012 21968 19068
rect 21968 19012 21972 19068
rect 21908 19008 21972 19012
rect 29028 19068 29092 19072
rect 29028 19012 29032 19068
rect 29032 19012 29088 19068
rect 29088 19012 29092 19068
rect 29028 19008 29092 19012
rect 29108 19068 29172 19072
rect 29108 19012 29112 19068
rect 29112 19012 29168 19068
rect 29168 19012 29172 19068
rect 29108 19008 29172 19012
rect 29188 19068 29252 19072
rect 29188 19012 29192 19068
rect 29192 19012 29248 19068
rect 29248 19012 29252 19068
rect 29188 19008 29252 19012
rect 29268 19068 29332 19072
rect 29268 19012 29272 19068
rect 29272 19012 29328 19068
rect 29328 19012 29332 19068
rect 29268 19008 29332 19012
rect 6288 18524 6352 18528
rect 6288 18468 6292 18524
rect 6292 18468 6348 18524
rect 6348 18468 6352 18524
rect 6288 18464 6352 18468
rect 6368 18524 6432 18528
rect 6368 18468 6372 18524
rect 6372 18468 6428 18524
rect 6428 18468 6432 18524
rect 6368 18464 6432 18468
rect 6448 18524 6512 18528
rect 6448 18468 6452 18524
rect 6452 18468 6508 18524
rect 6508 18468 6512 18524
rect 6448 18464 6512 18468
rect 6528 18524 6592 18528
rect 6528 18468 6532 18524
rect 6532 18468 6588 18524
rect 6588 18468 6592 18524
rect 6528 18464 6592 18468
rect 13648 18524 13712 18528
rect 13648 18468 13652 18524
rect 13652 18468 13708 18524
rect 13708 18468 13712 18524
rect 13648 18464 13712 18468
rect 13728 18524 13792 18528
rect 13728 18468 13732 18524
rect 13732 18468 13788 18524
rect 13788 18468 13792 18524
rect 13728 18464 13792 18468
rect 13808 18524 13872 18528
rect 13808 18468 13812 18524
rect 13812 18468 13868 18524
rect 13868 18468 13872 18524
rect 13808 18464 13872 18468
rect 13888 18524 13952 18528
rect 13888 18468 13892 18524
rect 13892 18468 13948 18524
rect 13948 18468 13952 18524
rect 13888 18464 13952 18468
rect 21008 18524 21072 18528
rect 21008 18468 21012 18524
rect 21012 18468 21068 18524
rect 21068 18468 21072 18524
rect 21008 18464 21072 18468
rect 21088 18524 21152 18528
rect 21088 18468 21092 18524
rect 21092 18468 21148 18524
rect 21148 18468 21152 18524
rect 21088 18464 21152 18468
rect 21168 18524 21232 18528
rect 21168 18468 21172 18524
rect 21172 18468 21228 18524
rect 21228 18468 21232 18524
rect 21168 18464 21232 18468
rect 21248 18524 21312 18528
rect 21248 18468 21252 18524
rect 21252 18468 21308 18524
rect 21308 18468 21312 18524
rect 21248 18464 21312 18468
rect 28368 18524 28432 18528
rect 28368 18468 28372 18524
rect 28372 18468 28428 18524
rect 28428 18468 28432 18524
rect 28368 18464 28432 18468
rect 28448 18524 28512 18528
rect 28448 18468 28452 18524
rect 28452 18468 28508 18524
rect 28508 18468 28512 18524
rect 28448 18464 28512 18468
rect 28528 18524 28592 18528
rect 28528 18468 28532 18524
rect 28532 18468 28588 18524
rect 28588 18468 28592 18524
rect 28528 18464 28592 18468
rect 28608 18524 28672 18528
rect 28608 18468 28612 18524
rect 28612 18468 28668 18524
rect 28668 18468 28672 18524
rect 28608 18464 28672 18468
rect 6948 17980 7012 17984
rect 6948 17924 6952 17980
rect 6952 17924 7008 17980
rect 7008 17924 7012 17980
rect 6948 17920 7012 17924
rect 7028 17980 7092 17984
rect 7028 17924 7032 17980
rect 7032 17924 7088 17980
rect 7088 17924 7092 17980
rect 7028 17920 7092 17924
rect 7108 17980 7172 17984
rect 7108 17924 7112 17980
rect 7112 17924 7168 17980
rect 7168 17924 7172 17980
rect 7108 17920 7172 17924
rect 7188 17980 7252 17984
rect 7188 17924 7192 17980
rect 7192 17924 7248 17980
rect 7248 17924 7252 17980
rect 7188 17920 7252 17924
rect 14308 17980 14372 17984
rect 14308 17924 14312 17980
rect 14312 17924 14368 17980
rect 14368 17924 14372 17980
rect 14308 17920 14372 17924
rect 14388 17980 14452 17984
rect 14388 17924 14392 17980
rect 14392 17924 14448 17980
rect 14448 17924 14452 17980
rect 14388 17920 14452 17924
rect 14468 17980 14532 17984
rect 14468 17924 14472 17980
rect 14472 17924 14528 17980
rect 14528 17924 14532 17980
rect 14468 17920 14532 17924
rect 14548 17980 14612 17984
rect 14548 17924 14552 17980
rect 14552 17924 14608 17980
rect 14608 17924 14612 17980
rect 14548 17920 14612 17924
rect 21668 17980 21732 17984
rect 21668 17924 21672 17980
rect 21672 17924 21728 17980
rect 21728 17924 21732 17980
rect 21668 17920 21732 17924
rect 21748 17980 21812 17984
rect 21748 17924 21752 17980
rect 21752 17924 21808 17980
rect 21808 17924 21812 17980
rect 21748 17920 21812 17924
rect 21828 17980 21892 17984
rect 21828 17924 21832 17980
rect 21832 17924 21888 17980
rect 21888 17924 21892 17980
rect 21828 17920 21892 17924
rect 21908 17980 21972 17984
rect 21908 17924 21912 17980
rect 21912 17924 21968 17980
rect 21968 17924 21972 17980
rect 21908 17920 21972 17924
rect 29028 17980 29092 17984
rect 29028 17924 29032 17980
rect 29032 17924 29088 17980
rect 29088 17924 29092 17980
rect 29028 17920 29092 17924
rect 29108 17980 29172 17984
rect 29108 17924 29112 17980
rect 29112 17924 29168 17980
rect 29168 17924 29172 17980
rect 29108 17920 29172 17924
rect 29188 17980 29252 17984
rect 29188 17924 29192 17980
rect 29192 17924 29248 17980
rect 29248 17924 29252 17980
rect 29188 17920 29252 17924
rect 29268 17980 29332 17984
rect 29268 17924 29272 17980
rect 29272 17924 29328 17980
rect 29328 17924 29332 17980
rect 29268 17920 29332 17924
rect 6288 17436 6352 17440
rect 6288 17380 6292 17436
rect 6292 17380 6348 17436
rect 6348 17380 6352 17436
rect 6288 17376 6352 17380
rect 6368 17436 6432 17440
rect 6368 17380 6372 17436
rect 6372 17380 6428 17436
rect 6428 17380 6432 17436
rect 6368 17376 6432 17380
rect 6448 17436 6512 17440
rect 6448 17380 6452 17436
rect 6452 17380 6508 17436
rect 6508 17380 6512 17436
rect 6448 17376 6512 17380
rect 6528 17436 6592 17440
rect 6528 17380 6532 17436
rect 6532 17380 6588 17436
rect 6588 17380 6592 17436
rect 6528 17376 6592 17380
rect 13648 17436 13712 17440
rect 13648 17380 13652 17436
rect 13652 17380 13708 17436
rect 13708 17380 13712 17436
rect 13648 17376 13712 17380
rect 13728 17436 13792 17440
rect 13728 17380 13732 17436
rect 13732 17380 13788 17436
rect 13788 17380 13792 17436
rect 13728 17376 13792 17380
rect 13808 17436 13872 17440
rect 13808 17380 13812 17436
rect 13812 17380 13868 17436
rect 13868 17380 13872 17436
rect 13808 17376 13872 17380
rect 13888 17436 13952 17440
rect 13888 17380 13892 17436
rect 13892 17380 13948 17436
rect 13948 17380 13952 17436
rect 13888 17376 13952 17380
rect 21008 17436 21072 17440
rect 21008 17380 21012 17436
rect 21012 17380 21068 17436
rect 21068 17380 21072 17436
rect 21008 17376 21072 17380
rect 21088 17436 21152 17440
rect 21088 17380 21092 17436
rect 21092 17380 21148 17436
rect 21148 17380 21152 17436
rect 21088 17376 21152 17380
rect 21168 17436 21232 17440
rect 21168 17380 21172 17436
rect 21172 17380 21228 17436
rect 21228 17380 21232 17436
rect 21168 17376 21232 17380
rect 21248 17436 21312 17440
rect 21248 17380 21252 17436
rect 21252 17380 21308 17436
rect 21308 17380 21312 17436
rect 21248 17376 21312 17380
rect 28368 17436 28432 17440
rect 28368 17380 28372 17436
rect 28372 17380 28428 17436
rect 28428 17380 28432 17436
rect 28368 17376 28432 17380
rect 28448 17436 28512 17440
rect 28448 17380 28452 17436
rect 28452 17380 28508 17436
rect 28508 17380 28512 17436
rect 28448 17376 28512 17380
rect 28528 17436 28592 17440
rect 28528 17380 28532 17436
rect 28532 17380 28588 17436
rect 28588 17380 28592 17436
rect 28528 17376 28592 17380
rect 28608 17436 28672 17440
rect 28608 17380 28612 17436
rect 28612 17380 28668 17436
rect 28668 17380 28672 17436
rect 28608 17376 28672 17380
rect 6948 16892 7012 16896
rect 6948 16836 6952 16892
rect 6952 16836 7008 16892
rect 7008 16836 7012 16892
rect 6948 16832 7012 16836
rect 7028 16892 7092 16896
rect 7028 16836 7032 16892
rect 7032 16836 7088 16892
rect 7088 16836 7092 16892
rect 7028 16832 7092 16836
rect 7108 16892 7172 16896
rect 7108 16836 7112 16892
rect 7112 16836 7168 16892
rect 7168 16836 7172 16892
rect 7108 16832 7172 16836
rect 7188 16892 7252 16896
rect 7188 16836 7192 16892
rect 7192 16836 7248 16892
rect 7248 16836 7252 16892
rect 7188 16832 7252 16836
rect 14308 16892 14372 16896
rect 14308 16836 14312 16892
rect 14312 16836 14368 16892
rect 14368 16836 14372 16892
rect 14308 16832 14372 16836
rect 14388 16892 14452 16896
rect 14388 16836 14392 16892
rect 14392 16836 14448 16892
rect 14448 16836 14452 16892
rect 14388 16832 14452 16836
rect 14468 16892 14532 16896
rect 14468 16836 14472 16892
rect 14472 16836 14528 16892
rect 14528 16836 14532 16892
rect 14468 16832 14532 16836
rect 14548 16892 14612 16896
rect 14548 16836 14552 16892
rect 14552 16836 14608 16892
rect 14608 16836 14612 16892
rect 14548 16832 14612 16836
rect 21668 16892 21732 16896
rect 21668 16836 21672 16892
rect 21672 16836 21728 16892
rect 21728 16836 21732 16892
rect 21668 16832 21732 16836
rect 21748 16892 21812 16896
rect 21748 16836 21752 16892
rect 21752 16836 21808 16892
rect 21808 16836 21812 16892
rect 21748 16832 21812 16836
rect 21828 16892 21892 16896
rect 21828 16836 21832 16892
rect 21832 16836 21888 16892
rect 21888 16836 21892 16892
rect 21828 16832 21892 16836
rect 21908 16892 21972 16896
rect 21908 16836 21912 16892
rect 21912 16836 21968 16892
rect 21968 16836 21972 16892
rect 21908 16832 21972 16836
rect 29028 16892 29092 16896
rect 29028 16836 29032 16892
rect 29032 16836 29088 16892
rect 29088 16836 29092 16892
rect 29028 16832 29092 16836
rect 29108 16892 29172 16896
rect 29108 16836 29112 16892
rect 29112 16836 29168 16892
rect 29168 16836 29172 16892
rect 29108 16832 29172 16836
rect 29188 16892 29252 16896
rect 29188 16836 29192 16892
rect 29192 16836 29248 16892
rect 29248 16836 29252 16892
rect 29188 16832 29252 16836
rect 29268 16892 29332 16896
rect 29268 16836 29272 16892
rect 29272 16836 29328 16892
rect 29328 16836 29332 16892
rect 29268 16832 29332 16836
rect 11100 16492 11164 16556
rect 16620 16492 16684 16556
rect 6288 16348 6352 16352
rect 6288 16292 6292 16348
rect 6292 16292 6348 16348
rect 6348 16292 6352 16348
rect 6288 16288 6352 16292
rect 6368 16348 6432 16352
rect 6368 16292 6372 16348
rect 6372 16292 6428 16348
rect 6428 16292 6432 16348
rect 6368 16288 6432 16292
rect 6448 16348 6512 16352
rect 6448 16292 6452 16348
rect 6452 16292 6508 16348
rect 6508 16292 6512 16348
rect 6448 16288 6512 16292
rect 6528 16348 6592 16352
rect 6528 16292 6532 16348
rect 6532 16292 6588 16348
rect 6588 16292 6592 16348
rect 6528 16288 6592 16292
rect 13648 16348 13712 16352
rect 13648 16292 13652 16348
rect 13652 16292 13708 16348
rect 13708 16292 13712 16348
rect 13648 16288 13712 16292
rect 13728 16348 13792 16352
rect 13728 16292 13732 16348
rect 13732 16292 13788 16348
rect 13788 16292 13792 16348
rect 13728 16288 13792 16292
rect 13808 16348 13872 16352
rect 13808 16292 13812 16348
rect 13812 16292 13868 16348
rect 13868 16292 13872 16348
rect 13808 16288 13872 16292
rect 13888 16348 13952 16352
rect 13888 16292 13892 16348
rect 13892 16292 13948 16348
rect 13948 16292 13952 16348
rect 13888 16288 13952 16292
rect 21008 16348 21072 16352
rect 21008 16292 21012 16348
rect 21012 16292 21068 16348
rect 21068 16292 21072 16348
rect 21008 16288 21072 16292
rect 21088 16348 21152 16352
rect 21088 16292 21092 16348
rect 21092 16292 21148 16348
rect 21148 16292 21152 16348
rect 21088 16288 21152 16292
rect 21168 16348 21232 16352
rect 21168 16292 21172 16348
rect 21172 16292 21228 16348
rect 21228 16292 21232 16348
rect 21168 16288 21232 16292
rect 21248 16348 21312 16352
rect 21248 16292 21252 16348
rect 21252 16292 21308 16348
rect 21308 16292 21312 16348
rect 21248 16288 21312 16292
rect 28368 16348 28432 16352
rect 28368 16292 28372 16348
rect 28372 16292 28428 16348
rect 28428 16292 28432 16348
rect 28368 16288 28432 16292
rect 28448 16348 28512 16352
rect 28448 16292 28452 16348
rect 28452 16292 28508 16348
rect 28508 16292 28512 16348
rect 28448 16288 28512 16292
rect 28528 16348 28592 16352
rect 28528 16292 28532 16348
rect 28532 16292 28588 16348
rect 28588 16292 28592 16348
rect 28528 16288 28592 16292
rect 28608 16348 28672 16352
rect 28608 16292 28612 16348
rect 28612 16292 28668 16348
rect 28668 16292 28672 16348
rect 28608 16288 28672 16292
rect 6948 15804 7012 15808
rect 6948 15748 6952 15804
rect 6952 15748 7008 15804
rect 7008 15748 7012 15804
rect 6948 15744 7012 15748
rect 7028 15804 7092 15808
rect 7028 15748 7032 15804
rect 7032 15748 7088 15804
rect 7088 15748 7092 15804
rect 7028 15744 7092 15748
rect 7108 15804 7172 15808
rect 7108 15748 7112 15804
rect 7112 15748 7168 15804
rect 7168 15748 7172 15804
rect 7108 15744 7172 15748
rect 7188 15804 7252 15808
rect 7188 15748 7192 15804
rect 7192 15748 7248 15804
rect 7248 15748 7252 15804
rect 7188 15744 7252 15748
rect 14308 15804 14372 15808
rect 14308 15748 14312 15804
rect 14312 15748 14368 15804
rect 14368 15748 14372 15804
rect 14308 15744 14372 15748
rect 14388 15804 14452 15808
rect 14388 15748 14392 15804
rect 14392 15748 14448 15804
rect 14448 15748 14452 15804
rect 14388 15744 14452 15748
rect 14468 15804 14532 15808
rect 14468 15748 14472 15804
rect 14472 15748 14528 15804
rect 14528 15748 14532 15804
rect 14468 15744 14532 15748
rect 14548 15804 14612 15808
rect 14548 15748 14552 15804
rect 14552 15748 14608 15804
rect 14608 15748 14612 15804
rect 14548 15744 14612 15748
rect 21668 15804 21732 15808
rect 21668 15748 21672 15804
rect 21672 15748 21728 15804
rect 21728 15748 21732 15804
rect 21668 15744 21732 15748
rect 21748 15804 21812 15808
rect 21748 15748 21752 15804
rect 21752 15748 21808 15804
rect 21808 15748 21812 15804
rect 21748 15744 21812 15748
rect 21828 15804 21892 15808
rect 21828 15748 21832 15804
rect 21832 15748 21888 15804
rect 21888 15748 21892 15804
rect 21828 15744 21892 15748
rect 21908 15804 21972 15808
rect 21908 15748 21912 15804
rect 21912 15748 21968 15804
rect 21968 15748 21972 15804
rect 21908 15744 21972 15748
rect 29028 15804 29092 15808
rect 29028 15748 29032 15804
rect 29032 15748 29088 15804
rect 29088 15748 29092 15804
rect 29028 15744 29092 15748
rect 29108 15804 29172 15808
rect 29108 15748 29112 15804
rect 29112 15748 29168 15804
rect 29168 15748 29172 15804
rect 29108 15744 29172 15748
rect 29188 15804 29252 15808
rect 29188 15748 29192 15804
rect 29192 15748 29248 15804
rect 29248 15748 29252 15804
rect 29188 15744 29252 15748
rect 29268 15804 29332 15808
rect 29268 15748 29272 15804
rect 29272 15748 29328 15804
rect 29328 15748 29332 15804
rect 29268 15744 29332 15748
rect 6288 15260 6352 15264
rect 6288 15204 6292 15260
rect 6292 15204 6348 15260
rect 6348 15204 6352 15260
rect 6288 15200 6352 15204
rect 6368 15260 6432 15264
rect 6368 15204 6372 15260
rect 6372 15204 6428 15260
rect 6428 15204 6432 15260
rect 6368 15200 6432 15204
rect 6448 15260 6512 15264
rect 6448 15204 6452 15260
rect 6452 15204 6508 15260
rect 6508 15204 6512 15260
rect 6448 15200 6512 15204
rect 6528 15260 6592 15264
rect 6528 15204 6532 15260
rect 6532 15204 6588 15260
rect 6588 15204 6592 15260
rect 6528 15200 6592 15204
rect 13648 15260 13712 15264
rect 13648 15204 13652 15260
rect 13652 15204 13708 15260
rect 13708 15204 13712 15260
rect 13648 15200 13712 15204
rect 13728 15260 13792 15264
rect 13728 15204 13732 15260
rect 13732 15204 13788 15260
rect 13788 15204 13792 15260
rect 13728 15200 13792 15204
rect 13808 15260 13872 15264
rect 13808 15204 13812 15260
rect 13812 15204 13868 15260
rect 13868 15204 13872 15260
rect 13808 15200 13872 15204
rect 13888 15260 13952 15264
rect 13888 15204 13892 15260
rect 13892 15204 13948 15260
rect 13948 15204 13952 15260
rect 13888 15200 13952 15204
rect 21008 15260 21072 15264
rect 21008 15204 21012 15260
rect 21012 15204 21068 15260
rect 21068 15204 21072 15260
rect 21008 15200 21072 15204
rect 21088 15260 21152 15264
rect 21088 15204 21092 15260
rect 21092 15204 21148 15260
rect 21148 15204 21152 15260
rect 21088 15200 21152 15204
rect 21168 15260 21232 15264
rect 21168 15204 21172 15260
rect 21172 15204 21228 15260
rect 21228 15204 21232 15260
rect 21168 15200 21232 15204
rect 21248 15260 21312 15264
rect 21248 15204 21252 15260
rect 21252 15204 21308 15260
rect 21308 15204 21312 15260
rect 21248 15200 21312 15204
rect 28368 15260 28432 15264
rect 28368 15204 28372 15260
rect 28372 15204 28428 15260
rect 28428 15204 28432 15260
rect 28368 15200 28432 15204
rect 28448 15260 28512 15264
rect 28448 15204 28452 15260
rect 28452 15204 28508 15260
rect 28508 15204 28512 15260
rect 28448 15200 28512 15204
rect 28528 15260 28592 15264
rect 28528 15204 28532 15260
rect 28532 15204 28588 15260
rect 28588 15204 28592 15260
rect 28528 15200 28592 15204
rect 28608 15260 28672 15264
rect 28608 15204 28612 15260
rect 28612 15204 28668 15260
rect 28668 15204 28672 15260
rect 28608 15200 28672 15204
rect 15332 15192 15396 15196
rect 15332 15136 15382 15192
rect 15382 15136 15396 15192
rect 15332 15132 15396 15136
rect 6948 14716 7012 14720
rect 6948 14660 6952 14716
rect 6952 14660 7008 14716
rect 7008 14660 7012 14716
rect 6948 14656 7012 14660
rect 7028 14716 7092 14720
rect 7028 14660 7032 14716
rect 7032 14660 7088 14716
rect 7088 14660 7092 14716
rect 7028 14656 7092 14660
rect 7108 14716 7172 14720
rect 7108 14660 7112 14716
rect 7112 14660 7168 14716
rect 7168 14660 7172 14716
rect 7108 14656 7172 14660
rect 7188 14716 7252 14720
rect 7188 14660 7192 14716
rect 7192 14660 7248 14716
rect 7248 14660 7252 14716
rect 7188 14656 7252 14660
rect 14308 14716 14372 14720
rect 14308 14660 14312 14716
rect 14312 14660 14368 14716
rect 14368 14660 14372 14716
rect 14308 14656 14372 14660
rect 14388 14716 14452 14720
rect 14388 14660 14392 14716
rect 14392 14660 14448 14716
rect 14448 14660 14452 14716
rect 14388 14656 14452 14660
rect 14468 14716 14532 14720
rect 14468 14660 14472 14716
rect 14472 14660 14528 14716
rect 14528 14660 14532 14716
rect 14468 14656 14532 14660
rect 14548 14716 14612 14720
rect 14548 14660 14552 14716
rect 14552 14660 14608 14716
rect 14608 14660 14612 14716
rect 14548 14656 14612 14660
rect 21668 14716 21732 14720
rect 21668 14660 21672 14716
rect 21672 14660 21728 14716
rect 21728 14660 21732 14716
rect 21668 14656 21732 14660
rect 21748 14716 21812 14720
rect 21748 14660 21752 14716
rect 21752 14660 21808 14716
rect 21808 14660 21812 14716
rect 21748 14656 21812 14660
rect 21828 14716 21892 14720
rect 21828 14660 21832 14716
rect 21832 14660 21888 14716
rect 21888 14660 21892 14716
rect 21828 14656 21892 14660
rect 21908 14716 21972 14720
rect 21908 14660 21912 14716
rect 21912 14660 21968 14716
rect 21968 14660 21972 14716
rect 21908 14656 21972 14660
rect 29028 14716 29092 14720
rect 29028 14660 29032 14716
rect 29032 14660 29088 14716
rect 29088 14660 29092 14716
rect 29028 14656 29092 14660
rect 29108 14716 29172 14720
rect 29108 14660 29112 14716
rect 29112 14660 29168 14716
rect 29168 14660 29172 14716
rect 29108 14656 29172 14660
rect 29188 14716 29252 14720
rect 29188 14660 29192 14716
rect 29192 14660 29248 14716
rect 29248 14660 29252 14716
rect 29188 14656 29252 14660
rect 29268 14716 29332 14720
rect 29268 14660 29272 14716
rect 29272 14660 29328 14716
rect 29328 14660 29332 14716
rect 29268 14656 29332 14660
rect 12204 14240 12268 14244
rect 12204 14184 12254 14240
rect 12254 14184 12268 14240
rect 12204 14180 12268 14184
rect 6288 14172 6352 14176
rect 6288 14116 6292 14172
rect 6292 14116 6348 14172
rect 6348 14116 6352 14172
rect 6288 14112 6352 14116
rect 6368 14172 6432 14176
rect 6368 14116 6372 14172
rect 6372 14116 6428 14172
rect 6428 14116 6432 14172
rect 6368 14112 6432 14116
rect 6448 14172 6512 14176
rect 6448 14116 6452 14172
rect 6452 14116 6508 14172
rect 6508 14116 6512 14172
rect 6448 14112 6512 14116
rect 6528 14172 6592 14176
rect 6528 14116 6532 14172
rect 6532 14116 6588 14172
rect 6588 14116 6592 14172
rect 6528 14112 6592 14116
rect 13648 14172 13712 14176
rect 13648 14116 13652 14172
rect 13652 14116 13708 14172
rect 13708 14116 13712 14172
rect 13648 14112 13712 14116
rect 13728 14172 13792 14176
rect 13728 14116 13732 14172
rect 13732 14116 13788 14172
rect 13788 14116 13792 14172
rect 13728 14112 13792 14116
rect 13808 14172 13872 14176
rect 13808 14116 13812 14172
rect 13812 14116 13868 14172
rect 13868 14116 13872 14172
rect 13808 14112 13872 14116
rect 13888 14172 13952 14176
rect 13888 14116 13892 14172
rect 13892 14116 13948 14172
rect 13948 14116 13952 14172
rect 13888 14112 13952 14116
rect 21008 14172 21072 14176
rect 21008 14116 21012 14172
rect 21012 14116 21068 14172
rect 21068 14116 21072 14172
rect 21008 14112 21072 14116
rect 21088 14172 21152 14176
rect 21088 14116 21092 14172
rect 21092 14116 21148 14172
rect 21148 14116 21152 14172
rect 21088 14112 21152 14116
rect 21168 14172 21232 14176
rect 21168 14116 21172 14172
rect 21172 14116 21228 14172
rect 21228 14116 21232 14172
rect 21168 14112 21232 14116
rect 21248 14172 21312 14176
rect 21248 14116 21252 14172
rect 21252 14116 21308 14172
rect 21308 14116 21312 14172
rect 21248 14112 21312 14116
rect 28368 14172 28432 14176
rect 28368 14116 28372 14172
rect 28372 14116 28428 14172
rect 28428 14116 28432 14172
rect 28368 14112 28432 14116
rect 28448 14172 28512 14176
rect 28448 14116 28452 14172
rect 28452 14116 28508 14172
rect 28508 14116 28512 14172
rect 28448 14112 28512 14116
rect 28528 14172 28592 14176
rect 28528 14116 28532 14172
rect 28532 14116 28588 14172
rect 28588 14116 28592 14172
rect 28528 14112 28592 14116
rect 28608 14172 28672 14176
rect 28608 14116 28612 14172
rect 28612 14116 28668 14172
rect 28668 14116 28672 14172
rect 28608 14112 28672 14116
rect 16436 13636 16500 13700
rect 6948 13628 7012 13632
rect 6948 13572 6952 13628
rect 6952 13572 7008 13628
rect 7008 13572 7012 13628
rect 6948 13568 7012 13572
rect 7028 13628 7092 13632
rect 7028 13572 7032 13628
rect 7032 13572 7088 13628
rect 7088 13572 7092 13628
rect 7028 13568 7092 13572
rect 7108 13628 7172 13632
rect 7108 13572 7112 13628
rect 7112 13572 7168 13628
rect 7168 13572 7172 13628
rect 7108 13568 7172 13572
rect 7188 13628 7252 13632
rect 7188 13572 7192 13628
rect 7192 13572 7248 13628
rect 7248 13572 7252 13628
rect 7188 13568 7252 13572
rect 14308 13628 14372 13632
rect 14308 13572 14312 13628
rect 14312 13572 14368 13628
rect 14368 13572 14372 13628
rect 14308 13568 14372 13572
rect 14388 13628 14452 13632
rect 14388 13572 14392 13628
rect 14392 13572 14448 13628
rect 14448 13572 14452 13628
rect 14388 13568 14452 13572
rect 14468 13628 14532 13632
rect 14468 13572 14472 13628
rect 14472 13572 14528 13628
rect 14528 13572 14532 13628
rect 14468 13568 14532 13572
rect 14548 13628 14612 13632
rect 14548 13572 14552 13628
rect 14552 13572 14608 13628
rect 14608 13572 14612 13628
rect 14548 13568 14612 13572
rect 21668 13628 21732 13632
rect 21668 13572 21672 13628
rect 21672 13572 21728 13628
rect 21728 13572 21732 13628
rect 21668 13568 21732 13572
rect 21748 13628 21812 13632
rect 21748 13572 21752 13628
rect 21752 13572 21808 13628
rect 21808 13572 21812 13628
rect 21748 13568 21812 13572
rect 21828 13628 21892 13632
rect 21828 13572 21832 13628
rect 21832 13572 21888 13628
rect 21888 13572 21892 13628
rect 21828 13568 21892 13572
rect 21908 13628 21972 13632
rect 21908 13572 21912 13628
rect 21912 13572 21968 13628
rect 21968 13572 21972 13628
rect 21908 13568 21972 13572
rect 29028 13628 29092 13632
rect 29028 13572 29032 13628
rect 29032 13572 29088 13628
rect 29088 13572 29092 13628
rect 29028 13568 29092 13572
rect 29108 13628 29172 13632
rect 29108 13572 29112 13628
rect 29112 13572 29168 13628
rect 29168 13572 29172 13628
rect 29108 13568 29172 13572
rect 29188 13628 29252 13632
rect 29188 13572 29192 13628
rect 29192 13572 29248 13628
rect 29248 13572 29252 13628
rect 29188 13568 29252 13572
rect 29268 13628 29332 13632
rect 29268 13572 29272 13628
rect 29272 13572 29328 13628
rect 29328 13572 29332 13628
rect 29268 13568 29332 13572
rect 6288 13084 6352 13088
rect 6288 13028 6292 13084
rect 6292 13028 6348 13084
rect 6348 13028 6352 13084
rect 6288 13024 6352 13028
rect 6368 13084 6432 13088
rect 6368 13028 6372 13084
rect 6372 13028 6428 13084
rect 6428 13028 6432 13084
rect 6368 13024 6432 13028
rect 6448 13084 6512 13088
rect 6448 13028 6452 13084
rect 6452 13028 6508 13084
rect 6508 13028 6512 13084
rect 6448 13024 6512 13028
rect 6528 13084 6592 13088
rect 6528 13028 6532 13084
rect 6532 13028 6588 13084
rect 6588 13028 6592 13084
rect 6528 13024 6592 13028
rect 13648 13084 13712 13088
rect 13648 13028 13652 13084
rect 13652 13028 13708 13084
rect 13708 13028 13712 13084
rect 13648 13024 13712 13028
rect 13728 13084 13792 13088
rect 13728 13028 13732 13084
rect 13732 13028 13788 13084
rect 13788 13028 13792 13084
rect 13728 13024 13792 13028
rect 13808 13084 13872 13088
rect 13808 13028 13812 13084
rect 13812 13028 13868 13084
rect 13868 13028 13872 13084
rect 13808 13024 13872 13028
rect 13888 13084 13952 13088
rect 13888 13028 13892 13084
rect 13892 13028 13948 13084
rect 13948 13028 13952 13084
rect 13888 13024 13952 13028
rect 21008 13084 21072 13088
rect 21008 13028 21012 13084
rect 21012 13028 21068 13084
rect 21068 13028 21072 13084
rect 21008 13024 21072 13028
rect 21088 13084 21152 13088
rect 21088 13028 21092 13084
rect 21092 13028 21148 13084
rect 21148 13028 21152 13084
rect 21088 13024 21152 13028
rect 21168 13084 21232 13088
rect 21168 13028 21172 13084
rect 21172 13028 21228 13084
rect 21228 13028 21232 13084
rect 21168 13024 21232 13028
rect 21248 13084 21312 13088
rect 21248 13028 21252 13084
rect 21252 13028 21308 13084
rect 21308 13028 21312 13084
rect 21248 13024 21312 13028
rect 28368 13084 28432 13088
rect 28368 13028 28372 13084
rect 28372 13028 28428 13084
rect 28428 13028 28432 13084
rect 28368 13024 28432 13028
rect 28448 13084 28512 13088
rect 28448 13028 28452 13084
rect 28452 13028 28508 13084
rect 28508 13028 28512 13084
rect 28448 13024 28512 13028
rect 28528 13084 28592 13088
rect 28528 13028 28532 13084
rect 28532 13028 28588 13084
rect 28588 13028 28592 13084
rect 28528 13024 28592 13028
rect 28608 13084 28672 13088
rect 28608 13028 28612 13084
rect 28612 13028 28668 13084
rect 28668 13028 28672 13084
rect 28608 13024 28672 13028
rect 6948 12540 7012 12544
rect 6948 12484 6952 12540
rect 6952 12484 7008 12540
rect 7008 12484 7012 12540
rect 6948 12480 7012 12484
rect 7028 12540 7092 12544
rect 7028 12484 7032 12540
rect 7032 12484 7088 12540
rect 7088 12484 7092 12540
rect 7028 12480 7092 12484
rect 7108 12540 7172 12544
rect 7108 12484 7112 12540
rect 7112 12484 7168 12540
rect 7168 12484 7172 12540
rect 7108 12480 7172 12484
rect 7188 12540 7252 12544
rect 7188 12484 7192 12540
rect 7192 12484 7248 12540
rect 7248 12484 7252 12540
rect 7188 12480 7252 12484
rect 14308 12540 14372 12544
rect 14308 12484 14312 12540
rect 14312 12484 14368 12540
rect 14368 12484 14372 12540
rect 14308 12480 14372 12484
rect 14388 12540 14452 12544
rect 14388 12484 14392 12540
rect 14392 12484 14448 12540
rect 14448 12484 14452 12540
rect 14388 12480 14452 12484
rect 14468 12540 14532 12544
rect 14468 12484 14472 12540
rect 14472 12484 14528 12540
rect 14528 12484 14532 12540
rect 14468 12480 14532 12484
rect 14548 12540 14612 12544
rect 14548 12484 14552 12540
rect 14552 12484 14608 12540
rect 14608 12484 14612 12540
rect 14548 12480 14612 12484
rect 21668 12540 21732 12544
rect 21668 12484 21672 12540
rect 21672 12484 21728 12540
rect 21728 12484 21732 12540
rect 21668 12480 21732 12484
rect 21748 12540 21812 12544
rect 21748 12484 21752 12540
rect 21752 12484 21808 12540
rect 21808 12484 21812 12540
rect 21748 12480 21812 12484
rect 21828 12540 21892 12544
rect 21828 12484 21832 12540
rect 21832 12484 21888 12540
rect 21888 12484 21892 12540
rect 21828 12480 21892 12484
rect 21908 12540 21972 12544
rect 21908 12484 21912 12540
rect 21912 12484 21968 12540
rect 21968 12484 21972 12540
rect 21908 12480 21972 12484
rect 29028 12540 29092 12544
rect 29028 12484 29032 12540
rect 29032 12484 29088 12540
rect 29088 12484 29092 12540
rect 29028 12480 29092 12484
rect 29108 12540 29172 12544
rect 29108 12484 29112 12540
rect 29112 12484 29168 12540
rect 29168 12484 29172 12540
rect 29108 12480 29172 12484
rect 29188 12540 29252 12544
rect 29188 12484 29192 12540
rect 29192 12484 29248 12540
rect 29248 12484 29252 12540
rect 29188 12480 29252 12484
rect 29268 12540 29332 12544
rect 29268 12484 29272 12540
rect 29272 12484 29328 12540
rect 29328 12484 29332 12540
rect 29268 12480 29332 12484
rect 6288 11996 6352 12000
rect 6288 11940 6292 11996
rect 6292 11940 6348 11996
rect 6348 11940 6352 11996
rect 6288 11936 6352 11940
rect 6368 11996 6432 12000
rect 6368 11940 6372 11996
rect 6372 11940 6428 11996
rect 6428 11940 6432 11996
rect 6368 11936 6432 11940
rect 6448 11996 6512 12000
rect 6448 11940 6452 11996
rect 6452 11940 6508 11996
rect 6508 11940 6512 11996
rect 6448 11936 6512 11940
rect 6528 11996 6592 12000
rect 6528 11940 6532 11996
rect 6532 11940 6588 11996
rect 6588 11940 6592 11996
rect 6528 11936 6592 11940
rect 13648 11996 13712 12000
rect 13648 11940 13652 11996
rect 13652 11940 13708 11996
rect 13708 11940 13712 11996
rect 13648 11936 13712 11940
rect 13728 11996 13792 12000
rect 13728 11940 13732 11996
rect 13732 11940 13788 11996
rect 13788 11940 13792 11996
rect 13728 11936 13792 11940
rect 13808 11996 13872 12000
rect 13808 11940 13812 11996
rect 13812 11940 13868 11996
rect 13868 11940 13872 11996
rect 13808 11936 13872 11940
rect 13888 11996 13952 12000
rect 13888 11940 13892 11996
rect 13892 11940 13948 11996
rect 13948 11940 13952 11996
rect 13888 11936 13952 11940
rect 21008 11996 21072 12000
rect 21008 11940 21012 11996
rect 21012 11940 21068 11996
rect 21068 11940 21072 11996
rect 21008 11936 21072 11940
rect 21088 11996 21152 12000
rect 21088 11940 21092 11996
rect 21092 11940 21148 11996
rect 21148 11940 21152 11996
rect 21088 11936 21152 11940
rect 21168 11996 21232 12000
rect 21168 11940 21172 11996
rect 21172 11940 21228 11996
rect 21228 11940 21232 11996
rect 21168 11936 21232 11940
rect 21248 11996 21312 12000
rect 21248 11940 21252 11996
rect 21252 11940 21308 11996
rect 21308 11940 21312 11996
rect 21248 11936 21312 11940
rect 28368 11996 28432 12000
rect 28368 11940 28372 11996
rect 28372 11940 28428 11996
rect 28428 11940 28432 11996
rect 28368 11936 28432 11940
rect 28448 11996 28512 12000
rect 28448 11940 28452 11996
rect 28452 11940 28508 11996
rect 28508 11940 28512 11996
rect 28448 11936 28512 11940
rect 28528 11996 28592 12000
rect 28528 11940 28532 11996
rect 28532 11940 28588 11996
rect 28588 11940 28592 11996
rect 28528 11936 28592 11940
rect 28608 11996 28672 12000
rect 28608 11940 28612 11996
rect 28612 11940 28668 11996
rect 28668 11940 28672 11996
rect 28608 11936 28672 11940
rect 24532 11928 24596 11932
rect 24532 11872 24546 11928
rect 24546 11872 24596 11928
rect 24532 11868 24596 11872
rect 6948 11452 7012 11456
rect 6948 11396 6952 11452
rect 6952 11396 7008 11452
rect 7008 11396 7012 11452
rect 6948 11392 7012 11396
rect 7028 11452 7092 11456
rect 7028 11396 7032 11452
rect 7032 11396 7088 11452
rect 7088 11396 7092 11452
rect 7028 11392 7092 11396
rect 7108 11452 7172 11456
rect 7108 11396 7112 11452
rect 7112 11396 7168 11452
rect 7168 11396 7172 11452
rect 7108 11392 7172 11396
rect 7188 11452 7252 11456
rect 7188 11396 7192 11452
rect 7192 11396 7248 11452
rect 7248 11396 7252 11452
rect 7188 11392 7252 11396
rect 14308 11452 14372 11456
rect 14308 11396 14312 11452
rect 14312 11396 14368 11452
rect 14368 11396 14372 11452
rect 14308 11392 14372 11396
rect 14388 11452 14452 11456
rect 14388 11396 14392 11452
rect 14392 11396 14448 11452
rect 14448 11396 14452 11452
rect 14388 11392 14452 11396
rect 14468 11452 14532 11456
rect 14468 11396 14472 11452
rect 14472 11396 14528 11452
rect 14528 11396 14532 11452
rect 14468 11392 14532 11396
rect 14548 11452 14612 11456
rect 14548 11396 14552 11452
rect 14552 11396 14608 11452
rect 14608 11396 14612 11452
rect 14548 11392 14612 11396
rect 21668 11452 21732 11456
rect 21668 11396 21672 11452
rect 21672 11396 21728 11452
rect 21728 11396 21732 11452
rect 21668 11392 21732 11396
rect 21748 11452 21812 11456
rect 21748 11396 21752 11452
rect 21752 11396 21808 11452
rect 21808 11396 21812 11452
rect 21748 11392 21812 11396
rect 21828 11452 21892 11456
rect 21828 11396 21832 11452
rect 21832 11396 21888 11452
rect 21888 11396 21892 11452
rect 21828 11392 21892 11396
rect 21908 11452 21972 11456
rect 21908 11396 21912 11452
rect 21912 11396 21968 11452
rect 21968 11396 21972 11452
rect 21908 11392 21972 11396
rect 29028 11452 29092 11456
rect 29028 11396 29032 11452
rect 29032 11396 29088 11452
rect 29088 11396 29092 11452
rect 29028 11392 29092 11396
rect 29108 11452 29172 11456
rect 29108 11396 29112 11452
rect 29112 11396 29168 11452
rect 29168 11396 29172 11452
rect 29108 11392 29172 11396
rect 29188 11452 29252 11456
rect 29188 11396 29192 11452
rect 29192 11396 29248 11452
rect 29248 11396 29252 11452
rect 29188 11392 29252 11396
rect 29268 11452 29332 11456
rect 29268 11396 29272 11452
rect 29272 11396 29328 11452
rect 29328 11396 29332 11452
rect 29268 11392 29332 11396
rect 14780 11188 14844 11252
rect 6288 10908 6352 10912
rect 6288 10852 6292 10908
rect 6292 10852 6348 10908
rect 6348 10852 6352 10908
rect 6288 10848 6352 10852
rect 6368 10908 6432 10912
rect 6368 10852 6372 10908
rect 6372 10852 6428 10908
rect 6428 10852 6432 10908
rect 6368 10848 6432 10852
rect 6448 10908 6512 10912
rect 6448 10852 6452 10908
rect 6452 10852 6508 10908
rect 6508 10852 6512 10908
rect 6448 10848 6512 10852
rect 6528 10908 6592 10912
rect 6528 10852 6532 10908
rect 6532 10852 6588 10908
rect 6588 10852 6592 10908
rect 6528 10848 6592 10852
rect 13648 10908 13712 10912
rect 13648 10852 13652 10908
rect 13652 10852 13708 10908
rect 13708 10852 13712 10908
rect 13648 10848 13712 10852
rect 13728 10908 13792 10912
rect 13728 10852 13732 10908
rect 13732 10852 13788 10908
rect 13788 10852 13792 10908
rect 13728 10848 13792 10852
rect 13808 10908 13872 10912
rect 13808 10852 13812 10908
rect 13812 10852 13868 10908
rect 13868 10852 13872 10908
rect 13808 10848 13872 10852
rect 13888 10908 13952 10912
rect 13888 10852 13892 10908
rect 13892 10852 13948 10908
rect 13948 10852 13952 10908
rect 13888 10848 13952 10852
rect 21008 10908 21072 10912
rect 21008 10852 21012 10908
rect 21012 10852 21068 10908
rect 21068 10852 21072 10908
rect 21008 10848 21072 10852
rect 21088 10908 21152 10912
rect 21088 10852 21092 10908
rect 21092 10852 21148 10908
rect 21148 10852 21152 10908
rect 21088 10848 21152 10852
rect 21168 10908 21232 10912
rect 21168 10852 21172 10908
rect 21172 10852 21228 10908
rect 21228 10852 21232 10908
rect 21168 10848 21232 10852
rect 21248 10908 21312 10912
rect 21248 10852 21252 10908
rect 21252 10852 21308 10908
rect 21308 10852 21312 10908
rect 21248 10848 21312 10852
rect 28368 10908 28432 10912
rect 28368 10852 28372 10908
rect 28372 10852 28428 10908
rect 28428 10852 28432 10908
rect 28368 10848 28432 10852
rect 28448 10908 28512 10912
rect 28448 10852 28452 10908
rect 28452 10852 28508 10908
rect 28508 10852 28512 10908
rect 28448 10848 28512 10852
rect 28528 10908 28592 10912
rect 28528 10852 28532 10908
rect 28532 10852 28588 10908
rect 28588 10852 28592 10908
rect 28528 10848 28592 10852
rect 28608 10908 28672 10912
rect 28608 10852 28612 10908
rect 28612 10852 28668 10908
rect 28668 10852 28672 10908
rect 28608 10848 28672 10852
rect 6948 10364 7012 10368
rect 6948 10308 6952 10364
rect 6952 10308 7008 10364
rect 7008 10308 7012 10364
rect 6948 10304 7012 10308
rect 7028 10364 7092 10368
rect 7028 10308 7032 10364
rect 7032 10308 7088 10364
rect 7088 10308 7092 10364
rect 7028 10304 7092 10308
rect 7108 10364 7172 10368
rect 7108 10308 7112 10364
rect 7112 10308 7168 10364
rect 7168 10308 7172 10364
rect 7108 10304 7172 10308
rect 7188 10364 7252 10368
rect 7188 10308 7192 10364
rect 7192 10308 7248 10364
rect 7248 10308 7252 10364
rect 7188 10304 7252 10308
rect 14308 10364 14372 10368
rect 14308 10308 14312 10364
rect 14312 10308 14368 10364
rect 14368 10308 14372 10364
rect 14308 10304 14372 10308
rect 14388 10364 14452 10368
rect 14388 10308 14392 10364
rect 14392 10308 14448 10364
rect 14448 10308 14452 10364
rect 14388 10304 14452 10308
rect 14468 10364 14532 10368
rect 14468 10308 14472 10364
rect 14472 10308 14528 10364
rect 14528 10308 14532 10364
rect 14468 10304 14532 10308
rect 14548 10364 14612 10368
rect 14548 10308 14552 10364
rect 14552 10308 14608 10364
rect 14608 10308 14612 10364
rect 14548 10304 14612 10308
rect 21668 10364 21732 10368
rect 21668 10308 21672 10364
rect 21672 10308 21728 10364
rect 21728 10308 21732 10364
rect 21668 10304 21732 10308
rect 21748 10364 21812 10368
rect 21748 10308 21752 10364
rect 21752 10308 21808 10364
rect 21808 10308 21812 10364
rect 21748 10304 21812 10308
rect 21828 10364 21892 10368
rect 21828 10308 21832 10364
rect 21832 10308 21888 10364
rect 21888 10308 21892 10364
rect 21828 10304 21892 10308
rect 21908 10364 21972 10368
rect 21908 10308 21912 10364
rect 21912 10308 21968 10364
rect 21968 10308 21972 10364
rect 21908 10304 21972 10308
rect 29028 10364 29092 10368
rect 29028 10308 29032 10364
rect 29032 10308 29088 10364
rect 29088 10308 29092 10364
rect 29028 10304 29092 10308
rect 29108 10364 29172 10368
rect 29108 10308 29112 10364
rect 29112 10308 29168 10364
rect 29168 10308 29172 10364
rect 29108 10304 29172 10308
rect 29188 10364 29252 10368
rect 29188 10308 29192 10364
rect 29192 10308 29248 10364
rect 29248 10308 29252 10364
rect 29188 10304 29252 10308
rect 29268 10364 29332 10368
rect 29268 10308 29272 10364
rect 29272 10308 29328 10364
rect 29328 10308 29332 10364
rect 29268 10304 29332 10308
rect 6288 9820 6352 9824
rect 6288 9764 6292 9820
rect 6292 9764 6348 9820
rect 6348 9764 6352 9820
rect 6288 9760 6352 9764
rect 6368 9820 6432 9824
rect 6368 9764 6372 9820
rect 6372 9764 6428 9820
rect 6428 9764 6432 9820
rect 6368 9760 6432 9764
rect 6448 9820 6512 9824
rect 6448 9764 6452 9820
rect 6452 9764 6508 9820
rect 6508 9764 6512 9820
rect 6448 9760 6512 9764
rect 6528 9820 6592 9824
rect 6528 9764 6532 9820
rect 6532 9764 6588 9820
rect 6588 9764 6592 9820
rect 6528 9760 6592 9764
rect 13648 9820 13712 9824
rect 13648 9764 13652 9820
rect 13652 9764 13708 9820
rect 13708 9764 13712 9820
rect 13648 9760 13712 9764
rect 13728 9820 13792 9824
rect 13728 9764 13732 9820
rect 13732 9764 13788 9820
rect 13788 9764 13792 9820
rect 13728 9760 13792 9764
rect 13808 9820 13872 9824
rect 13808 9764 13812 9820
rect 13812 9764 13868 9820
rect 13868 9764 13872 9820
rect 13808 9760 13872 9764
rect 13888 9820 13952 9824
rect 13888 9764 13892 9820
rect 13892 9764 13948 9820
rect 13948 9764 13952 9820
rect 13888 9760 13952 9764
rect 21008 9820 21072 9824
rect 21008 9764 21012 9820
rect 21012 9764 21068 9820
rect 21068 9764 21072 9820
rect 21008 9760 21072 9764
rect 21088 9820 21152 9824
rect 21088 9764 21092 9820
rect 21092 9764 21148 9820
rect 21148 9764 21152 9820
rect 21088 9760 21152 9764
rect 21168 9820 21232 9824
rect 21168 9764 21172 9820
rect 21172 9764 21228 9820
rect 21228 9764 21232 9820
rect 21168 9760 21232 9764
rect 21248 9820 21312 9824
rect 21248 9764 21252 9820
rect 21252 9764 21308 9820
rect 21308 9764 21312 9820
rect 21248 9760 21312 9764
rect 28368 9820 28432 9824
rect 28368 9764 28372 9820
rect 28372 9764 28428 9820
rect 28428 9764 28432 9820
rect 28368 9760 28432 9764
rect 28448 9820 28512 9824
rect 28448 9764 28452 9820
rect 28452 9764 28508 9820
rect 28508 9764 28512 9820
rect 28448 9760 28512 9764
rect 28528 9820 28592 9824
rect 28528 9764 28532 9820
rect 28532 9764 28588 9820
rect 28588 9764 28592 9820
rect 28528 9760 28592 9764
rect 28608 9820 28672 9824
rect 28608 9764 28612 9820
rect 28612 9764 28668 9820
rect 28668 9764 28672 9820
rect 28608 9760 28672 9764
rect 6948 9276 7012 9280
rect 6948 9220 6952 9276
rect 6952 9220 7008 9276
rect 7008 9220 7012 9276
rect 6948 9216 7012 9220
rect 7028 9276 7092 9280
rect 7028 9220 7032 9276
rect 7032 9220 7088 9276
rect 7088 9220 7092 9276
rect 7028 9216 7092 9220
rect 7108 9276 7172 9280
rect 7108 9220 7112 9276
rect 7112 9220 7168 9276
rect 7168 9220 7172 9276
rect 7108 9216 7172 9220
rect 7188 9276 7252 9280
rect 7188 9220 7192 9276
rect 7192 9220 7248 9276
rect 7248 9220 7252 9276
rect 7188 9216 7252 9220
rect 14308 9276 14372 9280
rect 14308 9220 14312 9276
rect 14312 9220 14368 9276
rect 14368 9220 14372 9276
rect 14308 9216 14372 9220
rect 14388 9276 14452 9280
rect 14388 9220 14392 9276
rect 14392 9220 14448 9276
rect 14448 9220 14452 9276
rect 14388 9216 14452 9220
rect 14468 9276 14532 9280
rect 14468 9220 14472 9276
rect 14472 9220 14528 9276
rect 14528 9220 14532 9276
rect 14468 9216 14532 9220
rect 14548 9276 14612 9280
rect 14548 9220 14552 9276
rect 14552 9220 14608 9276
rect 14608 9220 14612 9276
rect 14548 9216 14612 9220
rect 21668 9276 21732 9280
rect 21668 9220 21672 9276
rect 21672 9220 21728 9276
rect 21728 9220 21732 9276
rect 21668 9216 21732 9220
rect 21748 9276 21812 9280
rect 21748 9220 21752 9276
rect 21752 9220 21808 9276
rect 21808 9220 21812 9276
rect 21748 9216 21812 9220
rect 21828 9276 21892 9280
rect 21828 9220 21832 9276
rect 21832 9220 21888 9276
rect 21888 9220 21892 9276
rect 21828 9216 21892 9220
rect 21908 9276 21972 9280
rect 21908 9220 21912 9276
rect 21912 9220 21968 9276
rect 21968 9220 21972 9276
rect 21908 9216 21972 9220
rect 29028 9276 29092 9280
rect 29028 9220 29032 9276
rect 29032 9220 29088 9276
rect 29088 9220 29092 9276
rect 29028 9216 29092 9220
rect 29108 9276 29172 9280
rect 29108 9220 29112 9276
rect 29112 9220 29168 9276
rect 29168 9220 29172 9276
rect 29108 9216 29172 9220
rect 29188 9276 29252 9280
rect 29188 9220 29192 9276
rect 29192 9220 29248 9276
rect 29248 9220 29252 9276
rect 29188 9216 29252 9220
rect 29268 9276 29332 9280
rect 29268 9220 29272 9276
rect 29272 9220 29328 9276
rect 29328 9220 29332 9276
rect 29268 9216 29332 9220
rect 6288 8732 6352 8736
rect 6288 8676 6292 8732
rect 6292 8676 6348 8732
rect 6348 8676 6352 8732
rect 6288 8672 6352 8676
rect 6368 8732 6432 8736
rect 6368 8676 6372 8732
rect 6372 8676 6428 8732
rect 6428 8676 6432 8732
rect 6368 8672 6432 8676
rect 6448 8732 6512 8736
rect 6448 8676 6452 8732
rect 6452 8676 6508 8732
rect 6508 8676 6512 8732
rect 6448 8672 6512 8676
rect 6528 8732 6592 8736
rect 6528 8676 6532 8732
rect 6532 8676 6588 8732
rect 6588 8676 6592 8732
rect 6528 8672 6592 8676
rect 13648 8732 13712 8736
rect 13648 8676 13652 8732
rect 13652 8676 13708 8732
rect 13708 8676 13712 8732
rect 13648 8672 13712 8676
rect 13728 8732 13792 8736
rect 13728 8676 13732 8732
rect 13732 8676 13788 8732
rect 13788 8676 13792 8732
rect 13728 8672 13792 8676
rect 13808 8732 13872 8736
rect 13808 8676 13812 8732
rect 13812 8676 13868 8732
rect 13868 8676 13872 8732
rect 13808 8672 13872 8676
rect 13888 8732 13952 8736
rect 13888 8676 13892 8732
rect 13892 8676 13948 8732
rect 13948 8676 13952 8732
rect 13888 8672 13952 8676
rect 21008 8732 21072 8736
rect 21008 8676 21012 8732
rect 21012 8676 21068 8732
rect 21068 8676 21072 8732
rect 21008 8672 21072 8676
rect 21088 8732 21152 8736
rect 21088 8676 21092 8732
rect 21092 8676 21148 8732
rect 21148 8676 21152 8732
rect 21088 8672 21152 8676
rect 21168 8732 21232 8736
rect 21168 8676 21172 8732
rect 21172 8676 21228 8732
rect 21228 8676 21232 8732
rect 21168 8672 21232 8676
rect 21248 8732 21312 8736
rect 21248 8676 21252 8732
rect 21252 8676 21308 8732
rect 21308 8676 21312 8732
rect 21248 8672 21312 8676
rect 28368 8732 28432 8736
rect 28368 8676 28372 8732
rect 28372 8676 28428 8732
rect 28428 8676 28432 8732
rect 28368 8672 28432 8676
rect 28448 8732 28512 8736
rect 28448 8676 28452 8732
rect 28452 8676 28508 8732
rect 28508 8676 28512 8732
rect 28448 8672 28512 8676
rect 28528 8732 28592 8736
rect 28528 8676 28532 8732
rect 28532 8676 28588 8732
rect 28588 8676 28592 8732
rect 28528 8672 28592 8676
rect 28608 8732 28672 8736
rect 28608 8676 28612 8732
rect 28612 8676 28668 8732
rect 28668 8676 28672 8732
rect 28608 8672 28672 8676
rect 13124 8196 13188 8260
rect 6948 8188 7012 8192
rect 6948 8132 6952 8188
rect 6952 8132 7008 8188
rect 7008 8132 7012 8188
rect 6948 8128 7012 8132
rect 7028 8188 7092 8192
rect 7028 8132 7032 8188
rect 7032 8132 7088 8188
rect 7088 8132 7092 8188
rect 7028 8128 7092 8132
rect 7108 8188 7172 8192
rect 7108 8132 7112 8188
rect 7112 8132 7168 8188
rect 7168 8132 7172 8188
rect 7108 8128 7172 8132
rect 7188 8188 7252 8192
rect 7188 8132 7192 8188
rect 7192 8132 7248 8188
rect 7248 8132 7252 8188
rect 7188 8128 7252 8132
rect 14308 8188 14372 8192
rect 14308 8132 14312 8188
rect 14312 8132 14368 8188
rect 14368 8132 14372 8188
rect 14308 8128 14372 8132
rect 14388 8188 14452 8192
rect 14388 8132 14392 8188
rect 14392 8132 14448 8188
rect 14448 8132 14452 8188
rect 14388 8128 14452 8132
rect 14468 8188 14532 8192
rect 14468 8132 14472 8188
rect 14472 8132 14528 8188
rect 14528 8132 14532 8188
rect 14468 8128 14532 8132
rect 14548 8188 14612 8192
rect 14548 8132 14552 8188
rect 14552 8132 14608 8188
rect 14608 8132 14612 8188
rect 14548 8128 14612 8132
rect 21668 8188 21732 8192
rect 21668 8132 21672 8188
rect 21672 8132 21728 8188
rect 21728 8132 21732 8188
rect 21668 8128 21732 8132
rect 21748 8188 21812 8192
rect 21748 8132 21752 8188
rect 21752 8132 21808 8188
rect 21808 8132 21812 8188
rect 21748 8128 21812 8132
rect 21828 8188 21892 8192
rect 21828 8132 21832 8188
rect 21832 8132 21888 8188
rect 21888 8132 21892 8188
rect 21828 8128 21892 8132
rect 21908 8188 21972 8192
rect 21908 8132 21912 8188
rect 21912 8132 21968 8188
rect 21968 8132 21972 8188
rect 21908 8128 21972 8132
rect 29028 8188 29092 8192
rect 29028 8132 29032 8188
rect 29032 8132 29088 8188
rect 29088 8132 29092 8188
rect 29028 8128 29092 8132
rect 29108 8188 29172 8192
rect 29108 8132 29112 8188
rect 29112 8132 29168 8188
rect 29168 8132 29172 8188
rect 29108 8128 29172 8132
rect 29188 8188 29252 8192
rect 29188 8132 29192 8188
rect 29192 8132 29248 8188
rect 29248 8132 29252 8188
rect 29188 8128 29252 8132
rect 29268 8188 29332 8192
rect 29268 8132 29272 8188
rect 29272 8132 29328 8188
rect 29328 8132 29332 8188
rect 29268 8128 29332 8132
rect 6288 7644 6352 7648
rect 6288 7588 6292 7644
rect 6292 7588 6348 7644
rect 6348 7588 6352 7644
rect 6288 7584 6352 7588
rect 6368 7644 6432 7648
rect 6368 7588 6372 7644
rect 6372 7588 6428 7644
rect 6428 7588 6432 7644
rect 6368 7584 6432 7588
rect 6448 7644 6512 7648
rect 6448 7588 6452 7644
rect 6452 7588 6508 7644
rect 6508 7588 6512 7644
rect 6448 7584 6512 7588
rect 6528 7644 6592 7648
rect 6528 7588 6532 7644
rect 6532 7588 6588 7644
rect 6588 7588 6592 7644
rect 6528 7584 6592 7588
rect 13648 7644 13712 7648
rect 13648 7588 13652 7644
rect 13652 7588 13708 7644
rect 13708 7588 13712 7644
rect 13648 7584 13712 7588
rect 13728 7644 13792 7648
rect 13728 7588 13732 7644
rect 13732 7588 13788 7644
rect 13788 7588 13792 7644
rect 13728 7584 13792 7588
rect 13808 7644 13872 7648
rect 13808 7588 13812 7644
rect 13812 7588 13868 7644
rect 13868 7588 13872 7644
rect 13808 7584 13872 7588
rect 13888 7644 13952 7648
rect 13888 7588 13892 7644
rect 13892 7588 13948 7644
rect 13948 7588 13952 7644
rect 13888 7584 13952 7588
rect 21008 7644 21072 7648
rect 21008 7588 21012 7644
rect 21012 7588 21068 7644
rect 21068 7588 21072 7644
rect 21008 7584 21072 7588
rect 21088 7644 21152 7648
rect 21088 7588 21092 7644
rect 21092 7588 21148 7644
rect 21148 7588 21152 7644
rect 21088 7584 21152 7588
rect 21168 7644 21232 7648
rect 21168 7588 21172 7644
rect 21172 7588 21228 7644
rect 21228 7588 21232 7644
rect 21168 7584 21232 7588
rect 21248 7644 21312 7648
rect 21248 7588 21252 7644
rect 21252 7588 21308 7644
rect 21308 7588 21312 7644
rect 21248 7584 21312 7588
rect 28368 7644 28432 7648
rect 28368 7588 28372 7644
rect 28372 7588 28428 7644
rect 28428 7588 28432 7644
rect 28368 7584 28432 7588
rect 28448 7644 28512 7648
rect 28448 7588 28452 7644
rect 28452 7588 28508 7644
rect 28508 7588 28512 7644
rect 28448 7584 28512 7588
rect 28528 7644 28592 7648
rect 28528 7588 28532 7644
rect 28532 7588 28588 7644
rect 28588 7588 28592 7644
rect 28528 7584 28592 7588
rect 28608 7644 28672 7648
rect 28608 7588 28612 7644
rect 28612 7588 28668 7644
rect 28668 7588 28672 7644
rect 28608 7584 28672 7588
rect 6948 7100 7012 7104
rect 6948 7044 6952 7100
rect 6952 7044 7008 7100
rect 7008 7044 7012 7100
rect 6948 7040 7012 7044
rect 7028 7100 7092 7104
rect 7028 7044 7032 7100
rect 7032 7044 7088 7100
rect 7088 7044 7092 7100
rect 7028 7040 7092 7044
rect 7108 7100 7172 7104
rect 7108 7044 7112 7100
rect 7112 7044 7168 7100
rect 7168 7044 7172 7100
rect 7108 7040 7172 7044
rect 7188 7100 7252 7104
rect 7188 7044 7192 7100
rect 7192 7044 7248 7100
rect 7248 7044 7252 7100
rect 7188 7040 7252 7044
rect 14308 7100 14372 7104
rect 14308 7044 14312 7100
rect 14312 7044 14368 7100
rect 14368 7044 14372 7100
rect 14308 7040 14372 7044
rect 14388 7100 14452 7104
rect 14388 7044 14392 7100
rect 14392 7044 14448 7100
rect 14448 7044 14452 7100
rect 14388 7040 14452 7044
rect 14468 7100 14532 7104
rect 14468 7044 14472 7100
rect 14472 7044 14528 7100
rect 14528 7044 14532 7100
rect 14468 7040 14532 7044
rect 14548 7100 14612 7104
rect 14548 7044 14552 7100
rect 14552 7044 14608 7100
rect 14608 7044 14612 7100
rect 14548 7040 14612 7044
rect 21668 7100 21732 7104
rect 21668 7044 21672 7100
rect 21672 7044 21728 7100
rect 21728 7044 21732 7100
rect 21668 7040 21732 7044
rect 21748 7100 21812 7104
rect 21748 7044 21752 7100
rect 21752 7044 21808 7100
rect 21808 7044 21812 7100
rect 21748 7040 21812 7044
rect 21828 7100 21892 7104
rect 21828 7044 21832 7100
rect 21832 7044 21888 7100
rect 21888 7044 21892 7100
rect 21828 7040 21892 7044
rect 21908 7100 21972 7104
rect 21908 7044 21912 7100
rect 21912 7044 21968 7100
rect 21968 7044 21972 7100
rect 21908 7040 21972 7044
rect 29028 7100 29092 7104
rect 29028 7044 29032 7100
rect 29032 7044 29088 7100
rect 29088 7044 29092 7100
rect 29028 7040 29092 7044
rect 29108 7100 29172 7104
rect 29108 7044 29112 7100
rect 29112 7044 29168 7100
rect 29168 7044 29172 7100
rect 29108 7040 29172 7044
rect 29188 7100 29252 7104
rect 29188 7044 29192 7100
rect 29192 7044 29248 7100
rect 29248 7044 29252 7100
rect 29188 7040 29252 7044
rect 29268 7100 29332 7104
rect 29268 7044 29272 7100
rect 29272 7044 29328 7100
rect 29328 7044 29332 7100
rect 29268 7040 29332 7044
rect 13308 6836 13372 6900
rect 17724 6836 17788 6900
rect 6288 6556 6352 6560
rect 6288 6500 6292 6556
rect 6292 6500 6348 6556
rect 6348 6500 6352 6556
rect 6288 6496 6352 6500
rect 6368 6556 6432 6560
rect 6368 6500 6372 6556
rect 6372 6500 6428 6556
rect 6428 6500 6432 6556
rect 6368 6496 6432 6500
rect 6448 6556 6512 6560
rect 6448 6500 6452 6556
rect 6452 6500 6508 6556
rect 6508 6500 6512 6556
rect 6448 6496 6512 6500
rect 6528 6556 6592 6560
rect 6528 6500 6532 6556
rect 6532 6500 6588 6556
rect 6588 6500 6592 6556
rect 6528 6496 6592 6500
rect 13648 6556 13712 6560
rect 13648 6500 13652 6556
rect 13652 6500 13708 6556
rect 13708 6500 13712 6556
rect 13648 6496 13712 6500
rect 13728 6556 13792 6560
rect 13728 6500 13732 6556
rect 13732 6500 13788 6556
rect 13788 6500 13792 6556
rect 13728 6496 13792 6500
rect 13808 6556 13872 6560
rect 13808 6500 13812 6556
rect 13812 6500 13868 6556
rect 13868 6500 13872 6556
rect 13808 6496 13872 6500
rect 13888 6556 13952 6560
rect 13888 6500 13892 6556
rect 13892 6500 13948 6556
rect 13948 6500 13952 6556
rect 13888 6496 13952 6500
rect 21008 6556 21072 6560
rect 21008 6500 21012 6556
rect 21012 6500 21068 6556
rect 21068 6500 21072 6556
rect 21008 6496 21072 6500
rect 21088 6556 21152 6560
rect 21088 6500 21092 6556
rect 21092 6500 21148 6556
rect 21148 6500 21152 6556
rect 21088 6496 21152 6500
rect 21168 6556 21232 6560
rect 21168 6500 21172 6556
rect 21172 6500 21228 6556
rect 21228 6500 21232 6556
rect 21168 6496 21232 6500
rect 21248 6556 21312 6560
rect 21248 6500 21252 6556
rect 21252 6500 21308 6556
rect 21308 6500 21312 6556
rect 21248 6496 21312 6500
rect 28368 6556 28432 6560
rect 28368 6500 28372 6556
rect 28372 6500 28428 6556
rect 28428 6500 28432 6556
rect 28368 6496 28432 6500
rect 28448 6556 28512 6560
rect 28448 6500 28452 6556
rect 28452 6500 28508 6556
rect 28508 6500 28512 6556
rect 28448 6496 28512 6500
rect 28528 6556 28592 6560
rect 28528 6500 28532 6556
rect 28532 6500 28588 6556
rect 28588 6500 28592 6556
rect 28528 6496 28592 6500
rect 28608 6556 28672 6560
rect 28608 6500 28612 6556
rect 28612 6500 28668 6556
rect 28668 6500 28672 6556
rect 28608 6496 28672 6500
rect 6948 6012 7012 6016
rect 6948 5956 6952 6012
rect 6952 5956 7008 6012
rect 7008 5956 7012 6012
rect 6948 5952 7012 5956
rect 7028 6012 7092 6016
rect 7028 5956 7032 6012
rect 7032 5956 7088 6012
rect 7088 5956 7092 6012
rect 7028 5952 7092 5956
rect 7108 6012 7172 6016
rect 7108 5956 7112 6012
rect 7112 5956 7168 6012
rect 7168 5956 7172 6012
rect 7108 5952 7172 5956
rect 7188 6012 7252 6016
rect 7188 5956 7192 6012
rect 7192 5956 7248 6012
rect 7248 5956 7252 6012
rect 7188 5952 7252 5956
rect 14308 6012 14372 6016
rect 14308 5956 14312 6012
rect 14312 5956 14368 6012
rect 14368 5956 14372 6012
rect 14308 5952 14372 5956
rect 14388 6012 14452 6016
rect 14388 5956 14392 6012
rect 14392 5956 14448 6012
rect 14448 5956 14452 6012
rect 14388 5952 14452 5956
rect 14468 6012 14532 6016
rect 14468 5956 14472 6012
rect 14472 5956 14528 6012
rect 14528 5956 14532 6012
rect 14468 5952 14532 5956
rect 14548 6012 14612 6016
rect 14548 5956 14552 6012
rect 14552 5956 14608 6012
rect 14608 5956 14612 6012
rect 14548 5952 14612 5956
rect 21668 6012 21732 6016
rect 21668 5956 21672 6012
rect 21672 5956 21728 6012
rect 21728 5956 21732 6012
rect 21668 5952 21732 5956
rect 21748 6012 21812 6016
rect 21748 5956 21752 6012
rect 21752 5956 21808 6012
rect 21808 5956 21812 6012
rect 21748 5952 21812 5956
rect 21828 6012 21892 6016
rect 21828 5956 21832 6012
rect 21832 5956 21888 6012
rect 21888 5956 21892 6012
rect 21828 5952 21892 5956
rect 21908 6012 21972 6016
rect 21908 5956 21912 6012
rect 21912 5956 21968 6012
rect 21968 5956 21972 6012
rect 21908 5952 21972 5956
rect 29028 6012 29092 6016
rect 29028 5956 29032 6012
rect 29032 5956 29088 6012
rect 29088 5956 29092 6012
rect 29028 5952 29092 5956
rect 29108 6012 29172 6016
rect 29108 5956 29112 6012
rect 29112 5956 29168 6012
rect 29168 5956 29172 6012
rect 29108 5952 29172 5956
rect 29188 6012 29252 6016
rect 29188 5956 29192 6012
rect 29192 5956 29248 6012
rect 29248 5956 29252 6012
rect 29188 5952 29252 5956
rect 29268 6012 29332 6016
rect 29268 5956 29272 6012
rect 29272 5956 29328 6012
rect 29328 5956 29332 6012
rect 29268 5952 29332 5956
rect 12940 5536 13004 5540
rect 12940 5480 12990 5536
rect 12990 5480 13004 5536
rect 12940 5476 13004 5480
rect 6288 5468 6352 5472
rect 6288 5412 6292 5468
rect 6292 5412 6348 5468
rect 6348 5412 6352 5468
rect 6288 5408 6352 5412
rect 6368 5468 6432 5472
rect 6368 5412 6372 5468
rect 6372 5412 6428 5468
rect 6428 5412 6432 5468
rect 6368 5408 6432 5412
rect 6448 5468 6512 5472
rect 6448 5412 6452 5468
rect 6452 5412 6508 5468
rect 6508 5412 6512 5468
rect 6448 5408 6512 5412
rect 6528 5468 6592 5472
rect 6528 5412 6532 5468
rect 6532 5412 6588 5468
rect 6588 5412 6592 5468
rect 6528 5408 6592 5412
rect 13648 5468 13712 5472
rect 13648 5412 13652 5468
rect 13652 5412 13708 5468
rect 13708 5412 13712 5468
rect 13648 5408 13712 5412
rect 13728 5468 13792 5472
rect 13728 5412 13732 5468
rect 13732 5412 13788 5468
rect 13788 5412 13792 5468
rect 13728 5408 13792 5412
rect 13808 5468 13872 5472
rect 13808 5412 13812 5468
rect 13812 5412 13868 5468
rect 13868 5412 13872 5468
rect 13808 5408 13872 5412
rect 13888 5468 13952 5472
rect 13888 5412 13892 5468
rect 13892 5412 13948 5468
rect 13948 5412 13952 5468
rect 13888 5408 13952 5412
rect 21008 5468 21072 5472
rect 21008 5412 21012 5468
rect 21012 5412 21068 5468
rect 21068 5412 21072 5468
rect 21008 5408 21072 5412
rect 21088 5468 21152 5472
rect 21088 5412 21092 5468
rect 21092 5412 21148 5468
rect 21148 5412 21152 5468
rect 21088 5408 21152 5412
rect 21168 5468 21232 5472
rect 21168 5412 21172 5468
rect 21172 5412 21228 5468
rect 21228 5412 21232 5468
rect 21168 5408 21232 5412
rect 21248 5468 21312 5472
rect 21248 5412 21252 5468
rect 21252 5412 21308 5468
rect 21308 5412 21312 5468
rect 21248 5408 21312 5412
rect 28368 5468 28432 5472
rect 28368 5412 28372 5468
rect 28372 5412 28428 5468
rect 28428 5412 28432 5468
rect 28368 5408 28432 5412
rect 28448 5468 28512 5472
rect 28448 5412 28452 5468
rect 28452 5412 28508 5468
rect 28508 5412 28512 5468
rect 28448 5408 28512 5412
rect 28528 5468 28592 5472
rect 28528 5412 28532 5468
rect 28532 5412 28588 5468
rect 28588 5412 28592 5468
rect 28528 5408 28592 5412
rect 28608 5468 28672 5472
rect 28608 5412 28612 5468
rect 28612 5412 28668 5468
rect 28668 5412 28672 5468
rect 28608 5408 28672 5412
rect 6948 4924 7012 4928
rect 6948 4868 6952 4924
rect 6952 4868 7008 4924
rect 7008 4868 7012 4924
rect 6948 4864 7012 4868
rect 7028 4924 7092 4928
rect 7028 4868 7032 4924
rect 7032 4868 7088 4924
rect 7088 4868 7092 4924
rect 7028 4864 7092 4868
rect 7108 4924 7172 4928
rect 7108 4868 7112 4924
rect 7112 4868 7168 4924
rect 7168 4868 7172 4924
rect 7108 4864 7172 4868
rect 7188 4924 7252 4928
rect 7188 4868 7192 4924
rect 7192 4868 7248 4924
rect 7248 4868 7252 4924
rect 7188 4864 7252 4868
rect 14308 4924 14372 4928
rect 14308 4868 14312 4924
rect 14312 4868 14368 4924
rect 14368 4868 14372 4924
rect 14308 4864 14372 4868
rect 14388 4924 14452 4928
rect 14388 4868 14392 4924
rect 14392 4868 14448 4924
rect 14448 4868 14452 4924
rect 14388 4864 14452 4868
rect 14468 4924 14532 4928
rect 14468 4868 14472 4924
rect 14472 4868 14528 4924
rect 14528 4868 14532 4924
rect 14468 4864 14532 4868
rect 14548 4924 14612 4928
rect 14548 4868 14552 4924
rect 14552 4868 14608 4924
rect 14608 4868 14612 4924
rect 14548 4864 14612 4868
rect 21668 4924 21732 4928
rect 21668 4868 21672 4924
rect 21672 4868 21728 4924
rect 21728 4868 21732 4924
rect 21668 4864 21732 4868
rect 21748 4924 21812 4928
rect 21748 4868 21752 4924
rect 21752 4868 21808 4924
rect 21808 4868 21812 4924
rect 21748 4864 21812 4868
rect 21828 4924 21892 4928
rect 21828 4868 21832 4924
rect 21832 4868 21888 4924
rect 21888 4868 21892 4924
rect 21828 4864 21892 4868
rect 21908 4924 21972 4928
rect 21908 4868 21912 4924
rect 21912 4868 21968 4924
rect 21968 4868 21972 4924
rect 21908 4864 21972 4868
rect 29028 4924 29092 4928
rect 29028 4868 29032 4924
rect 29032 4868 29088 4924
rect 29088 4868 29092 4924
rect 29028 4864 29092 4868
rect 29108 4924 29172 4928
rect 29108 4868 29112 4924
rect 29112 4868 29168 4924
rect 29168 4868 29172 4924
rect 29108 4864 29172 4868
rect 29188 4924 29252 4928
rect 29188 4868 29192 4924
rect 29192 4868 29248 4924
rect 29248 4868 29252 4924
rect 29188 4864 29252 4868
rect 29268 4924 29332 4928
rect 29268 4868 29272 4924
rect 29272 4868 29328 4924
rect 29328 4868 29332 4924
rect 29268 4864 29332 4868
rect 6288 4380 6352 4384
rect 6288 4324 6292 4380
rect 6292 4324 6348 4380
rect 6348 4324 6352 4380
rect 6288 4320 6352 4324
rect 6368 4380 6432 4384
rect 6368 4324 6372 4380
rect 6372 4324 6428 4380
rect 6428 4324 6432 4380
rect 6368 4320 6432 4324
rect 6448 4380 6512 4384
rect 6448 4324 6452 4380
rect 6452 4324 6508 4380
rect 6508 4324 6512 4380
rect 6448 4320 6512 4324
rect 6528 4380 6592 4384
rect 6528 4324 6532 4380
rect 6532 4324 6588 4380
rect 6588 4324 6592 4380
rect 6528 4320 6592 4324
rect 13648 4380 13712 4384
rect 13648 4324 13652 4380
rect 13652 4324 13708 4380
rect 13708 4324 13712 4380
rect 13648 4320 13712 4324
rect 13728 4380 13792 4384
rect 13728 4324 13732 4380
rect 13732 4324 13788 4380
rect 13788 4324 13792 4380
rect 13728 4320 13792 4324
rect 13808 4380 13872 4384
rect 13808 4324 13812 4380
rect 13812 4324 13868 4380
rect 13868 4324 13872 4380
rect 13808 4320 13872 4324
rect 13888 4380 13952 4384
rect 13888 4324 13892 4380
rect 13892 4324 13948 4380
rect 13948 4324 13952 4380
rect 13888 4320 13952 4324
rect 21008 4380 21072 4384
rect 21008 4324 21012 4380
rect 21012 4324 21068 4380
rect 21068 4324 21072 4380
rect 21008 4320 21072 4324
rect 21088 4380 21152 4384
rect 21088 4324 21092 4380
rect 21092 4324 21148 4380
rect 21148 4324 21152 4380
rect 21088 4320 21152 4324
rect 21168 4380 21232 4384
rect 21168 4324 21172 4380
rect 21172 4324 21228 4380
rect 21228 4324 21232 4380
rect 21168 4320 21232 4324
rect 21248 4380 21312 4384
rect 21248 4324 21252 4380
rect 21252 4324 21308 4380
rect 21308 4324 21312 4380
rect 21248 4320 21312 4324
rect 28368 4380 28432 4384
rect 28368 4324 28372 4380
rect 28372 4324 28428 4380
rect 28428 4324 28432 4380
rect 28368 4320 28432 4324
rect 28448 4380 28512 4384
rect 28448 4324 28452 4380
rect 28452 4324 28508 4380
rect 28508 4324 28512 4380
rect 28448 4320 28512 4324
rect 28528 4380 28592 4384
rect 28528 4324 28532 4380
rect 28532 4324 28588 4380
rect 28588 4324 28592 4380
rect 28528 4320 28592 4324
rect 28608 4380 28672 4384
rect 28608 4324 28612 4380
rect 28612 4324 28668 4380
rect 28668 4324 28672 4380
rect 28608 4320 28672 4324
rect 6948 3836 7012 3840
rect 6948 3780 6952 3836
rect 6952 3780 7008 3836
rect 7008 3780 7012 3836
rect 6948 3776 7012 3780
rect 7028 3836 7092 3840
rect 7028 3780 7032 3836
rect 7032 3780 7088 3836
rect 7088 3780 7092 3836
rect 7028 3776 7092 3780
rect 7108 3836 7172 3840
rect 7108 3780 7112 3836
rect 7112 3780 7168 3836
rect 7168 3780 7172 3836
rect 7108 3776 7172 3780
rect 7188 3836 7252 3840
rect 7188 3780 7192 3836
rect 7192 3780 7248 3836
rect 7248 3780 7252 3836
rect 7188 3776 7252 3780
rect 14308 3836 14372 3840
rect 14308 3780 14312 3836
rect 14312 3780 14368 3836
rect 14368 3780 14372 3836
rect 14308 3776 14372 3780
rect 14388 3836 14452 3840
rect 14388 3780 14392 3836
rect 14392 3780 14448 3836
rect 14448 3780 14452 3836
rect 14388 3776 14452 3780
rect 14468 3836 14532 3840
rect 14468 3780 14472 3836
rect 14472 3780 14528 3836
rect 14528 3780 14532 3836
rect 14468 3776 14532 3780
rect 14548 3836 14612 3840
rect 14548 3780 14552 3836
rect 14552 3780 14608 3836
rect 14608 3780 14612 3836
rect 14548 3776 14612 3780
rect 21668 3836 21732 3840
rect 21668 3780 21672 3836
rect 21672 3780 21728 3836
rect 21728 3780 21732 3836
rect 21668 3776 21732 3780
rect 21748 3836 21812 3840
rect 21748 3780 21752 3836
rect 21752 3780 21808 3836
rect 21808 3780 21812 3836
rect 21748 3776 21812 3780
rect 21828 3836 21892 3840
rect 21828 3780 21832 3836
rect 21832 3780 21888 3836
rect 21888 3780 21892 3836
rect 21828 3776 21892 3780
rect 21908 3836 21972 3840
rect 21908 3780 21912 3836
rect 21912 3780 21968 3836
rect 21968 3780 21972 3836
rect 21908 3776 21972 3780
rect 29028 3836 29092 3840
rect 29028 3780 29032 3836
rect 29032 3780 29088 3836
rect 29088 3780 29092 3836
rect 29028 3776 29092 3780
rect 29108 3836 29172 3840
rect 29108 3780 29112 3836
rect 29112 3780 29168 3836
rect 29168 3780 29172 3836
rect 29108 3776 29172 3780
rect 29188 3836 29252 3840
rect 29188 3780 29192 3836
rect 29192 3780 29248 3836
rect 29248 3780 29252 3836
rect 29188 3776 29252 3780
rect 29268 3836 29332 3840
rect 29268 3780 29272 3836
rect 29272 3780 29328 3836
rect 29328 3780 29332 3836
rect 29268 3776 29332 3780
rect 6288 3292 6352 3296
rect 6288 3236 6292 3292
rect 6292 3236 6348 3292
rect 6348 3236 6352 3292
rect 6288 3232 6352 3236
rect 6368 3292 6432 3296
rect 6368 3236 6372 3292
rect 6372 3236 6428 3292
rect 6428 3236 6432 3292
rect 6368 3232 6432 3236
rect 6448 3292 6512 3296
rect 6448 3236 6452 3292
rect 6452 3236 6508 3292
rect 6508 3236 6512 3292
rect 6448 3232 6512 3236
rect 6528 3292 6592 3296
rect 6528 3236 6532 3292
rect 6532 3236 6588 3292
rect 6588 3236 6592 3292
rect 6528 3232 6592 3236
rect 13648 3292 13712 3296
rect 13648 3236 13652 3292
rect 13652 3236 13708 3292
rect 13708 3236 13712 3292
rect 13648 3232 13712 3236
rect 13728 3292 13792 3296
rect 13728 3236 13732 3292
rect 13732 3236 13788 3292
rect 13788 3236 13792 3292
rect 13728 3232 13792 3236
rect 13808 3292 13872 3296
rect 13808 3236 13812 3292
rect 13812 3236 13868 3292
rect 13868 3236 13872 3292
rect 13808 3232 13872 3236
rect 13888 3292 13952 3296
rect 13888 3236 13892 3292
rect 13892 3236 13948 3292
rect 13948 3236 13952 3292
rect 13888 3232 13952 3236
rect 21008 3292 21072 3296
rect 21008 3236 21012 3292
rect 21012 3236 21068 3292
rect 21068 3236 21072 3292
rect 21008 3232 21072 3236
rect 21088 3292 21152 3296
rect 21088 3236 21092 3292
rect 21092 3236 21148 3292
rect 21148 3236 21152 3292
rect 21088 3232 21152 3236
rect 21168 3292 21232 3296
rect 21168 3236 21172 3292
rect 21172 3236 21228 3292
rect 21228 3236 21232 3292
rect 21168 3232 21232 3236
rect 21248 3292 21312 3296
rect 21248 3236 21252 3292
rect 21252 3236 21308 3292
rect 21308 3236 21312 3292
rect 21248 3232 21312 3236
rect 28368 3292 28432 3296
rect 28368 3236 28372 3292
rect 28372 3236 28428 3292
rect 28428 3236 28432 3292
rect 28368 3232 28432 3236
rect 28448 3292 28512 3296
rect 28448 3236 28452 3292
rect 28452 3236 28508 3292
rect 28508 3236 28512 3292
rect 28448 3232 28512 3236
rect 28528 3292 28592 3296
rect 28528 3236 28532 3292
rect 28532 3236 28588 3292
rect 28588 3236 28592 3292
rect 28528 3232 28592 3236
rect 28608 3292 28672 3296
rect 28608 3236 28612 3292
rect 28612 3236 28668 3292
rect 28668 3236 28672 3292
rect 28608 3232 28672 3236
rect 6948 2748 7012 2752
rect 6948 2692 6952 2748
rect 6952 2692 7008 2748
rect 7008 2692 7012 2748
rect 6948 2688 7012 2692
rect 7028 2748 7092 2752
rect 7028 2692 7032 2748
rect 7032 2692 7088 2748
rect 7088 2692 7092 2748
rect 7028 2688 7092 2692
rect 7108 2748 7172 2752
rect 7108 2692 7112 2748
rect 7112 2692 7168 2748
rect 7168 2692 7172 2748
rect 7108 2688 7172 2692
rect 7188 2748 7252 2752
rect 7188 2692 7192 2748
rect 7192 2692 7248 2748
rect 7248 2692 7252 2748
rect 7188 2688 7252 2692
rect 14308 2748 14372 2752
rect 14308 2692 14312 2748
rect 14312 2692 14368 2748
rect 14368 2692 14372 2748
rect 14308 2688 14372 2692
rect 14388 2748 14452 2752
rect 14388 2692 14392 2748
rect 14392 2692 14448 2748
rect 14448 2692 14452 2748
rect 14388 2688 14452 2692
rect 14468 2748 14532 2752
rect 14468 2692 14472 2748
rect 14472 2692 14528 2748
rect 14528 2692 14532 2748
rect 14468 2688 14532 2692
rect 14548 2748 14612 2752
rect 14548 2692 14552 2748
rect 14552 2692 14608 2748
rect 14608 2692 14612 2748
rect 14548 2688 14612 2692
rect 21668 2748 21732 2752
rect 21668 2692 21672 2748
rect 21672 2692 21728 2748
rect 21728 2692 21732 2748
rect 21668 2688 21732 2692
rect 21748 2748 21812 2752
rect 21748 2692 21752 2748
rect 21752 2692 21808 2748
rect 21808 2692 21812 2748
rect 21748 2688 21812 2692
rect 21828 2748 21892 2752
rect 21828 2692 21832 2748
rect 21832 2692 21888 2748
rect 21888 2692 21892 2748
rect 21828 2688 21892 2692
rect 21908 2748 21972 2752
rect 21908 2692 21912 2748
rect 21912 2692 21968 2748
rect 21968 2692 21972 2748
rect 21908 2688 21972 2692
rect 29028 2748 29092 2752
rect 29028 2692 29032 2748
rect 29032 2692 29088 2748
rect 29088 2692 29092 2748
rect 29028 2688 29092 2692
rect 29108 2748 29172 2752
rect 29108 2692 29112 2748
rect 29112 2692 29168 2748
rect 29168 2692 29172 2748
rect 29108 2688 29172 2692
rect 29188 2748 29252 2752
rect 29188 2692 29192 2748
rect 29192 2692 29248 2748
rect 29248 2692 29252 2748
rect 29188 2688 29252 2692
rect 29268 2748 29332 2752
rect 29268 2692 29272 2748
rect 29272 2692 29328 2748
rect 29328 2692 29332 2748
rect 29268 2688 29332 2692
<< metal4 >>
rect 6280 31584 6600 32144
rect 6280 31520 6288 31584
rect 6352 31520 6368 31584
rect 6432 31520 6448 31584
rect 6512 31520 6528 31584
rect 6592 31520 6600 31584
rect 6280 30496 6600 31520
rect 6280 30432 6288 30496
rect 6352 30432 6368 30496
rect 6432 30432 6448 30496
rect 6512 30432 6528 30496
rect 6592 30432 6600 30496
rect 6280 29408 6600 30432
rect 6280 29344 6288 29408
rect 6352 29344 6368 29408
rect 6432 29344 6448 29408
rect 6512 29344 6528 29408
rect 6592 29344 6600 29408
rect 6280 28320 6600 29344
rect 6280 28256 6288 28320
rect 6352 28256 6368 28320
rect 6432 28256 6448 28320
rect 6512 28256 6528 28320
rect 6592 28256 6600 28320
rect 6280 27232 6600 28256
rect 6280 27168 6288 27232
rect 6352 27168 6368 27232
rect 6432 27168 6448 27232
rect 6512 27168 6528 27232
rect 6592 27168 6600 27232
rect 6280 26144 6600 27168
rect 6280 26080 6288 26144
rect 6352 26080 6368 26144
rect 6432 26080 6448 26144
rect 6512 26080 6528 26144
rect 6592 26080 6600 26144
rect 6280 25056 6600 26080
rect 6280 24992 6288 25056
rect 6352 24992 6368 25056
rect 6432 24992 6448 25056
rect 6512 24992 6528 25056
rect 6592 24992 6600 25056
rect 6280 23968 6600 24992
rect 6280 23904 6288 23968
rect 6352 23904 6368 23968
rect 6432 23904 6448 23968
rect 6512 23904 6528 23968
rect 6592 23904 6600 23968
rect 6280 22880 6600 23904
rect 6280 22816 6288 22880
rect 6352 22816 6368 22880
rect 6432 22816 6448 22880
rect 6512 22816 6528 22880
rect 6592 22816 6600 22880
rect 6280 21792 6600 22816
rect 6280 21728 6288 21792
rect 6352 21728 6368 21792
rect 6432 21728 6448 21792
rect 6512 21728 6528 21792
rect 6592 21728 6600 21792
rect 6280 20704 6600 21728
rect 6280 20640 6288 20704
rect 6352 20640 6368 20704
rect 6432 20640 6448 20704
rect 6512 20640 6528 20704
rect 6592 20640 6600 20704
rect 6280 19616 6600 20640
rect 6280 19552 6288 19616
rect 6352 19552 6368 19616
rect 6432 19552 6448 19616
rect 6512 19552 6528 19616
rect 6592 19552 6600 19616
rect 6280 18528 6600 19552
rect 6280 18464 6288 18528
rect 6352 18464 6368 18528
rect 6432 18464 6448 18528
rect 6512 18464 6528 18528
rect 6592 18464 6600 18528
rect 6280 17440 6600 18464
rect 6280 17376 6288 17440
rect 6352 17376 6368 17440
rect 6432 17376 6448 17440
rect 6512 17376 6528 17440
rect 6592 17376 6600 17440
rect 6280 16352 6600 17376
rect 6280 16288 6288 16352
rect 6352 16288 6368 16352
rect 6432 16288 6448 16352
rect 6512 16288 6528 16352
rect 6592 16288 6600 16352
rect 6280 15264 6600 16288
rect 6280 15200 6288 15264
rect 6352 15200 6368 15264
rect 6432 15200 6448 15264
rect 6512 15200 6528 15264
rect 6592 15200 6600 15264
rect 6280 14176 6600 15200
rect 6280 14112 6288 14176
rect 6352 14112 6368 14176
rect 6432 14112 6448 14176
rect 6512 14112 6528 14176
rect 6592 14112 6600 14176
rect 6280 13088 6600 14112
rect 6280 13024 6288 13088
rect 6352 13024 6368 13088
rect 6432 13024 6448 13088
rect 6512 13024 6528 13088
rect 6592 13024 6600 13088
rect 6280 12000 6600 13024
rect 6280 11936 6288 12000
rect 6352 11936 6368 12000
rect 6432 11936 6448 12000
rect 6512 11936 6528 12000
rect 6592 11936 6600 12000
rect 6280 10912 6600 11936
rect 6280 10848 6288 10912
rect 6352 10848 6368 10912
rect 6432 10848 6448 10912
rect 6512 10848 6528 10912
rect 6592 10848 6600 10912
rect 6280 9824 6600 10848
rect 6280 9760 6288 9824
rect 6352 9760 6368 9824
rect 6432 9760 6448 9824
rect 6512 9760 6528 9824
rect 6592 9760 6600 9824
rect 6280 8736 6600 9760
rect 6280 8672 6288 8736
rect 6352 8672 6368 8736
rect 6432 8672 6448 8736
rect 6512 8672 6528 8736
rect 6592 8672 6600 8736
rect 6280 7648 6600 8672
rect 6280 7584 6288 7648
rect 6352 7584 6368 7648
rect 6432 7584 6448 7648
rect 6512 7584 6528 7648
rect 6592 7584 6600 7648
rect 6280 6560 6600 7584
rect 6280 6496 6288 6560
rect 6352 6496 6368 6560
rect 6432 6496 6448 6560
rect 6512 6496 6528 6560
rect 6592 6496 6600 6560
rect 6280 5472 6600 6496
rect 6280 5408 6288 5472
rect 6352 5408 6368 5472
rect 6432 5408 6448 5472
rect 6512 5408 6528 5472
rect 6592 5408 6600 5472
rect 6280 4384 6600 5408
rect 6280 4320 6288 4384
rect 6352 4320 6368 4384
rect 6432 4320 6448 4384
rect 6512 4320 6528 4384
rect 6592 4320 6600 4384
rect 6280 3296 6600 4320
rect 6280 3232 6288 3296
rect 6352 3232 6368 3296
rect 6432 3232 6448 3296
rect 6512 3232 6528 3296
rect 6592 3232 6600 3296
rect 6280 2672 6600 3232
rect 6940 32128 7260 32144
rect 6940 32064 6948 32128
rect 7012 32064 7028 32128
rect 7092 32064 7108 32128
rect 7172 32064 7188 32128
rect 7252 32064 7260 32128
rect 6940 31040 7260 32064
rect 13307 31924 13373 31925
rect 13307 31860 13308 31924
rect 13372 31860 13373 31924
rect 13307 31859 13373 31860
rect 6940 30976 6948 31040
rect 7012 30976 7028 31040
rect 7092 30976 7108 31040
rect 7172 30976 7188 31040
rect 7252 30976 7260 31040
rect 6940 29952 7260 30976
rect 6940 29888 6948 29952
rect 7012 29888 7028 29952
rect 7092 29888 7108 29952
rect 7172 29888 7188 29952
rect 7252 29888 7260 29952
rect 6940 28864 7260 29888
rect 6940 28800 6948 28864
rect 7012 28800 7028 28864
rect 7092 28800 7108 28864
rect 7172 28800 7188 28864
rect 7252 28800 7260 28864
rect 6940 27776 7260 28800
rect 6940 27712 6948 27776
rect 7012 27712 7028 27776
rect 7092 27712 7108 27776
rect 7172 27712 7188 27776
rect 7252 27712 7260 27776
rect 6940 26688 7260 27712
rect 11099 27708 11165 27709
rect 11099 27644 11100 27708
rect 11164 27644 11165 27708
rect 11099 27643 11165 27644
rect 6940 26624 6948 26688
rect 7012 26624 7028 26688
rect 7092 26624 7108 26688
rect 7172 26624 7188 26688
rect 7252 26624 7260 26688
rect 6940 25600 7260 26624
rect 6940 25536 6948 25600
rect 7012 25536 7028 25600
rect 7092 25536 7108 25600
rect 7172 25536 7188 25600
rect 7252 25536 7260 25600
rect 6940 24512 7260 25536
rect 6940 24448 6948 24512
rect 7012 24448 7028 24512
rect 7092 24448 7108 24512
rect 7172 24448 7188 24512
rect 7252 24448 7260 24512
rect 6940 23424 7260 24448
rect 6940 23360 6948 23424
rect 7012 23360 7028 23424
rect 7092 23360 7108 23424
rect 7172 23360 7188 23424
rect 7252 23360 7260 23424
rect 6940 22336 7260 23360
rect 6940 22272 6948 22336
rect 7012 22272 7028 22336
rect 7092 22272 7108 22336
rect 7172 22272 7188 22336
rect 7252 22272 7260 22336
rect 6940 21248 7260 22272
rect 6940 21184 6948 21248
rect 7012 21184 7028 21248
rect 7092 21184 7108 21248
rect 7172 21184 7188 21248
rect 7252 21184 7260 21248
rect 6940 20160 7260 21184
rect 6940 20096 6948 20160
rect 7012 20096 7028 20160
rect 7092 20096 7108 20160
rect 7172 20096 7188 20160
rect 7252 20096 7260 20160
rect 6940 19072 7260 20096
rect 6940 19008 6948 19072
rect 7012 19008 7028 19072
rect 7092 19008 7108 19072
rect 7172 19008 7188 19072
rect 7252 19008 7260 19072
rect 6940 17984 7260 19008
rect 6940 17920 6948 17984
rect 7012 17920 7028 17984
rect 7092 17920 7108 17984
rect 7172 17920 7188 17984
rect 7252 17920 7260 17984
rect 6940 16896 7260 17920
rect 6940 16832 6948 16896
rect 7012 16832 7028 16896
rect 7092 16832 7108 16896
rect 7172 16832 7188 16896
rect 7252 16832 7260 16896
rect 6940 15808 7260 16832
rect 11102 16557 11162 27643
rect 11283 25804 11349 25805
rect 11283 25740 11284 25804
rect 11348 25740 11349 25804
rect 11283 25739 11349 25740
rect 11286 20501 11346 25739
rect 13123 23764 13189 23765
rect 13123 23700 13124 23764
rect 13188 23700 13189 23764
rect 13123 23699 13189 23700
rect 11283 20500 11349 20501
rect 11283 20436 11284 20500
rect 11348 20436 11349 20500
rect 11283 20435 11349 20436
rect 12939 19412 13005 19413
rect 12939 19348 12940 19412
rect 13004 19348 13005 19412
rect 12939 19347 13005 19348
rect 12203 19276 12269 19277
rect 12203 19212 12204 19276
rect 12268 19212 12269 19276
rect 12203 19211 12269 19212
rect 11099 16556 11165 16557
rect 11099 16492 11100 16556
rect 11164 16492 11165 16556
rect 11099 16491 11165 16492
rect 6940 15744 6948 15808
rect 7012 15744 7028 15808
rect 7092 15744 7108 15808
rect 7172 15744 7188 15808
rect 7252 15744 7260 15808
rect 6940 14720 7260 15744
rect 6940 14656 6948 14720
rect 7012 14656 7028 14720
rect 7092 14656 7108 14720
rect 7172 14656 7188 14720
rect 7252 14656 7260 14720
rect 6940 13632 7260 14656
rect 12206 14245 12266 19211
rect 12203 14244 12269 14245
rect 12203 14180 12204 14244
rect 12268 14180 12269 14244
rect 12203 14179 12269 14180
rect 6940 13568 6948 13632
rect 7012 13568 7028 13632
rect 7092 13568 7108 13632
rect 7172 13568 7188 13632
rect 7252 13568 7260 13632
rect 6940 12544 7260 13568
rect 6940 12480 6948 12544
rect 7012 12480 7028 12544
rect 7092 12480 7108 12544
rect 7172 12480 7188 12544
rect 7252 12480 7260 12544
rect 6940 11456 7260 12480
rect 6940 11392 6948 11456
rect 7012 11392 7028 11456
rect 7092 11392 7108 11456
rect 7172 11392 7188 11456
rect 7252 11392 7260 11456
rect 6940 10368 7260 11392
rect 6940 10304 6948 10368
rect 7012 10304 7028 10368
rect 7092 10304 7108 10368
rect 7172 10304 7188 10368
rect 7252 10304 7260 10368
rect 6940 9280 7260 10304
rect 6940 9216 6948 9280
rect 7012 9216 7028 9280
rect 7092 9216 7108 9280
rect 7172 9216 7188 9280
rect 7252 9216 7260 9280
rect 6940 8192 7260 9216
rect 6940 8128 6948 8192
rect 7012 8128 7028 8192
rect 7092 8128 7108 8192
rect 7172 8128 7188 8192
rect 7252 8128 7260 8192
rect 6940 7104 7260 8128
rect 6940 7040 6948 7104
rect 7012 7040 7028 7104
rect 7092 7040 7108 7104
rect 7172 7040 7188 7104
rect 7252 7040 7260 7104
rect 6940 6016 7260 7040
rect 6940 5952 6948 6016
rect 7012 5952 7028 6016
rect 7092 5952 7108 6016
rect 7172 5952 7188 6016
rect 7252 5952 7260 6016
rect 6940 4928 7260 5952
rect 12942 5541 13002 19347
rect 13126 8261 13186 23699
rect 13123 8260 13189 8261
rect 13123 8196 13124 8260
rect 13188 8196 13189 8260
rect 13123 8195 13189 8196
rect 13310 6901 13370 31859
rect 13640 31584 13960 32144
rect 13640 31520 13648 31584
rect 13712 31520 13728 31584
rect 13792 31520 13808 31584
rect 13872 31520 13888 31584
rect 13952 31520 13960 31584
rect 13640 30496 13960 31520
rect 13640 30432 13648 30496
rect 13712 30432 13728 30496
rect 13792 30432 13808 30496
rect 13872 30432 13888 30496
rect 13952 30432 13960 30496
rect 13640 29408 13960 30432
rect 13640 29344 13648 29408
rect 13712 29344 13728 29408
rect 13792 29344 13808 29408
rect 13872 29344 13888 29408
rect 13952 29344 13960 29408
rect 13640 28320 13960 29344
rect 13640 28256 13648 28320
rect 13712 28256 13728 28320
rect 13792 28256 13808 28320
rect 13872 28256 13888 28320
rect 13952 28256 13960 28320
rect 13640 27232 13960 28256
rect 13640 27168 13648 27232
rect 13712 27168 13728 27232
rect 13792 27168 13808 27232
rect 13872 27168 13888 27232
rect 13952 27168 13960 27232
rect 13640 26144 13960 27168
rect 13640 26080 13648 26144
rect 13712 26080 13728 26144
rect 13792 26080 13808 26144
rect 13872 26080 13888 26144
rect 13952 26080 13960 26144
rect 13640 25056 13960 26080
rect 13640 24992 13648 25056
rect 13712 24992 13728 25056
rect 13792 24992 13808 25056
rect 13872 24992 13888 25056
rect 13952 24992 13960 25056
rect 13640 23968 13960 24992
rect 13640 23904 13648 23968
rect 13712 23904 13728 23968
rect 13792 23904 13808 23968
rect 13872 23904 13888 23968
rect 13952 23904 13960 23968
rect 13640 22880 13960 23904
rect 13640 22816 13648 22880
rect 13712 22816 13728 22880
rect 13792 22816 13808 22880
rect 13872 22816 13888 22880
rect 13952 22816 13960 22880
rect 13640 21792 13960 22816
rect 13640 21728 13648 21792
rect 13712 21728 13728 21792
rect 13792 21728 13808 21792
rect 13872 21728 13888 21792
rect 13952 21728 13960 21792
rect 13640 20704 13960 21728
rect 13640 20640 13648 20704
rect 13712 20640 13728 20704
rect 13792 20640 13808 20704
rect 13872 20640 13888 20704
rect 13952 20640 13960 20704
rect 13640 19616 13960 20640
rect 13640 19552 13648 19616
rect 13712 19552 13728 19616
rect 13792 19552 13808 19616
rect 13872 19552 13888 19616
rect 13952 19552 13960 19616
rect 13640 18528 13960 19552
rect 13640 18464 13648 18528
rect 13712 18464 13728 18528
rect 13792 18464 13808 18528
rect 13872 18464 13888 18528
rect 13952 18464 13960 18528
rect 13640 17440 13960 18464
rect 13640 17376 13648 17440
rect 13712 17376 13728 17440
rect 13792 17376 13808 17440
rect 13872 17376 13888 17440
rect 13952 17376 13960 17440
rect 13640 16352 13960 17376
rect 13640 16288 13648 16352
rect 13712 16288 13728 16352
rect 13792 16288 13808 16352
rect 13872 16288 13888 16352
rect 13952 16288 13960 16352
rect 13640 15264 13960 16288
rect 13640 15200 13648 15264
rect 13712 15200 13728 15264
rect 13792 15200 13808 15264
rect 13872 15200 13888 15264
rect 13952 15200 13960 15264
rect 13640 14176 13960 15200
rect 13640 14112 13648 14176
rect 13712 14112 13728 14176
rect 13792 14112 13808 14176
rect 13872 14112 13888 14176
rect 13952 14112 13960 14176
rect 13640 13088 13960 14112
rect 13640 13024 13648 13088
rect 13712 13024 13728 13088
rect 13792 13024 13808 13088
rect 13872 13024 13888 13088
rect 13952 13024 13960 13088
rect 13640 12000 13960 13024
rect 13640 11936 13648 12000
rect 13712 11936 13728 12000
rect 13792 11936 13808 12000
rect 13872 11936 13888 12000
rect 13952 11936 13960 12000
rect 13640 10912 13960 11936
rect 13640 10848 13648 10912
rect 13712 10848 13728 10912
rect 13792 10848 13808 10912
rect 13872 10848 13888 10912
rect 13952 10848 13960 10912
rect 13640 9824 13960 10848
rect 13640 9760 13648 9824
rect 13712 9760 13728 9824
rect 13792 9760 13808 9824
rect 13872 9760 13888 9824
rect 13952 9760 13960 9824
rect 13640 8736 13960 9760
rect 13640 8672 13648 8736
rect 13712 8672 13728 8736
rect 13792 8672 13808 8736
rect 13872 8672 13888 8736
rect 13952 8672 13960 8736
rect 13640 7648 13960 8672
rect 13640 7584 13648 7648
rect 13712 7584 13728 7648
rect 13792 7584 13808 7648
rect 13872 7584 13888 7648
rect 13952 7584 13960 7648
rect 13307 6900 13373 6901
rect 13307 6836 13308 6900
rect 13372 6836 13373 6900
rect 13307 6835 13373 6836
rect 13640 6560 13960 7584
rect 13640 6496 13648 6560
rect 13712 6496 13728 6560
rect 13792 6496 13808 6560
rect 13872 6496 13888 6560
rect 13952 6496 13960 6560
rect 12939 5540 13005 5541
rect 12939 5476 12940 5540
rect 13004 5476 13005 5540
rect 12939 5475 13005 5476
rect 6940 4864 6948 4928
rect 7012 4864 7028 4928
rect 7092 4864 7108 4928
rect 7172 4864 7188 4928
rect 7252 4864 7260 4928
rect 6940 3840 7260 4864
rect 6940 3776 6948 3840
rect 7012 3776 7028 3840
rect 7092 3776 7108 3840
rect 7172 3776 7188 3840
rect 7252 3776 7260 3840
rect 6940 2752 7260 3776
rect 6940 2688 6948 2752
rect 7012 2688 7028 2752
rect 7092 2688 7108 2752
rect 7172 2688 7188 2752
rect 7252 2688 7260 2752
rect 6940 2672 7260 2688
rect 13640 5472 13960 6496
rect 13640 5408 13648 5472
rect 13712 5408 13728 5472
rect 13792 5408 13808 5472
rect 13872 5408 13888 5472
rect 13952 5408 13960 5472
rect 13640 4384 13960 5408
rect 13640 4320 13648 4384
rect 13712 4320 13728 4384
rect 13792 4320 13808 4384
rect 13872 4320 13888 4384
rect 13952 4320 13960 4384
rect 13640 3296 13960 4320
rect 13640 3232 13648 3296
rect 13712 3232 13728 3296
rect 13792 3232 13808 3296
rect 13872 3232 13888 3296
rect 13952 3232 13960 3296
rect 13640 2672 13960 3232
rect 14300 32128 14620 32144
rect 14300 32064 14308 32128
rect 14372 32064 14388 32128
rect 14452 32064 14468 32128
rect 14532 32064 14548 32128
rect 14612 32064 14620 32128
rect 14300 31040 14620 32064
rect 17723 31788 17789 31789
rect 17723 31724 17724 31788
rect 17788 31724 17789 31788
rect 17723 31723 17789 31724
rect 14300 30976 14308 31040
rect 14372 30976 14388 31040
rect 14452 30976 14468 31040
rect 14532 30976 14548 31040
rect 14612 30976 14620 31040
rect 14300 29952 14620 30976
rect 14300 29888 14308 29952
rect 14372 29888 14388 29952
rect 14452 29888 14468 29952
rect 14532 29888 14548 29952
rect 14612 29888 14620 29952
rect 14300 28864 14620 29888
rect 14300 28800 14308 28864
rect 14372 28800 14388 28864
rect 14452 28800 14468 28864
rect 14532 28800 14548 28864
rect 14612 28800 14620 28864
rect 14300 27776 14620 28800
rect 16619 28116 16685 28117
rect 16619 28052 16620 28116
rect 16684 28052 16685 28116
rect 16619 28051 16685 28052
rect 14300 27712 14308 27776
rect 14372 27712 14388 27776
rect 14452 27712 14468 27776
rect 14532 27712 14548 27776
rect 14612 27712 14620 27776
rect 14300 26688 14620 27712
rect 14300 26624 14308 26688
rect 14372 26624 14388 26688
rect 14452 26624 14468 26688
rect 14532 26624 14548 26688
rect 14612 26624 14620 26688
rect 14300 25600 14620 26624
rect 14300 25536 14308 25600
rect 14372 25536 14388 25600
rect 14452 25536 14468 25600
rect 14532 25536 14548 25600
rect 14612 25536 14620 25600
rect 14300 24512 14620 25536
rect 14300 24448 14308 24512
rect 14372 24448 14388 24512
rect 14452 24448 14468 24512
rect 14532 24448 14548 24512
rect 14612 24448 14620 24512
rect 14300 23424 14620 24448
rect 14300 23360 14308 23424
rect 14372 23360 14388 23424
rect 14452 23360 14468 23424
rect 14532 23360 14548 23424
rect 14612 23360 14620 23424
rect 14300 22336 14620 23360
rect 14300 22272 14308 22336
rect 14372 22272 14388 22336
rect 14452 22272 14468 22336
rect 14532 22272 14548 22336
rect 14612 22272 14620 22336
rect 14300 21248 14620 22272
rect 14300 21184 14308 21248
rect 14372 21184 14388 21248
rect 14452 21184 14468 21248
rect 14532 21184 14548 21248
rect 14612 21184 14620 21248
rect 14300 20160 14620 21184
rect 14779 20772 14845 20773
rect 14779 20708 14780 20772
rect 14844 20708 14845 20772
rect 14779 20707 14845 20708
rect 16435 20772 16501 20773
rect 16435 20708 16436 20772
rect 16500 20708 16501 20772
rect 16435 20707 16501 20708
rect 14300 20096 14308 20160
rect 14372 20096 14388 20160
rect 14452 20096 14468 20160
rect 14532 20096 14548 20160
rect 14612 20096 14620 20160
rect 14300 19072 14620 20096
rect 14300 19008 14308 19072
rect 14372 19008 14388 19072
rect 14452 19008 14468 19072
rect 14532 19008 14548 19072
rect 14612 19008 14620 19072
rect 14300 17984 14620 19008
rect 14300 17920 14308 17984
rect 14372 17920 14388 17984
rect 14452 17920 14468 17984
rect 14532 17920 14548 17984
rect 14612 17920 14620 17984
rect 14300 16896 14620 17920
rect 14300 16832 14308 16896
rect 14372 16832 14388 16896
rect 14452 16832 14468 16896
rect 14532 16832 14548 16896
rect 14612 16832 14620 16896
rect 14300 15808 14620 16832
rect 14300 15744 14308 15808
rect 14372 15744 14388 15808
rect 14452 15744 14468 15808
rect 14532 15744 14548 15808
rect 14612 15744 14620 15808
rect 14300 14720 14620 15744
rect 14300 14656 14308 14720
rect 14372 14656 14388 14720
rect 14452 14656 14468 14720
rect 14532 14656 14548 14720
rect 14612 14656 14620 14720
rect 14300 13632 14620 14656
rect 14300 13568 14308 13632
rect 14372 13568 14388 13632
rect 14452 13568 14468 13632
rect 14532 13568 14548 13632
rect 14612 13568 14620 13632
rect 14300 12544 14620 13568
rect 14300 12480 14308 12544
rect 14372 12480 14388 12544
rect 14452 12480 14468 12544
rect 14532 12480 14548 12544
rect 14612 12480 14620 12544
rect 14300 11456 14620 12480
rect 14300 11392 14308 11456
rect 14372 11392 14388 11456
rect 14452 11392 14468 11456
rect 14532 11392 14548 11456
rect 14612 11392 14620 11456
rect 14300 10368 14620 11392
rect 14782 11253 14842 20707
rect 15331 19956 15397 19957
rect 15331 19892 15332 19956
rect 15396 19892 15397 19956
rect 15331 19891 15397 19892
rect 15334 15197 15394 19891
rect 15331 15196 15397 15197
rect 15331 15132 15332 15196
rect 15396 15132 15397 15196
rect 15331 15131 15397 15132
rect 16438 13701 16498 20707
rect 16622 16557 16682 28051
rect 16619 16556 16685 16557
rect 16619 16492 16620 16556
rect 16684 16492 16685 16556
rect 16619 16491 16685 16492
rect 16435 13700 16501 13701
rect 16435 13636 16436 13700
rect 16500 13636 16501 13700
rect 16435 13635 16501 13636
rect 14779 11252 14845 11253
rect 14779 11188 14780 11252
rect 14844 11188 14845 11252
rect 14779 11187 14845 11188
rect 14300 10304 14308 10368
rect 14372 10304 14388 10368
rect 14452 10304 14468 10368
rect 14532 10304 14548 10368
rect 14612 10304 14620 10368
rect 14300 9280 14620 10304
rect 14300 9216 14308 9280
rect 14372 9216 14388 9280
rect 14452 9216 14468 9280
rect 14532 9216 14548 9280
rect 14612 9216 14620 9280
rect 14300 8192 14620 9216
rect 14300 8128 14308 8192
rect 14372 8128 14388 8192
rect 14452 8128 14468 8192
rect 14532 8128 14548 8192
rect 14612 8128 14620 8192
rect 14300 7104 14620 8128
rect 14300 7040 14308 7104
rect 14372 7040 14388 7104
rect 14452 7040 14468 7104
rect 14532 7040 14548 7104
rect 14612 7040 14620 7104
rect 14300 6016 14620 7040
rect 17726 6901 17786 31723
rect 21000 31584 21320 32144
rect 21000 31520 21008 31584
rect 21072 31520 21088 31584
rect 21152 31520 21168 31584
rect 21232 31520 21248 31584
rect 21312 31520 21320 31584
rect 21000 30496 21320 31520
rect 21000 30432 21008 30496
rect 21072 30432 21088 30496
rect 21152 30432 21168 30496
rect 21232 30432 21248 30496
rect 21312 30432 21320 30496
rect 21000 29408 21320 30432
rect 21000 29344 21008 29408
rect 21072 29344 21088 29408
rect 21152 29344 21168 29408
rect 21232 29344 21248 29408
rect 21312 29344 21320 29408
rect 21000 28320 21320 29344
rect 21000 28256 21008 28320
rect 21072 28256 21088 28320
rect 21152 28256 21168 28320
rect 21232 28256 21248 28320
rect 21312 28256 21320 28320
rect 21000 27232 21320 28256
rect 21000 27168 21008 27232
rect 21072 27168 21088 27232
rect 21152 27168 21168 27232
rect 21232 27168 21248 27232
rect 21312 27168 21320 27232
rect 21000 26144 21320 27168
rect 21000 26080 21008 26144
rect 21072 26080 21088 26144
rect 21152 26080 21168 26144
rect 21232 26080 21248 26144
rect 21312 26080 21320 26144
rect 21000 25056 21320 26080
rect 21000 24992 21008 25056
rect 21072 24992 21088 25056
rect 21152 24992 21168 25056
rect 21232 24992 21248 25056
rect 21312 24992 21320 25056
rect 21000 23968 21320 24992
rect 21000 23904 21008 23968
rect 21072 23904 21088 23968
rect 21152 23904 21168 23968
rect 21232 23904 21248 23968
rect 21312 23904 21320 23968
rect 21000 22880 21320 23904
rect 21000 22816 21008 22880
rect 21072 22816 21088 22880
rect 21152 22816 21168 22880
rect 21232 22816 21248 22880
rect 21312 22816 21320 22880
rect 21000 21792 21320 22816
rect 21000 21728 21008 21792
rect 21072 21728 21088 21792
rect 21152 21728 21168 21792
rect 21232 21728 21248 21792
rect 21312 21728 21320 21792
rect 21000 20704 21320 21728
rect 21000 20640 21008 20704
rect 21072 20640 21088 20704
rect 21152 20640 21168 20704
rect 21232 20640 21248 20704
rect 21312 20640 21320 20704
rect 21000 19616 21320 20640
rect 21000 19552 21008 19616
rect 21072 19552 21088 19616
rect 21152 19552 21168 19616
rect 21232 19552 21248 19616
rect 21312 19552 21320 19616
rect 21000 18528 21320 19552
rect 21000 18464 21008 18528
rect 21072 18464 21088 18528
rect 21152 18464 21168 18528
rect 21232 18464 21248 18528
rect 21312 18464 21320 18528
rect 21000 17440 21320 18464
rect 21000 17376 21008 17440
rect 21072 17376 21088 17440
rect 21152 17376 21168 17440
rect 21232 17376 21248 17440
rect 21312 17376 21320 17440
rect 21000 16352 21320 17376
rect 21000 16288 21008 16352
rect 21072 16288 21088 16352
rect 21152 16288 21168 16352
rect 21232 16288 21248 16352
rect 21312 16288 21320 16352
rect 21000 15264 21320 16288
rect 21000 15200 21008 15264
rect 21072 15200 21088 15264
rect 21152 15200 21168 15264
rect 21232 15200 21248 15264
rect 21312 15200 21320 15264
rect 21000 14176 21320 15200
rect 21000 14112 21008 14176
rect 21072 14112 21088 14176
rect 21152 14112 21168 14176
rect 21232 14112 21248 14176
rect 21312 14112 21320 14176
rect 21000 13088 21320 14112
rect 21000 13024 21008 13088
rect 21072 13024 21088 13088
rect 21152 13024 21168 13088
rect 21232 13024 21248 13088
rect 21312 13024 21320 13088
rect 21000 12000 21320 13024
rect 21000 11936 21008 12000
rect 21072 11936 21088 12000
rect 21152 11936 21168 12000
rect 21232 11936 21248 12000
rect 21312 11936 21320 12000
rect 21000 10912 21320 11936
rect 21000 10848 21008 10912
rect 21072 10848 21088 10912
rect 21152 10848 21168 10912
rect 21232 10848 21248 10912
rect 21312 10848 21320 10912
rect 21000 9824 21320 10848
rect 21000 9760 21008 9824
rect 21072 9760 21088 9824
rect 21152 9760 21168 9824
rect 21232 9760 21248 9824
rect 21312 9760 21320 9824
rect 21000 8736 21320 9760
rect 21000 8672 21008 8736
rect 21072 8672 21088 8736
rect 21152 8672 21168 8736
rect 21232 8672 21248 8736
rect 21312 8672 21320 8736
rect 21000 7648 21320 8672
rect 21000 7584 21008 7648
rect 21072 7584 21088 7648
rect 21152 7584 21168 7648
rect 21232 7584 21248 7648
rect 21312 7584 21320 7648
rect 17723 6900 17789 6901
rect 17723 6836 17724 6900
rect 17788 6836 17789 6900
rect 17723 6835 17789 6836
rect 14300 5952 14308 6016
rect 14372 5952 14388 6016
rect 14452 5952 14468 6016
rect 14532 5952 14548 6016
rect 14612 5952 14620 6016
rect 14300 4928 14620 5952
rect 14300 4864 14308 4928
rect 14372 4864 14388 4928
rect 14452 4864 14468 4928
rect 14532 4864 14548 4928
rect 14612 4864 14620 4928
rect 14300 3840 14620 4864
rect 14300 3776 14308 3840
rect 14372 3776 14388 3840
rect 14452 3776 14468 3840
rect 14532 3776 14548 3840
rect 14612 3776 14620 3840
rect 14300 2752 14620 3776
rect 14300 2688 14308 2752
rect 14372 2688 14388 2752
rect 14452 2688 14468 2752
rect 14532 2688 14548 2752
rect 14612 2688 14620 2752
rect 14300 2672 14620 2688
rect 21000 6560 21320 7584
rect 21000 6496 21008 6560
rect 21072 6496 21088 6560
rect 21152 6496 21168 6560
rect 21232 6496 21248 6560
rect 21312 6496 21320 6560
rect 21000 5472 21320 6496
rect 21000 5408 21008 5472
rect 21072 5408 21088 5472
rect 21152 5408 21168 5472
rect 21232 5408 21248 5472
rect 21312 5408 21320 5472
rect 21000 4384 21320 5408
rect 21000 4320 21008 4384
rect 21072 4320 21088 4384
rect 21152 4320 21168 4384
rect 21232 4320 21248 4384
rect 21312 4320 21320 4384
rect 21000 3296 21320 4320
rect 21000 3232 21008 3296
rect 21072 3232 21088 3296
rect 21152 3232 21168 3296
rect 21232 3232 21248 3296
rect 21312 3232 21320 3296
rect 21000 2672 21320 3232
rect 21660 32128 21980 32144
rect 21660 32064 21668 32128
rect 21732 32064 21748 32128
rect 21812 32064 21828 32128
rect 21892 32064 21908 32128
rect 21972 32064 21980 32128
rect 21660 31040 21980 32064
rect 21660 30976 21668 31040
rect 21732 30976 21748 31040
rect 21812 30976 21828 31040
rect 21892 30976 21908 31040
rect 21972 30976 21980 31040
rect 21660 29952 21980 30976
rect 21660 29888 21668 29952
rect 21732 29888 21748 29952
rect 21812 29888 21828 29952
rect 21892 29888 21908 29952
rect 21972 29888 21980 29952
rect 21660 28864 21980 29888
rect 21660 28800 21668 28864
rect 21732 28800 21748 28864
rect 21812 28800 21828 28864
rect 21892 28800 21908 28864
rect 21972 28800 21980 28864
rect 21660 27776 21980 28800
rect 21660 27712 21668 27776
rect 21732 27712 21748 27776
rect 21812 27712 21828 27776
rect 21892 27712 21908 27776
rect 21972 27712 21980 27776
rect 21660 26688 21980 27712
rect 21660 26624 21668 26688
rect 21732 26624 21748 26688
rect 21812 26624 21828 26688
rect 21892 26624 21908 26688
rect 21972 26624 21980 26688
rect 21660 25600 21980 26624
rect 21660 25536 21668 25600
rect 21732 25536 21748 25600
rect 21812 25536 21828 25600
rect 21892 25536 21908 25600
rect 21972 25536 21980 25600
rect 21660 24512 21980 25536
rect 21660 24448 21668 24512
rect 21732 24448 21748 24512
rect 21812 24448 21828 24512
rect 21892 24448 21908 24512
rect 21972 24448 21980 24512
rect 21660 23424 21980 24448
rect 21660 23360 21668 23424
rect 21732 23360 21748 23424
rect 21812 23360 21828 23424
rect 21892 23360 21908 23424
rect 21972 23360 21980 23424
rect 21660 22336 21980 23360
rect 21660 22272 21668 22336
rect 21732 22272 21748 22336
rect 21812 22272 21828 22336
rect 21892 22272 21908 22336
rect 21972 22272 21980 22336
rect 21660 21248 21980 22272
rect 21660 21184 21668 21248
rect 21732 21184 21748 21248
rect 21812 21184 21828 21248
rect 21892 21184 21908 21248
rect 21972 21184 21980 21248
rect 21660 20160 21980 21184
rect 28360 31584 28680 32144
rect 28360 31520 28368 31584
rect 28432 31520 28448 31584
rect 28512 31520 28528 31584
rect 28592 31520 28608 31584
rect 28672 31520 28680 31584
rect 28360 30496 28680 31520
rect 28360 30432 28368 30496
rect 28432 30432 28448 30496
rect 28512 30432 28528 30496
rect 28592 30432 28608 30496
rect 28672 30432 28680 30496
rect 28360 29408 28680 30432
rect 28360 29344 28368 29408
rect 28432 29344 28448 29408
rect 28512 29344 28528 29408
rect 28592 29344 28608 29408
rect 28672 29344 28680 29408
rect 28360 28320 28680 29344
rect 28360 28256 28368 28320
rect 28432 28256 28448 28320
rect 28512 28256 28528 28320
rect 28592 28256 28608 28320
rect 28672 28256 28680 28320
rect 28360 27232 28680 28256
rect 28360 27168 28368 27232
rect 28432 27168 28448 27232
rect 28512 27168 28528 27232
rect 28592 27168 28608 27232
rect 28672 27168 28680 27232
rect 28360 26144 28680 27168
rect 28360 26080 28368 26144
rect 28432 26080 28448 26144
rect 28512 26080 28528 26144
rect 28592 26080 28608 26144
rect 28672 26080 28680 26144
rect 28360 25056 28680 26080
rect 28360 24992 28368 25056
rect 28432 24992 28448 25056
rect 28512 24992 28528 25056
rect 28592 24992 28608 25056
rect 28672 24992 28680 25056
rect 28360 23968 28680 24992
rect 28360 23904 28368 23968
rect 28432 23904 28448 23968
rect 28512 23904 28528 23968
rect 28592 23904 28608 23968
rect 28672 23904 28680 23968
rect 28360 22880 28680 23904
rect 28360 22816 28368 22880
rect 28432 22816 28448 22880
rect 28512 22816 28528 22880
rect 28592 22816 28608 22880
rect 28672 22816 28680 22880
rect 28360 21792 28680 22816
rect 28360 21728 28368 21792
rect 28432 21728 28448 21792
rect 28512 21728 28528 21792
rect 28592 21728 28608 21792
rect 28672 21728 28680 21792
rect 24531 20908 24597 20909
rect 24531 20844 24532 20908
rect 24596 20844 24597 20908
rect 24531 20843 24597 20844
rect 21660 20096 21668 20160
rect 21732 20096 21748 20160
rect 21812 20096 21828 20160
rect 21892 20096 21908 20160
rect 21972 20096 21980 20160
rect 21660 19072 21980 20096
rect 21660 19008 21668 19072
rect 21732 19008 21748 19072
rect 21812 19008 21828 19072
rect 21892 19008 21908 19072
rect 21972 19008 21980 19072
rect 21660 17984 21980 19008
rect 21660 17920 21668 17984
rect 21732 17920 21748 17984
rect 21812 17920 21828 17984
rect 21892 17920 21908 17984
rect 21972 17920 21980 17984
rect 21660 16896 21980 17920
rect 21660 16832 21668 16896
rect 21732 16832 21748 16896
rect 21812 16832 21828 16896
rect 21892 16832 21908 16896
rect 21972 16832 21980 16896
rect 21660 15808 21980 16832
rect 21660 15744 21668 15808
rect 21732 15744 21748 15808
rect 21812 15744 21828 15808
rect 21892 15744 21908 15808
rect 21972 15744 21980 15808
rect 21660 14720 21980 15744
rect 21660 14656 21668 14720
rect 21732 14656 21748 14720
rect 21812 14656 21828 14720
rect 21892 14656 21908 14720
rect 21972 14656 21980 14720
rect 21660 13632 21980 14656
rect 21660 13568 21668 13632
rect 21732 13568 21748 13632
rect 21812 13568 21828 13632
rect 21892 13568 21908 13632
rect 21972 13568 21980 13632
rect 21660 12544 21980 13568
rect 21660 12480 21668 12544
rect 21732 12480 21748 12544
rect 21812 12480 21828 12544
rect 21892 12480 21908 12544
rect 21972 12480 21980 12544
rect 21660 11456 21980 12480
rect 24534 11933 24594 20843
rect 28360 20704 28680 21728
rect 28360 20640 28368 20704
rect 28432 20640 28448 20704
rect 28512 20640 28528 20704
rect 28592 20640 28608 20704
rect 28672 20640 28680 20704
rect 28360 19616 28680 20640
rect 28360 19552 28368 19616
rect 28432 19552 28448 19616
rect 28512 19552 28528 19616
rect 28592 19552 28608 19616
rect 28672 19552 28680 19616
rect 28360 18528 28680 19552
rect 28360 18464 28368 18528
rect 28432 18464 28448 18528
rect 28512 18464 28528 18528
rect 28592 18464 28608 18528
rect 28672 18464 28680 18528
rect 28360 17440 28680 18464
rect 28360 17376 28368 17440
rect 28432 17376 28448 17440
rect 28512 17376 28528 17440
rect 28592 17376 28608 17440
rect 28672 17376 28680 17440
rect 28360 16352 28680 17376
rect 28360 16288 28368 16352
rect 28432 16288 28448 16352
rect 28512 16288 28528 16352
rect 28592 16288 28608 16352
rect 28672 16288 28680 16352
rect 28360 15264 28680 16288
rect 28360 15200 28368 15264
rect 28432 15200 28448 15264
rect 28512 15200 28528 15264
rect 28592 15200 28608 15264
rect 28672 15200 28680 15264
rect 28360 14176 28680 15200
rect 28360 14112 28368 14176
rect 28432 14112 28448 14176
rect 28512 14112 28528 14176
rect 28592 14112 28608 14176
rect 28672 14112 28680 14176
rect 28360 13088 28680 14112
rect 28360 13024 28368 13088
rect 28432 13024 28448 13088
rect 28512 13024 28528 13088
rect 28592 13024 28608 13088
rect 28672 13024 28680 13088
rect 28360 12000 28680 13024
rect 28360 11936 28368 12000
rect 28432 11936 28448 12000
rect 28512 11936 28528 12000
rect 28592 11936 28608 12000
rect 28672 11936 28680 12000
rect 24531 11932 24597 11933
rect 24531 11868 24532 11932
rect 24596 11868 24597 11932
rect 24531 11867 24597 11868
rect 21660 11392 21668 11456
rect 21732 11392 21748 11456
rect 21812 11392 21828 11456
rect 21892 11392 21908 11456
rect 21972 11392 21980 11456
rect 21660 10368 21980 11392
rect 21660 10304 21668 10368
rect 21732 10304 21748 10368
rect 21812 10304 21828 10368
rect 21892 10304 21908 10368
rect 21972 10304 21980 10368
rect 21660 9280 21980 10304
rect 21660 9216 21668 9280
rect 21732 9216 21748 9280
rect 21812 9216 21828 9280
rect 21892 9216 21908 9280
rect 21972 9216 21980 9280
rect 21660 8192 21980 9216
rect 21660 8128 21668 8192
rect 21732 8128 21748 8192
rect 21812 8128 21828 8192
rect 21892 8128 21908 8192
rect 21972 8128 21980 8192
rect 21660 7104 21980 8128
rect 21660 7040 21668 7104
rect 21732 7040 21748 7104
rect 21812 7040 21828 7104
rect 21892 7040 21908 7104
rect 21972 7040 21980 7104
rect 21660 6016 21980 7040
rect 21660 5952 21668 6016
rect 21732 5952 21748 6016
rect 21812 5952 21828 6016
rect 21892 5952 21908 6016
rect 21972 5952 21980 6016
rect 21660 4928 21980 5952
rect 21660 4864 21668 4928
rect 21732 4864 21748 4928
rect 21812 4864 21828 4928
rect 21892 4864 21908 4928
rect 21972 4864 21980 4928
rect 21660 3840 21980 4864
rect 21660 3776 21668 3840
rect 21732 3776 21748 3840
rect 21812 3776 21828 3840
rect 21892 3776 21908 3840
rect 21972 3776 21980 3840
rect 21660 2752 21980 3776
rect 21660 2688 21668 2752
rect 21732 2688 21748 2752
rect 21812 2688 21828 2752
rect 21892 2688 21908 2752
rect 21972 2688 21980 2752
rect 21660 2672 21980 2688
rect 28360 10912 28680 11936
rect 28360 10848 28368 10912
rect 28432 10848 28448 10912
rect 28512 10848 28528 10912
rect 28592 10848 28608 10912
rect 28672 10848 28680 10912
rect 28360 9824 28680 10848
rect 28360 9760 28368 9824
rect 28432 9760 28448 9824
rect 28512 9760 28528 9824
rect 28592 9760 28608 9824
rect 28672 9760 28680 9824
rect 28360 8736 28680 9760
rect 28360 8672 28368 8736
rect 28432 8672 28448 8736
rect 28512 8672 28528 8736
rect 28592 8672 28608 8736
rect 28672 8672 28680 8736
rect 28360 7648 28680 8672
rect 28360 7584 28368 7648
rect 28432 7584 28448 7648
rect 28512 7584 28528 7648
rect 28592 7584 28608 7648
rect 28672 7584 28680 7648
rect 28360 6560 28680 7584
rect 28360 6496 28368 6560
rect 28432 6496 28448 6560
rect 28512 6496 28528 6560
rect 28592 6496 28608 6560
rect 28672 6496 28680 6560
rect 28360 5472 28680 6496
rect 28360 5408 28368 5472
rect 28432 5408 28448 5472
rect 28512 5408 28528 5472
rect 28592 5408 28608 5472
rect 28672 5408 28680 5472
rect 28360 4384 28680 5408
rect 28360 4320 28368 4384
rect 28432 4320 28448 4384
rect 28512 4320 28528 4384
rect 28592 4320 28608 4384
rect 28672 4320 28680 4384
rect 28360 3296 28680 4320
rect 28360 3232 28368 3296
rect 28432 3232 28448 3296
rect 28512 3232 28528 3296
rect 28592 3232 28608 3296
rect 28672 3232 28680 3296
rect 28360 2672 28680 3232
rect 29020 32128 29340 32144
rect 29020 32064 29028 32128
rect 29092 32064 29108 32128
rect 29172 32064 29188 32128
rect 29252 32064 29268 32128
rect 29332 32064 29340 32128
rect 29020 31040 29340 32064
rect 29020 30976 29028 31040
rect 29092 30976 29108 31040
rect 29172 30976 29188 31040
rect 29252 30976 29268 31040
rect 29332 30976 29340 31040
rect 29020 29952 29340 30976
rect 29020 29888 29028 29952
rect 29092 29888 29108 29952
rect 29172 29888 29188 29952
rect 29252 29888 29268 29952
rect 29332 29888 29340 29952
rect 29020 28864 29340 29888
rect 29020 28800 29028 28864
rect 29092 28800 29108 28864
rect 29172 28800 29188 28864
rect 29252 28800 29268 28864
rect 29332 28800 29340 28864
rect 29020 27776 29340 28800
rect 29020 27712 29028 27776
rect 29092 27712 29108 27776
rect 29172 27712 29188 27776
rect 29252 27712 29268 27776
rect 29332 27712 29340 27776
rect 29020 26688 29340 27712
rect 29020 26624 29028 26688
rect 29092 26624 29108 26688
rect 29172 26624 29188 26688
rect 29252 26624 29268 26688
rect 29332 26624 29340 26688
rect 29020 25600 29340 26624
rect 29020 25536 29028 25600
rect 29092 25536 29108 25600
rect 29172 25536 29188 25600
rect 29252 25536 29268 25600
rect 29332 25536 29340 25600
rect 29020 24512 29340 25536
rect 29020 24448 29028 24512
rect 29092 24448 29108 24512
rect 29172 24448 29188 24512
rect 29252 24448 29268 24512
rect 29332 24448 29340 24512
rect 29020 23424 29340 24448
rect 29020 23360 29028 23424
rect 29092 23360 29108 23424
rect 29172 23360 29188 23424
rect 29252 23360 29268 23424
rect 29332 23360 29340 23424
rect 29020 22336 29340 23360
rect 29020 22272 29028 22336
rect 29092 22272 29108 22336
rect 29172 22272 29188 22336
rect 29252 22272 29268 22336
rect 29332 22272 29340 22336
rect 29020 21248 29340 22272
rect 29020 21184 29028 21248
rect 29092 21184 29108 21248
rect 29172 21184 29188 21248
rect 29252 21184 29268 21248
rect 29332 21184 29340 21248
rect 29020 20160 29340 21184
rect 29020 20096 29028 20160
rect 29092 20096 29108 20160
rect 29172 20096 29188 20160
rect 29252 20096 29268 20160
rect 29332 20096 29340 20160
rect 29020 19072 29340 20096
rect 29020 19008 29028 19072
rect 29092 19008 29108 19072
rect 29172 19008 29188 19072
rect 29252 19008 29268 19072
rect 29332 19008 29340 19072
rect 29020 17984 29340 19008
rect 29020 17920 29028 17984
rect 29092 17920 29108 17984
rect 29172 17920 29188 17984
rect 29252 17920 29268 17984
rect 29332 17920 29340 17984
rect 29020 16896 29340 17920
rect 29020 16832 29028 16896
rect 29092 16832 29108 16896
rect 29172 16832 29188 16896
rect 29252 16832 29268 16896
rect 29332 16832 29340 16896
rect 29020 15808 29340 16832
rect 29020 15744 29028 15808
rect 29092 15744 29108 15808
rect 29172 15744 29188 15808
rect 29252 15744 29268 15808
rect 29332 15744 29340 15808
rect 29020 14720 29340 15744
rect 29020 14656 29028 14720
rect 29092 14656 29108 14720
rect 29172 14656 29188 14720
rect 29252 14656 29268 14720
rect 29332 14656 29340 14720
rect 29020 13632 29340 14656
rect 29020 13568 29028 13632
rect 29092 13568 29108 13632
rect 29172 13568 29188 13632
rect 29252 13568 29268 13632
rect 29332 13568 29340 13632
rect 29020 12544 29340 13568
rect 29020 12480 29028 12544
rect 29092 12480 29108 12544
rect 29172 12480 29188 12544
rect 29252 12480 29268 12544
rect 29332 12480 29340 12544
rect 29020 11456 29340 12480
rect 29020 11392 29028 11456
rect 29092 11392 29108 11456
rect 29172 11392 29188 11456
rect 29252 11392 29268 11456
rect 29332 11392 29340 11456
rect 29020 10368 29340 11392
rect 29020 10304 29028 10368
rect 29092 10304 29108 10368
rect 29172 10304 29188 10368
rect 29252 10304 29268 10368
rect 29332 10304 29340 10368
rect 29020 9280 29340 10304
rect 29020 9216 29028 9280
rect 29092 9216 29108 9280
rect 29172 9216 29188 9280
rect 29252 9216 29268 9280
rect 29332 9216 29340 9280
rect 29020 8192 29340 9216
rect 29020 8128 29028 8192
rect 29092 8128 29108 8192
rect 29172 8128 29188 8192
rect 29252 8128 29268 8192
rect 29332 8128 29340 8192
rect 29020 7104 29340 8128
rect 29020 7040 29028 7104
rect 29092 7040 29108 7104
rect 29172 7040 29188 7104
rect 29252 7040 29268 7104
rect 29332 7040 29340 7104
rect 29020 6016 29340 7040
rect 29020 5952 29028 6016
rect 29092 5952 29108 6016
rect 29172 5952 29188 6016
rect 29252 5952 29268 6016
rect 29332 5952 29340 6016
rect 29020 4928 29340 5952
rect 29020 4864 29028 4928
rect 29092 4864 29108 4928
rect 29172 4864 29188 4928
rect 29252 4864 29268 4928
rect 29332 4864 29340 4928
rect 29020 3840 29340 4864
rect 29020 3776 29028 3840
rect 29092 3776 29108 3840
rect 29172 3776 29188 3840
rect 29252 3776 29268 3840
rect 29332 3776 29340 3840
rect 29020 2752 29340 3776
rect 29020 2688 29028 2752
rect 29092 2688 29108 2752
rect 29172 2688 29188 2752
rect 29252 2688 29268 2752
rect 29332 2688 29340 2752
rect 29020 2672 29340 2688
use sky130_fd_sc_hd__inv_2  _0617_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31648 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0618_
timestamp 1688980957
transform 1 0 14076 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0619_
timestamp 1688980957
transform 1 0 23644 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0620_
timestamp 1688980957
transform -1 0 26128 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0621_
timestamp 1688980957
transform 1 0 26036 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0622_
timestamp 1688980957
transform -1 0 23736 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0623_
timestamp 1688980957
transform 1 0 29532 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0624_
timestamp 1688980957
transform 1 0 16192 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0625_
timestamp 1688980957
transform -1 0 12052 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0626_
timestamp 1688980957
transform -1 0 12972 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0627_
timestamp 1688980957
transform -1 0 18032 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0628_
timestamp 1688980957
transform -1 0 22816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0629_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23368 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0630_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24564 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _0631_
timestamp 1688980957
transform 1 0 22908 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0632_
timestamp 1688980957
transform -1 0 27692 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0633_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0634_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26864 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0635_
timestamp 1688980957
transform 1 0 23460 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0636_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29808 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0637_
timestamp 1688980957
transform 1 0 25392 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _0638_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26496 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0639_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26588 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0640_
timestamp 1688980957
transform -1 0 27968 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__or4bb_1  _0641_
timestamp 1688980957
transform 1 0 24472 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0642_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25576 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_4  _0643_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26312 0 -1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__o31a_1  _0644_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0645_
timestamp 1688980957
transform -1 0 24472 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0646_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24288 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0647_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24288 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0648_
timestamp 1688980957
transform 1 0 24196 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0649_
timestamp 1688980957
transform -1 0 24840 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0650_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24380 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1688980957
transform -1 0 26496 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0652_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28428 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0653_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25944 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0654_
timestamp 1688980957
transform 1 0 25392 0 -1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0655_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22724 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0656_
timestamp 1688980957
transform -1 0 24656 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0657_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26680 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0658_
timestamp 1688980957
transform 1 0 22356 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _0659_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25116 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _0660_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25760 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0661_
timestamp 1688980957
transform 1 0 23920 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0662_
timestamp 1688980957
transform -1 0 22724 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0663_
timestamp 1688980957
transform 1 0 23092 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0664_
timestamp 1688980957
transform -1 0 28336 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0665_
timestamp 1688980957
transform 1 0 27508 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o41a_1  _0666_
timestamp 1688980957
transform 1 0 23552 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0667_
timestamp 1688980957
transform 1 0 23460 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _0668_
timestamp 1688980957
transform -1 0 25024 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0669_
timestamp 1688980957
transform -1 0 22540 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0670_
timestamp 1688980957
transform 1 0 21712 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0671_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21436 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _0672_
timestamp 1688980957
transform -1 0 30360 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__or4bb_1  _0673_
timestamp 1688980957
transform 1 0 27692 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0674_
timestamp 1688980957
transform 1 0 27692 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0675_
timestamp 1688980957
transform 1 0 27048 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor4_1  _0676_
timestamp 1688980957
transform 1 0 27508 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0677_
timestamp 1688980957
transform -1 0 24288 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0678_
timestamp 1688980957
transform -1 0 24656 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0679_
timestamp 1688980957
transform -1 0 20792 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _0680_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23644 0 1 13600
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_1  _0681_
timestamp 1688980957
transform 1 0 27968 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0682_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28428 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0683_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29256 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0684_
timestamp 1688980957
transform -1 0 26496 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0685_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25024 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _0686_
timestamp 1688980957
transform -1 0 23184 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0687_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24012 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0688_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20792 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0689_
timestamp 1688980957
transform 1 0 24564 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0690_
timestamp 1688980957
transform -1 0 25668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0691_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0692_
timestamp 1688980957
transform 1 0 22264 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and4_2  _0693_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27876 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0694_
timestamp 1688980957
transform 1 0 25116 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 1688980957
transform 1 0 24932 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0696_
timestamp 1688980957
transform -1 0 27784 0 -1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1688980957
transform 1 0 26588 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0698_
timestamp 1688980957
transform -1 0 28244 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0699_
timestamp 1688980957
transform 1 0 27968 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0700_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29716 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0701_
timestamp 1688980957
transform -1 0 29532 0 1 10336
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0702_
timestamp 1688980957
transform -1 0 30176 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _0703_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24932 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  _0704_
timestamp 1688980957
transform -1 0 23920 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a41oi_2  _0705_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29072 0 -1 12512
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _0706_
timestamp 1688980957
transform 1 0 30452 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0707_
timestamp 1688980957
transform -1 0 31648 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0708_
timestamp 1688980957
transform -1 0 29256 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_1  _0709_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29072 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0710_
timestamp 1688980957
transform 1 0 30820 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0711_
timestamp 1688980957
transform -1 0 30360 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0712_
timestamp 1688980957
transform 1 0 31464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0713_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28704 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0714_
timestamp 1688980957
transform 1 0 27140 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0715_
timestamp 1688980957
transform 1 0 28612 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0716_
timestamp 1688980957
transform 1 0 30820 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0717_
timestamp 1688980957
transform 1 0 30544 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0718_
timestamp 1688980957
transform -1 0 30544 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0719_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28612 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0720_
timestamp 1688980957
transform -1 0 29072 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0721_
timestamp 1688980957
transform -1 0 30084 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0722_
timestamp 1688980957
transform -1 0 28520 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_1  _0723_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28980 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0724_
timestamp 1688980957
transform 1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0725_
timestamp 1688980957
transform -1 0 28060 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0726_
timestamp 1688980957
transform -1 0 25944 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0727_
timestamp 1688980957
transform 1 0 26772 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0728_
timestamp 1688980957
transform 1 0 26036 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0729_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27508 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0730_
timestamp 1688980957
transform 1 0 27416 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0731_
timestamp 1688980957
transform -1 0 26220 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0732_
timestamp 1688980957
transform -1 0 27324 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0733_
timestamp 1688980957
transform -1 0 29072 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1688980957
transform 1 0 29072 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0735_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0736_
timestamp 1688980957
transform 1 0 27876 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0737_
timestamp 1688980957
transform -1 0 26128 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0738_
timestamp 1688980957
transform -1 0 29072 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0739_
timestamp 1688980957
transform -1 0 26312 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0740_
timestamp 1688980957
transform 1 0 26312 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0741_
timestamp 1688980957
transform -1 0 28336 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0742_
timestamp 1688980957
transform -1 0 28152 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0743_
timestamp 1688980957
transform 1 0 25944 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0744_
timestamp 1688980957
transform 1 0 21252 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0745_
timestamp 1688980957
transform 1 0 22080 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0746_
timestamp 1688980957
transform -1 0 21712 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0747_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23552 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0748_
timestamp 1688980957
transform 1 0 23460 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0749_
timestamp 1688980957
transform -1 0 22724 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0750_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19136 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _0751_
timestamp 1688980957
transform 1 0 21620 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0752_
timestamp 1688980957
transform 1 0 22724 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0753_
timestamp 1688980957
transform 1 0 23092 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0754_
timestamp 1688980957
transform 1 0 24288 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0755_
timestamp 1688980957
transform -1 0 24288 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0756_
timestamp 1688980957
transform 1 0 17204 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0757_
timestamp 1688980957
transform 1 0 17204 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0758_
timestamp 1688980957
transform -1 0 23000 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0759_
timestamp 1688980957
transform 1 0 16836 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0760_
timestamp 1688980957
transform 1 0 18860 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0761_
timestamp 1688980957
transform 1 0 19780 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0762_
timestamp 1688980957
transform 1 0 20884 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__and2_2  _0763_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27692 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _0764_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27140 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1688980957
transform -1 0 19780 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0766_
timestamp 1688980957
transform -1 0 26404 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0767_
timestamp 1688980957
transform 1 0 20884 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0768_
timestamp 1688980957
transform -1 0 21804 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0769_
timestamp 1688980957
transform -1 0 29440 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0770_
timestamp 1688980957
transform -1 0 20148 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0771_
timestamp 1688980957
transform -1 0 27416 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0772_
timestamp 1688980957
transform 1 0 19964 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0773_
timestamp 1688980957
transform -1 0 20424 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_2  _0774_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29532 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _0775_
timestamp 1688980957
transform -1 0 27876 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0776_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27140 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _0777_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25944 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0778_
timestamp 1688980957
transform -1 0 24380 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _0779_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26036 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0780_
timestamp 1688980957
transform -1 0 28244 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0781_
timestamp 1688980957
transform -1 0 25852 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0782_
timestamp 1688980957
transform 1 0 26864 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0783_
timestamp 1688980957
transform -1 0 24748 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0784_
timestamp 1688980957
transform 1 0 24840 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0785_
timestamp 1688980957
transform -1 0 24840 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0786_
timestamp 1688980957
transform -1 0 28336 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0787_
timestamp 1688980957
transform 1 0 30452 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0788_
timestamp 1688980957
transform -1 0 31188 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0789_
timestamp 1688980957
transform -1 0 29256 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1688980957
transform -1 0 28152 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0791_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27416 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0792_
timestamp 1688980957
transform -1 0 25116 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0793_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23000 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0794_
timestamp 1688980957
transform 1 0 24932 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0795_
timestamp 1688980957
transform 1 0 23552 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0796_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27876 0 -1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0797_
timestamp 1688980957
transform -1 0 24012 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0798_
timestamp 1688980957
transform 1 0 24196 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0799_
timestamp 1688980957
transform 1 0 25576 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0800_
timestamp 1688980957
transform 1 0 25392 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0801_
timestamp 1688980957
transform -1 0 24840 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0802_
timestamp 1688980957
transform 1 0 26036 0 -1 31008
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0803_
timestamp 1688980957
transform -1 0 26956 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0804_
timestamp 1688980957
transform -1 0 26772 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0805_
timestamp 1688980957
transform -1 0 28336 0 1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _0806_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29348 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0807_
timestamp 1688980957
transform -1 0 28796 0 1 28832
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0808_
timestamp 1688980957
transform -1 0 25944 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1688980957
transform 1 0 29808 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _0810_
timestamp 1688980957
transform 1 0 28796 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0811_
timestamp 1688980957
transform 1 0 30636 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0812_
timestamp 1688980957
transform 1 0 31096 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0813_
timestamp 1688980957
transform 1 0 27140 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0814_
timestamp 1688980957
transform -1 0 30544 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0815_
timestamp 1688980957
transform -1 0 28888 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1688980957
transform -1 0 29716 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _0817_
timestamp 1688980957
transform -1 0 28244 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0818_
timestamp 1688980957
transform -1 0 28520 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0819_
timestamp 1688980957
transform 1 0 28244 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0820_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27784 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0821_
timestamp 1688980957
transform -1 0 27416 0 1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0822_
timestamp 1688980957
transform 1 0 26220 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0823_
timestamp 1688980957
transform 1 0 24932 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0824_
timestamp 1688980957
transform -1 0 25944 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _0825_
timestamp 1688980957
transform 1 0 24932 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0826_
timestamp 1688980957
transform 1 0 24288 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0827_
timestamp 1688980957
transform 1 0 23460 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0828_
timestamp 1688980957
transform 1 0 23000 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0829_
timestamp 1688980957
transform -1 0 21988 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0830_
timestamp 1688980957
transform 1 0 23184 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0831_
timestamp 1688980957
transform 1 0 14720 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0832_
timestamp 1688980957
transform -1 0 14720 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _0833_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0834_
timestamp 1688980957
transform 1 0 14260 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _0835_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21344 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0836_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17480 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_2  _0837_
timestamp 1688980957
transform 1 0 17204 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_4  _0838_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2b_1  _0839_
timestamp 1688980957
transform 1 0 12236 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__or2_4  _0840_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12236 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _0841_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0842_
timestamp 1688980957
transform -1 0 14168 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_4  _0843_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 17952
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _0844_
timestamp 1688980957
transform -1 0 19504 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_2  _0845_
timestamp 1688980957
transform 1 0 14904 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _0846_
timestamp 1688980957
transform -1 0 13800 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0847_
timestamp 1688980957
transform 1 0 14352 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _0848_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 -1 16864
box -38 -48 958 592
use sky130_fd_sc_hd__nor3_1  _0849_
timestamp 1688980957
transform 1 0 14076 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _0850_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17388 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0851_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0852_
timestamp 1688980957
transform 1 0 13524 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0853_
timestamp 1688980957
transform 1 0 9844 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _0854_
timestamp 1688980957
transform 1 0 11960 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0855_
timestamp 1688980957
transform -1 0 12328 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0856_
timestamp 1688980957
transform 1 0 13156 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0857_
timestamp 1688980957
transform -1 0 13524 0 1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0858_
timestamp 1688980957
transform -1 0 16468 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0859_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12880 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _0860_
timestamp 1688980957
transform 1 0 8924 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _0861_
timestamp 1688980957
transform -1 0 13800 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0862_
timestamp 1688980957
transform -1 0 15364 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0863_
timestamp 1688980957
transform -1 0 14628 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0864_
timestamp 1688980957
transform 1 0 13524 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0865_
timestamp 1688980957
transform 1 0 14996 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0866_
timestamp 1688980957
transform 1 0 13984 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 1688980957
transform 1 0 13156 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0868_
timestamp 1688980957
transform -1 0 15088 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _0869_
timestamp 1688980957
transform -1 0 13064 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0870_
timestamp 1688980957
transform 1 0 12420 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _0871_
timestamp 1688980957
transform 1 0 13984 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_2  _0872_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16744 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__a2111oi_4  _0873_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 -1 15776
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _0874_
timestamp 1688980957
transform 1 0 13984 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0875_
timestamp 1688980957
transform -1 0 12696 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0876_
timestamp 1688980957
transform -1 0 11776 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0877_
timestamp 1688980957
transform 1 0 11316 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0878_
timestamp 1688980957
transform 1 0 11684 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0879_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11316 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0880_
timestamp 1688980957
transform -1 0 11408 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0881_
timestamp 1688980957
transform 1 0 12420 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0882_
timestamp 1688980957
transform -1 0 12604 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0883_
timestamp 1688980957
transform -1 0 15916 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0884_
timestamp 1688980957
transform 1 0 13156 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0885_
timestamp 1688980957
transform -1 0 13708 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0886_
timestamp 1688980957
transform 1 0 14168 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0887_
timestamp 1688980957
transform -1 0 14996 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0888_
timestamp 1688980957
transform 1 0 14996 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _0889_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _0890_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0891_
timestamp 1688980957
transform -1 0 14720 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0892_
timestamp 1688980957
transform 1 0 15364 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0893_
timestamp 1688980957
transform 1 0 14352 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0894_
timestamp 1688980957
transform -1 0 11868 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0895_
timestamp 1688980957
transform 1 0 11868 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0896_
timestamp 1688980957
transform -1 0 11316 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0897_
timestamp 1688980957
transform -1 0 10212 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0898_
timestamp 1688980957
transform -1 0 11960 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0899_
timestamp 1688980957
transform 1 0 9844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0900_
timestamp 1688980957
transform 1 0 14260 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0901_
timestamp 1688980957
transform 1 0 14904 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0902_
timestamp 1688980957
transform 1 0 12420 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0903_
timestamp 1688980957
transform 1 0 13984 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0904_
timestamp 1688980957
transform -1 0 11224 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0905_
timestamp 1688980957
transform 1 0 10672 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0906_
timestamp 1688980957
transform -1 0 15364 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0907_
timestamp 1688980957
transform 1 0 13708 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_4  _0908_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10856 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0909_
timestamp 1688980957
transform -1 0 7544 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0910_
timestamp 1688980957
transform -1 0 13800 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0911_
timestamp 1688980957
transform -1 0 10028 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0912_
timestamp 1688980957
transform -1 0 6072 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0913_
timestamp 1688980957
transform 1 0 6256 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0914_
timestamp 1688980957
transform 1 0 18308 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0915_
timestamp 1688980957
transform -1 0 9476 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0916_
timestamp 1688980957
transform 1 0 18124 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0917_
timestamp 1688980957
transform -1 0 12604 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0918_
timestamp 1688980957
transform -1 0 10212 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0919_
timestamp 1688980957
transform -1 0 10856 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0920_
timestamp 1688980957
transform -1 0 7084 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0921_
timestamp 1688980957
transform 1 0 10304 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0922_
timestamp 1688980957
transform 1 0 17296 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0923_
timestamp 1688980957
transform 1 0 10212 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0924_
timestamp 1688980957
transform -1 0 11316 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1688980957
transform -1 0 15548 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0926_
timestamp 1688980957
transform 1 0 15732 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 1688980957
transform -1 0 12144 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0928_
timestamp 1688980957
transform -1 0 9384 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0929_
timestamp 1688980957
transform -1 0 10948 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0930_
timestamp 1688980957
transform -1 0 11224 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0931_
timestamp 1688980957
transform 1 0 14720 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0932_
timestamp 1688980957
transform -1 0 8372 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_4  _0933_
timestamp 1688980957
transform 1 0 10856 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0934_
timestamp 1688980957
transform -1 0 11960 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0935_
timestamp 1688980957
transform -1 0 6164 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0936_
timestamp 1688980957
transform -1 0 7176 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0937_
timestamp 1688980957
transform -1 0 7360 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0938_
timestamp 1688980957
transform 1 0 16836 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0939_
timestamp 1688980957
transform -1 0 13800 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0940_
timestamp 1688980957
transform -1 0 17480 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0941_
timestamp 1688980957
transform -1 0 18952 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0942_
timestamp 1688980957
transform -1 0 8648 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0943_
timestamp 1688980957
transform -1 0 9476 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0944_
timestamp 1688980957
transform 1 0 17204 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0945_
timestamp 1688980957
transform -1 0 8924 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0946_
timestamp 1688980957
transform 1 0 14996 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0947_
timestamp 1688980957
transform -1 0 10028 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0948_
timestamp 1688980957
transform 1 0 11316 0 -1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0949_
timestamp 1688980957
transform 1 0 14352 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0950_
timestamp 1688980957
transform 1 0 8096 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0951_
timestamp 1688980957
transform 1 0 7268 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0952_
timestamp 1688980957
transform 1 0 9292 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0953_
timestamp 1688980957
transform 1 0 8740 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0954_
timestamp 1688980957
transform 1 0 10120 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0955_
timestamp 1688980957
transform 1 0 11960 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0956_
timestamp 1688980957
transform 1 0 10580 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0957_
timestamp 1688980957
transform -1 0 13984 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0958_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16836 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__nor3_4  _0959_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13984 0 1 14688
box -38 -48 1234 592
use sky130_fd_sc_hd__mux4_1  _0960_
timestamp 1688980957
transform -1 0 31924 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0961_
timestamp 1688980957
transform -1 0 23184 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0962_
timestamp 1688980957
transform 1 0 21988 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0963_
timestamp 1688980957
transform 1 0 13616 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0964_
timestamp 1688980957
transform 1 0 14996 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0965_
timestamp 1688980957
transform 1 0 16468 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0966_
timestamp 1688980957
transform -1 0 14812 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0967_
timestamp 1688980957
transform 1 0 13984 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0968_
timestamp 1688980957
transform -1 0 14996 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0969_
timestamp 1688980957
transform -1 0 31924 0 -1 20128
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0970_
timestamp 1688980957
transform 1 0 22540 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0971_
timestamp 1688980957
transform 1 0 24196 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0972_
timestamp 1688980957
transform 1 0 10672 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0973_
timestamp 1688980957
transform 1 0 14168 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0974_
timestamp 1688980957
transform 1 0 14996 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0975_
timestamp 1688980957
transform 1 0 13156 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0976_
timestamp 1688980957
transform 1 0 15732 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0977_
timestamp 1688980957
transform 1 0 15732 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0978_
timestamp 1688980957
transform -1 0 19320 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0979_
timestamp 1688980957
transform -1 0 21528 0 1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0980_
timestamp 1688980957
transform 1 0 20240 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _0981_
timestamp 1688980957
transform 1 0 18400 0 -1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__and3b_1  _0982_
timestamp 1688980957
transform 1 0 19412 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0983_
timestamp 1688980957
transform 1 0 20884 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0984_
timestamp 1688980957
transform 1 0 15824 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 1688980957
transform -1 0 20332 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0986_
timestamp 1688980957
transform 1 0 19044 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0987_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17112 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0988_
timestamp 1688980957
transform 1 0 16836 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0989_
timestamp 1688980957
transform -1 0 12880 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0990_
timestamp 1688980957
transform 1 0 29348 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0991_
timestamp 1688980957
transform 1 0 4416 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0992_
timestamp 1688980957
transform 1 0 6440 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0993_
timestamp 1688980957
transform 1 0 29532 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0994_
timestamp 1688980957
transform 1 0 5428 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0995_
timestamp 1688980957
transform 1 0 28612 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0996_
timestamp 1688980957
transform 1 0 20884 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0997_
timestamp 1688980957
transform 1 0 14352 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1688980957
transform 1 0 16008 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 1688980957
transform 1 0 13524 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1000_
timestamp 1688980957
transform -1 0 6256 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1001_
timestamp 1688980957
transform 1 0 5704 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1002_
timestamp 1688980957
transform -1 0 18124 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1003_
timestamp 1688980957
transform -1 0 17296 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1004_
timestamp 1688980957
transform 1 0 11040 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 1688980957
transform 1 0 14628 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1006_
timestamp 1688980957
transform -1 0 6440 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1007_
timestamp 1688980957
transform 1 0 13800 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1008_
timestamp 1688980957
transform -1 0 11776 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1009_
timestamp 1688980957
transform -1 0 4968 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1010_
timestamp 1688980957
transform -1 0 6256 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1011_
timestamp 1688980957
transform -1 0 24748 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1012_
timestamp 1688980957
transform 1 0 8004 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1013_
timestamp 1688980957
transform 1 0 20976 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1688980957
transform 1 0 8004 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1015_
timestamp 1688980957
transform -1 0 5336 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1016_
timestamp 1688980957
transform 1 0 19688 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1017_
timestamp 1688980957
transform 1 0 14628 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1018_
timestamp 1688980957
transform 1 0 16928 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1688980957
transform 1 0 9384 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1020_
timestamp 1688980957
transform 1 0 3404 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1021_
timestamp 1688980957
transform 1 0 6532 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__o2bb2a_1  _1022_
timestamp 1688980957
transform 1 0 15824 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1023_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1024_
timestamp 1688980957
transform -1 0 18216 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and4_4  _1025_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17204 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp 1688980957
transform -1 0 12880 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1027_
timestamp 1688980957
transform 1 0 4692 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1688980957
transform -1 0 6256 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1029_
timestamp 1688980957
transform -1 0 6624 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1030_
timestamp 1688980957
transform 1 0 18584 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1031_
timestamp 1688980957
transform 1 0 13432 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1032_
timestamp 1688980957
transform -1 0 19596 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1033_
timestamp 1688980957
transform -1 0 19780 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1034_
timestamp 1688980957
transform 1 0 5428 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1035_
timestamp 1688980957
transform 1 0 8004 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1036_
timestamp 1688980957
transform 1 0 19780 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1037_
timestamp 1688980957
transform 1 0 8464 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1038_
timestamp 1688980957
transform 1 0 18860 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1039_
timestamp 1688980957
transform 1 0 8004 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1040_
timestamp 1688980957
transform 1 0 19504 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1041_
timestamp 1688980957
transform 1 0 15732 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1042_
timestamp 1688980957
transform 1 0 18308 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1043_
timestamp 1688980957
transform 1 0 17296 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1044_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22724 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1045_
timestamp 1688980957
transform 1 0 21988 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1046_
timestamp 1688980957
transform 1 0 28888 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1047_
timestamp 1688980957
transform 1 0 28704 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1048_
timestamp 1688980957
transform 1 0 22816 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1049_
timestamp 1688980957
transform -1 0 18584 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1050_
timestamp 1688980957
transform 1 0 19136 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1051_
timestamp 1688980957
transform 1 0 15916 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1052_
timestamp 1688980957
transform -1 0 21620 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1688980957
transform -1 0 7912 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1054_
timestamp 1688980957
transform -1 0 18124 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1055_
timestamp 1688980957
transform 1 0 7544 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1056_
timestamp 1688980957
transform -1 0 19228 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1688980957
transform -1 0 6900 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1058_
timestamp 1688980957
transform -1 0 6532 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1059_
timestamp 1688980957
transform -1 0 21896 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1688980957
transform 1 0 18860 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1061_
timestamp 1688980957
transform -1 0 15272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1688980957
transform -1 0 20332 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1063_
timestamp 1688980957
transform -1 0 5244 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1064_
timestamp 1688980957
transform -1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1065_
timestamp 1688980957
transform -1 0 6440 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1066_
timestamp 1688980957
transform -1 0 12788 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1688980957
transform -1 0 7636 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1688980957
transform -1 0 5244 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1688980957
transform 1 0 9660 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1688980957
transform 1 0 18308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1688980957
transform 1 0 12788 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1688980957
transform 1 0 20424 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1688980957
transform -1 0 5704 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1688980957
transform 1 0 8188 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1688980957
transform 1 0 21804 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1688980957
transform 1 0 7636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1688980957
transform -1 0 25668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1688980957
transform -1 0 6900 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1688980957
transform -1 0 5244 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1688980957
transform -1 0 12696 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1688980957
transform -1 0 16008 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1688980957
transform -1 0 7544 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1688980957
transform -1 0 16284 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1688980957
transform -1 0 12144 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1688980957
transform -1 0 19320 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1086_
timestamp 1688980957
transform -1 0 19320 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1688980957
transform -1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1688980957
transform -1 0 6348 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1688980957
transform -1 0 15456 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1688980957
transform 1 0 16836 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1688980957
transform -1 0 13892 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1688980957
transform 1 0 21252 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1688980957
transform -1 0 30176 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1688980957
transform -1 0 5244 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1688980957
transform 1 0 31188 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1688980957
transform 1 0 6440 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1688980957
transform -1 0 5612 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1688980957
transform 1 0 30176 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1688980957
transform 1 0 17848 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1688980957
transform -1 0 20608 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1688980957
transform -1 0 21620 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1688980957
transform -1 0 16284 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1688980957
transform -1 0 16744 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1688980957
transform -1 0 23736 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1688980957
transform -1 0 16744 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1106_
timestamp 1688980957
transform -1 0 17296 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1688980957
transform -1 0 23276 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1688980957
transform -1 0 13064 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1688980957
transform -1 0 10120 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1688980957
transform 1 0 11684 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1688980957
transform 1 0 10672 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1688980957
transform 1 0 9016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1688980957
transform 1 0 8740 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1688980957
transform -1 0 8372 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1688980957
transform 1 0 8464 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1688980957
transform -1 0 16744 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1688980957
transform -1 0 13432 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1688980957
transform -1 0 10304 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1688980957
transform 1 0 15732 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1688980957
transform 1 0 8004 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1688980957
transform -1 0 18584 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1688980957
transform -1 0 7912 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1688980957
transform 1 0 6992 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1688980957
transform -1 0 19228 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1688980957
transform -1 0 18124 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1688980957
transform -1 0 14168 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1688980957
transform 1 0 18584 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1688980957
transform -1 0 6440 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1688980957
transform 1 0 5704 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1688980957
transform -1 0 5888 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1688980957
transform -1 0 12236 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1688980957
transform -1 0 10212 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1688980957
transform 1 0 10212 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1134_
timestamp 1688980957
transform -1 0 10488 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1688980957
transform 1 0 18124 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1688980957
transform -1 0 12972 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1688980957
transform -1 0 19780 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1688980957
transform -1 0 9844 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1688980957
transform 1 0 7636 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1688980957
transform -1 0 21436 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1688980957
transform 1 0 7820 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1688980957
transform -1 0 18216 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 1688980957
transform -1 0 7360 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1688980957
transform 1 0 5704 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1688980957
transform -1 0 10304 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1688980957
transform 1 0 13432 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1688980957
transform -1 0 8280 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1688980957
transform 1 0 13984 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1149_
timestamp 1688980957
transform -1 0 10488 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1688980957
transform -1 0 16376 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1688980957
transform -1 0 16100 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1688980957
transform -1 0 9936 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1153_
timestamp 1688980957
transform -1 0 10304 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1154_
timestamp 1688980957
transform -1 0 13432 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1155_
timestamp 1688980957
transform -1 0 16008 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 1688980957
transform -1 0 15548 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1688980957
transform -1 0 14260 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1158_
timestamp 1688980957
transform -1 0 12972 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1159_
timestamp 1688980957
transform 1 0 10580 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1688980957
transform 1 0 12052 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1688980957
transform -1 0 14076 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1688980957
transform -1 0 17112 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1163_
timestamp 1688980957
transform -1 0 30360 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1688980957
transform -1 0 29992 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1688980957
transform 1 0 21988 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1688980957
transform 1 0 22356 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1167_
timestamp 1688980957
transform -1 0 23460 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1688980957
transform 1 0 25576 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1688980957
transform -1 0 28888 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1688980957
transform -1 0 28888 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1171_
timestamp 1688980957
transform -1 0 30360 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1688980957
transform -1 0 31004 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1688980957
transform -1 0 31004 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1174_
timestamp 1688980957
transform -1 0 31464 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1688980957
transform -1 0 31096 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1176_
timestamp 1688980957
transform -1 0 28888 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1177_
timestamp 1688980957
transform 1 0 25668 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1688980957
transform -1 0 25668 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1688980957
transform 1 0 22632 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1688980957
transform 1 0 22540 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1688980957
transform -1 0 28796 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1688980957
transform -1 0 28520 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1688980957
transform -1 0 25208 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1688980957
transform 1 0 23000 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1688980957
transform -1 0 19964 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1688980957
transform -1 0 21712 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1688980957
transform -1 0 28428 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1688980957
transform 1 0 19044 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1688980957
transform -1 0 29716 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190_
timestamp 1688980957
transform -1 0 21160 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1688980957
transform -1 0 20516 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1688980957
transform -1 0 27508 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1688980957
transform -1 0 20056 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1194_
timestamp 1688980957
transform -1 0 21988 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1195_
timestamp 1688980957
transform -1 0 21160 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1196_
timestamp 1688980957
transform -1 0 18584 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1197_
timestamp 1688980957
transform -1 0 18584 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198_
timestamp 1688980957
transform -1 0 24012 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1199_
timestamp 1688980957
transform -1 0 18584 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1688980957
transform -1 0 18584 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1688980957
transform -1 0 23736 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1688980957
transform 1 0 25116 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1688980957
transform 1 0 28888 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1688980957
transform -1 0 24196 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1688980957
transform 1 0 24380 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1688980957
transform -1 0 28612 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1207_
timestamp 1688980957
transform -1 0 28428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1688980957
transform 1 0 25668 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 1688980957
transform 1 0 25668 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1688980957
transform 1 0 25668 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1688980957
transform 1 0 26312 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1212_
timestamp 1688980957
transform -1 0 25944 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1213_
timestamp 1688980957
transform -1 0 28888 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1688980957
transform 1 0 27692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1688980957
transform 1 0 29440 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1216_
timestamp 1688980957
transform -1 0 30636 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1688980957
transform -1 0 31464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1218_
timestamp 1688980957
transform -1 0 31464 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1688980957
transform -1 0 31740 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1220_
timestamp 1688980957
transform 1 0 28704 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1688980957
transform 1 0 31648 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1222_
timestamp 1688980957
transform 1 0 22632 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1223_
timestamp 1688980957
transform -1 0 25208 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1688980957
transform 1 0 19780 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1688980957
transform 1 0 20976 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1226_
timestamp 1688980957
transform 1 0 20516 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1227_
timestamp 1688980957
transform -1 0 22816 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1228_
timestamp 1688980957
transform 1 0 24932 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1688980957
transform -1 0 22264 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1688980957
transform -1 0 28704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1231_
timestamp 1688980957
transform -1 0 23368 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1232_
timestamp 1688980957
transform 1 0 21528 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1233_
timestamp 1688980957
transform -1 0 25024 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _1234_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21436 0 -1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1235_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 1 19040
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1236_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18124 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1237_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1238_
timestamp 1688980957
transform 1 0 18676 0 -1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 1688980957
transform -1 0 8556 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1240_
timestamp 1688980957
transform 1 0 16928 0 1 22304
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1241_
timestamp 1688980957
transform 1 0 6624 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1242_
timestamp 1688980957
transform -1 0 20148 0 1 26656
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1243_
timestamp 1688980957
transform -1 0 7452 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 1688980957
transform 1 0 4692 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1245_
timestamp 1688980957
transform -1 0 20608 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1246_
timestamp 1688980957
transform -1 0 20240 0 -1 11424
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1247_
timestamp 1688980957
transform 1 0 12880 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1248_
timestamp 1688980957
transform 1 0 18216 0 1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1249_
timestamp 1688980957
transform -1 0 5796 0 -1 23392
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1250_
timestamp 1688980957
transform -1 0 6164 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1251_
timestamp 1688980957
transform -1 0 5336 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1252_
timestamp 1688980957
transform -1 0 12512 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1253_
timestamp 1688980957
transform 1 0 6072 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1254_
timestamp 1688980957
transform -1 0 4968 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1255_
timestamp 1688980957
transform 1 0 8648 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1256_
timestamp 1688980957
transform 1 0 16284 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1257_
timestamp 1688980957
transform -1 0 14628 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1258_
timestamp 1688980957
transform 1 0 19412 0 -1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1259_
timestamp 1688980957
transform -1 0 5336 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1260_
timestamp 1688980957
transform 1 0 8004 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1261_
timestamp 1688980957
transform 1 0 20884 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 1688980957
transform -1 0 8556 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1263_
timestamp 1688980957
transform -1 0 25392 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1264_
timestamp 1688980957
transform -1 0 5244 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1265_
timestamp 1688980957
transform -1 0 4968 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1266_
timestamp 1688980957
transform 1 0 10580 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1267_
timestamp 1688980957
transform 1 0 13892 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 1688980957
transform -1 0 6440 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1269_
timestamp 1688980957
transform 1 0 13800 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1270_
timestamp 1688980957
transform 1 0 10580 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1271_
timestamp 1688980957
transform 1 0 17204 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1272_
timestamp 1688980957
transform 1 0 17020 0 1 28832
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1273_
timestamp 1688980957
transform -1 0 5704 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1274_
timestamp 1688980957
transform -1 0 6072 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1275_
timestamp 1688980957
transform 1 0 13248 0 -1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1276_
timestamp 1688980957
transform 1 0 15640 0 -1 31008
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1277_
timestamp 1688980957
transform 1 0 11960 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1278_
timestamp 1688980957
transform 1 0 20332 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1279_
timestamp 1688980957
transform 1 0 28060 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1280_
timestamp 1688980957
transform 1 0 3956 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1281_
timestamp 1688980957
transform 1 0 29348 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1282_
timestamp 1688980957
transform 1 0 5428 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1283_
timestamp 1688980957
transform -1 0 5336 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1284_
timestamp 1688980957
transform 1 0 29256 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1285_
timestamp 1688980957
transform 1 0 15732 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1286_
timestamp 1688980957
transform 1 0 18952 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1287_
timestamp 1688980957
transform 1 0 18768 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1288_
timestamp 1688980957
transform 1 0 13800 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1289_
timestamp 1688980957
transform 1 0 14628 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1290_
timestamp 1688980957
transform 1 0 21528 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1291_
timestamp 1688980957
transform 1 0 14628 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1292_
timestamp 1688980957
transform 1 0 15548 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1293_
timestamp 1688980957
transform 1 0 21528 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1294_
timestamp 1688980957
transform -1 0 13800 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1295_
timestamp 1688980957
transform 1 0 8648 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1296_
timestamp 1688980957
transform 1 0 10948 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1297_
timestamp 1688980957
transform 1 0 9752 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1298_
timestamp 1688980957
transform 1 0 8096 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1299_
timestamp 1688980957
transform 1 0 8004 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1300_
timestamp 1688980957
transform 1 0 6072 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1301_
timestamp 1688980957
transform 1 0 7452 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1302_
timestamp 1688980957
transform 1 0 14444 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1303_
timestamp 1688980957
transform 1 0 11224 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1304_
timestamp 1688980957
transform 1 0 7544 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1305_
timestamp 1688980957
transform 1 0 15824 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1306_
timestamp 1688980957
transform 1 0 6992 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1307_
timestamp 1688980957
transform 1 0 16376 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1308_
timestamp 1688980957
transform -1 0 8832 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1309_
timestamp 1688980957
transform 1 0 6072 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1310_
timestamp 1688980957
transform 1 0 17664 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1311_
timestamp 1688980957
transform -1 0 18768 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1312_
timestamp 1688980957
transform 1 0 12604 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1313_
timestamp 1688980957
transform 1 0 17664 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1314_
timestamp 1688980957
transform 1 0 4232 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1315_
timestamp 1688980957
transform 1 0 4968 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1316_
timestamp 1688980957
transform 1 0 4232 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1317_
timestamp 1688980957
transform 1 0 10212 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1318_
timestamp 1688980957
transform 1 0 7360 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1319_
timestamp 1688980957
transform -1 0 11224 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1320_
timestamp 1688980957
transform 1 0 8372 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1321_
timestamp 1688980957
transform 1 0 15824 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1322_
timestamp 1688980957
transform 1 0 10856 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1323_
timestamp 1688980957
transform 1 0 17664 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1324_
timestamp 1688980957
transform 1 0 7268 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1325_
timestamp 1688980957
transform -1 0 9844 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1326_
timestamp 1688980957
transform -1 0 20608 0 -1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1327_
timestamp 1688980957
transform 1 0 8004 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1328_
timestamp 1688980957
transform 1 0 18768 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1329_
timestamp 1688980957
transform -1 0 7084 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1330_
timestamp 1688980957
transform 1 0 4692 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1331_
timestamp 1688980957
transform 1 0 8648 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1332_
timestamp 1688980957
transform 1 0 12512 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1333_
timestamp 1688980957
transform 1 0 6072 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1334_
timestamp 1688980957
transform 1 0 13064 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1335_
timestamp 1688980957
transform 1 0 10028 0 -1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1336_
timestamp 1688980957
transform 1 0 13800 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1337_
timestamp 1688980957
transform 1 0 14720 0 -1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1338_
timestamp 1688980957
transform -1 0 10120 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1339_
timestamp 1688980957
transform -1 0 10488 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1340_
timestamp 1688980957
transform 1 0 11316 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1341_
timestamp 1688980957
transform 1 0 13984 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1342_
timestamp 1688980957
transform -1 0 16376 0 -1 12512
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1343_
timestamp 1688980957
transform -1 0 15088 0 1 12512
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1344_
timestamp 1688980957
transform 1 0 11592 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1345_
timestamp 1688980957
transform 1 0 10580 0 -1 13600
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1346_
timestamp 1688980957
transform 1 0 12328 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1347_
timestamp 1688980957
transform 1 0 12512 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1348_
timestamp 1688980957
transform 1 0 15180 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1349_
timestamp 1688980957
transform 1 0 29072 0 1 15776
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1350_
timestamp 1688980957
transform 1 0 28612 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1351_
timestamp 1688980957
transform 1 0 21344 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1352_
timestamp 1688980957
transform 1 0 21528 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1353_
timestamp 1688980957
transform 1 0 22080 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1354_
timestamp 1688980957
transform 1 0 23460 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1355_
timestamp 1688980957
transform 1 0 26036 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1356_
timestamp 1688980957
transform 1 0 27508 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1357_
timestamp 1688980957
transform 1 0 28244 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1358_
timestamp 1688980957
transform 1 0 28888 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1359_
timestamp 1688980957
transform 1 0 29256 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1360_
timestamp 1688980957
transform 1 0 28888 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1361_
timestamp 1688980957
transform 1 0 26496 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1362_
timestamp 1688980957
transform 1 0 25852 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1363_
timestamp 1688980957
transform -1 0 27876 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1364_
timestamp 1688980957
transform 1 0 23552 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1365_
timestamp 1688980957
transform 1 0 21712 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1366_
timestamp 1688980957
transform 1 0 21712 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1367_
timestamp 1688980957
transform 1 0 26404 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1368_
timestamp 1688980957
transform 1 0 25760 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1369_
timestamp 1688980957
transform -1 0 25392 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1370_
timestamp 1688980957
transform 1 0 22540 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1371_
timestamp 1688980957
transform -1 0 20608 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1372_
timestamp 1688980957
transform 1 0 19320 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1373_
timestamp 1688980957
transform -1 0 28520 0 -1 17952
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1374_
timestamp 1688980957
transform -1 0 20424 0 -1 21216
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1375_
timestamp 1688980957
transform -1 0 30360 0 1 20128
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1376_
timestamp 1688980957
transform -1 0 22080 0 -1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1377_
timestamp 1688980957
transform -1 0 21344 0 -1 23392
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1378_
timestamp 1688980957
transform -1 0 28244 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1379_
timestamp 1688980957
transform -1 0 20700 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1380_
timestamp 1688980957
transform 1 0 19596 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1381_
timestamp 1688980957
transform 1 0 18952 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1382_
timestamp 1688980957
transform -1 0 18860 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1383_
timestamp 1688980957
transform 1 0 16284 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1384_
timestamp 1688980957
transform 1 0 21344 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1385_
timestamp 1688980957
transform 1 0 16376 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1386_
timestamp 1688980957
transform 1 0 16376 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1387_
timestamp 1688980957
transform 1 0 22172 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1388_
timestamp 1688980957
transform 1 0 22540 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1389_
timestamp 1688980957
transform -1 0 31096 0 1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1390_
timestamp 1688980957
transform 1 0 22540 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1391_
timestamp 1688980957
transform 1 0 23736 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1392_
timestamp 1688980957
transform 1 0 25484 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1393_
timestamp 1688980957
transform 1 0 25852 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1394_
timestamp 1688980957
transform 1 0 26036 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1395_
timestamp 1688980957
transform 1 0 26036 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1396_
timestamp 1688980957
transform 1 0 24840 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1397_
timestamp 1688980957
transform -1 0 27876 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1398_
timestamp 1688980957
transform -1 0 26864 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1399_
timestamp 1688980957
transform 1 0 26036 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1400_
timestamp 1688980957
transform 1 0 26680 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1401_
timestamp 1688980957
transform 1 0 28520 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1402_
timestamp 1688980957
transform 1 0 29072 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1403_
timestamp 1688980957
transform 1 0 29532 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1404_
timestamp 1688980957
transform 1 0 29348 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1405_
timestamp 1688980957
transform 1 0 29256 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1406_
timestamp 1688980957
transform 1 0 29072 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1407_
timestamp 1688980957
transform 1 0 28980 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1408_
timestamp 1688980957
transform 1 0 21620 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1409_
timestamp 1688980957
transform 1 0 21436 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1410_
timestamp 1688980957
transform 1 0 19412 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1411_
timestamp 1688980957
transform -1 0 22356 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1412_
timestamp 1688980957
transform -1 0 22724 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1413_
timestamp 1688980957
transform -1 0 23460 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1414_
timestamp 1688980957
transform 1 0 24840 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1415_
timestamp 1688980957
transform -1 0 22908 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1416_
timestamp 1688980957
transform 1 0 26404 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1417_
timestamp 1688980957
transform -1 0 23092 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1418_
timestamp 1688980957
transform -1 0 23184 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1419_
timestamp 1688980957
transform 1 0 23736 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _1420_ Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B1
timestamp 1688980957
transform 1 0 28888 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1688980957
transform -1 0 31832 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1688980957
transform 1 0 29164 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1688980957
transform 1 0 28612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1688980957
transform 1 0 25300 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B
timestamp 1688980957
transform 1 0 24932 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__S
timestamp 1688980957
transform 1 0 25944 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__S
timestamp 1688980957
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__S
timestamp 1688980957
transform 1 0 18860 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__S
timestamp 1688980957
transform 1 0 24656 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__S
timestamp 1688980957
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__S
timestamp 1688980957
transform 1 0 19872 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__S
timestamp 1688980957
transform 1 0 20608 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__S
timestamp 1688980957
transform 1 0 21712 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1
timestamp 1688980957
transform 1 0 25392 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1
timestamp 1688980957
transform -1 0 21712 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A1
timestamp 1688980957
transform 1 0 28888 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A1
timestamp 1688980957
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A1
timestamp 1688980957
transform 1 0 27784 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__C
timestamp 1688980957
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B
timestamp 1688980957
transform 1 0 12236 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__D_N
timestamp 1688980957
transform 1 0 11132 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A
timestamp 1688980957
transform 1 0 15824 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B
timestamp 1688980957
transform 1 0 15364 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__D_N
timestamp 1688980957
transform 1 0 15548 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A_N
timestamp 1688980957
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__B
timestamp 1688980957
transform 1 0 13340 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__C
timestamp 1688980957
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__D
timestamp 1688980957
transform -1 0 14260 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A1
timestamp 1688980957
transform 1 0 15180 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A2
timestamp 1688980957
transform 1 0 16192 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B
timestamp 1688980957
transform -1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1688980957
transform 1 0 15272 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B1
timestamp 1688980957
transform 1 0 12788 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__C_N
timestamp 1688980957
transform -1 0 13248 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A1_N
timestamp 1688980957
transform 1 0 13800 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B1
timestamp 1688980957
transform 1 0 13340 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A1_N
timestamp 1688980957
transform 1 0 12788 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B
timestamp 1688980957
transform -1 0 11040 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__C_N
timestamp 1688980957
transform 1 0 10488 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A1_N
timestamp 1688980957
transform -1 0 10672 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B1
timestamp 1688980957
transform 1 0 10304 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B
timestamp 1688980957
transform 1 0 11500 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__C_N
timestamp 1688980957
transform 1 0 11868 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A1_N
timestamp 1688980957
transform 1 0 10764 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B1
timestamp 1688980957
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B
timestamp 1688980957
transform -1 0 13984 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A1_N
timestamp 1688980957
transform -1 0 16468 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B1
timestamp 1688980957
transform 1 0 15916 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B
timestamp 1688980957
transform 1 0 11868 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__C_N
timestamp 1688980957
transform -1 0 11684 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A1_N
timestamp 1688980957
transform 1 0 13432 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B1
timestamp 1688980957
transform 1 0 13800 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__C_N
timestamp 1688980957
transform 1 0 11868 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A1_N
timestamp 1688980957
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B1
timestamp 1688980957
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__C_N
timestamp 1688980957
transform 1 0 15916 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A1_N
timestamp 1688980957
transform 1 0 13524 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__B1
timestamp 1688980957
transform 1 0 14628 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B
timestamp 1688980957
transform 1 0 11776 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A2
timestamp 1688980957
transform 1 0 7728 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1688980957
transform 1 0 7544 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B2
timestamp 1688980957
transform -1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A2
timestamp 1688980957
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B1
timestamp 1688980957
transform 1 0 12512 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B2
timestamp 1688980957
transform 1 0 13248 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1
timestamp 1688980957
transform 1 0 10028 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B2
timestamp 1688980957
transform 1 0 10488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B1
timestamp 1688980957
transform -1 0 5336 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B2
timestamp 1688980957
transform 1 0 6716 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A2
timestamp 1688980957
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1688980957
transform 1 0 6072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B2
timestamp 1688980957
transform 1 0 7636 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A2
timestamp 1688980957
transform 1 0 17664 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B1
timestamp 1688980957
transform 1 0 18032 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B2
timestamp 1688980957
transform -1 0 19136 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A2
timestamp 1688980957
transform 1 0 8924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B1
timestamp 1688980957
transform 1 0 9476 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B2
timestamp 1688980957
transform -1 0 10028 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A2
timestamp 1688980957
transform -1 0 16744 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B1
timestamp 1688980957
transform -1 0 16376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B2
timestamp 1688980957
transform -1 0 18768 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A2
timestamp 1688980957
transform 1 0 10396 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__B2
timestamp 1688980957
transform 1 0 11040 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B2
timestamp 1688980957
transform -1 0 7268 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A2
timestamp 1688980957
transform 1 0 17112 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B2
timestamp 1688980957
transform -1 0 18676 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1688980957
transform 1 0 12328 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B2
timestamp 1688980957
transform -1 0 13800 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A2
timestamp 1688980957
transform 1 0 16928 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B2
timestamp 1688980957
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B2
timestamp 1688980957
transform 1 0 8556 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__B2
timestamp 1688980957
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A2
timestamp 1688980957
transform 1 0 12512 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B1
timestamp 1688980957
transform 1 0 11132 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B2
timestamp 1688980957
transform 1 0 12144 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A2
timestamp 1688980957
transform 1 0 6624 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B1
timestamp 1688980957
transform -1 0 6348 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B2
timestamp 1688980957
transform 1 0 6992 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A2
timestamp 1688980957
transform 1 0 7360 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B1
timestamp 1688980957
transform 1 0 6992 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1
timestamp 1688980957
transform 1 0 8188 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B2
timestamp 1688980957
transform -1 0 8004 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A2
timestamp 1688980957
transform 1 0 17756 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B1
timestamp 1688980957
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B2
timestamp 1688980957
transform -1 0 17848 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A2
timestamp 1688980957
transform 1 0 12880 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B1
timestamp 1688980957
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B2
timestamp 1688980957
transform 1 0 12512 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A2
timestamp 1688980957
transform 1 0 16560 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B1
timestamp 1688980957
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A2
timestamp 1688980957
transform 1 0 17480 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B1
timestamp 1688980957
transform 1 0 18032 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__B2
timestamp 1688980957
transform -1 0 19596 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A2
timestamp 1688980957
transform 1 0 9660 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A2
timestamp 1688980957
transform 1 0 18032 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A2
timestamp 1688980957
transform 1 0 9108 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A2
timestamp 1688980957
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A2
timestamp 1688980957
transform 1 0 10212 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A2
timestamp 1688980957
transform 1 0 12144 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A0
timestamp 1688980957
transform 1 0 7728 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A0
timestamp 1688980957
transform 1 0 10304 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A0
timestamp 1688980957
transform 1 0 9200 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A0
timestamp 1688980957
transform -1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A0
timestamp 1688980957
transform 1 0 11592 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A0
timestamp 1688980957
transform 1 0 13984 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__S0
timestamp 1688980957
transform 1 0 29624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__S1
timestamp 1688980957
transform -1 0 30544 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A0
timestamp 1688980957
transform 1 0 12696 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A1
timestamp 1688980957
transform -1 0 13064 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__S0
timestamp 1688980957
transform 1 0 13432 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__S1
timestamp 1688980957
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A1
timestamp 1688980957
transform 1 0 13432 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__S0
timestamp 1688980957
transform 1 0 13800 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__S1
timestamp 1688980957
transform 1 0 13984 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A1
timestamp 1688980957
transform -1 0 30728 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__S0
timestamp 1688980957
transform -1 0 31556 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__S1
timestamp 1688980957
transform 1 0 30912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1688980957
transform -1 0 10672 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__S0
timestamp 1688980957
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__S1
timestamp 1688980957
transform 1 0 12604 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1688980957
transform -1 0 13800 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__S0
timestamp 1688980957
transform 1 0 15456 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__S1
timestamp 1688980957
transform 1 0 14260 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A0
timestamp 1688980957
transform -1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__S0
timestamp 1688980957
transform -1 0 16744 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__S1
timestamp 1688980957
transform 1 0 15456 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__S0
timestamp 1688980957
transform -1 0 18216 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__S1
timestamp 1688980957
transform -1 0 18584 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B
timestamp 1688980957
transform -1 0 20700 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B
timestamp 1688980957
transform 1 0 12236 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1688980957
transform 1 0 28980 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__S
timestamp 1688980957
transform 1 0 29164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__S
timestamp 1688980957
transform 1 0 5612 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A1
timestamp 1688980957
transform -1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__S
timestamp 1688980957
transform 1 0 6256 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1688980957
transform -1 0 28980 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__S
timestamp 1688980957
transform -1 0 28888 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__S
timestamp 1688980957
transform 1 0 6440 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1688980957
transform 1 0 28244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__S
timestamp 1688980957
transform 1 0 28428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1688980957
transform -1 0 19688 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__S
timestamp 1688980957
transform 1 0 21528 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A1
timestamp 1688980957
transform -1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__S
timestamp 1688980957
transform 1 0 12328 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__S
timestamp 1688980957
transform 1 0 15456 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__S
timestamp 1688980957
transform 1 0 13156 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__S
timestamp 1688980957
transform 1 0 6256 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__S
timestamp 1688980957
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__S
timestamp 1688980957
transform 1 0 15548 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__S
timestamp 1688980957
transform 1 0 16560 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__S
timestamp 1688980957
transform 1 0 10856 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__S
timestamp 1688980957
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__S
timestamp 1688980957
transform 1 0 6900 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__S
timestamp 1688980957
transform 1 0 12144 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__S
timestamp 1688980957
transform 1 0 10764 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__S
timestamp 1688980957
transform 1 0 4784 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__S
timestamp 1688980957
transform 1 0 6256 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__S
timestamp 1688980957
transform 1 0 23736 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__S
timestamp 1688980957
transform 1 0 7452 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__S
timestamp 1688980957
transform 1 0 20792 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__S
timestamp 1688980957
transform 1 0 9752 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__S
timestamp 1688980957
transform 1 0 5428 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__S
timestamp 1688980957
transform 1 0 19504 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__S
timestamp 1688980957
transform -1 0 14168 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__S
timestamp 1688980957
transform -1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__S
timestamp 1688980957
transform 1 0 9200 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__S
timestamp 1688980957
transform -1 0 3404 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__S
timestamp 1688980957
transform 1 0 6992 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A2
timestamp 1688980957
transform 1 0 15824 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__S
timestamp 1688980957
transform -1 0 13064 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__S
timestamp 1688980957
transform 1 0 5612 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__S
timestamp 1688980957
transform -1 0 6532 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__S
timestamp 1688980957
transform 1 0 6624 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__S
timestamp 1688980957
transform 1 0 16652 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__S
timestamp 1688980957
transform -1 0 15640 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__S
timestamp 1688980957
transform 1 0 17664 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__S
timestamp 1688980957
transform 1 0 18492 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__S
timestamp 1688980957
transform 1 0 6716 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__S
timestamp 1688980957
transform -1 0 10212 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__S
timestamp 1688980957
transform -1 0 18952 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__S
timestamp 1688980957
transform 1 0 9292 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__S
timestamp 1688980957
transform 1 0 18584 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__S
timestamp 1688980957
transform 1 0 9016 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__S
timestamp 1688980957
transform 1 0 19780 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__S
timestamp 1688980957
transform 1 0 15456 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A
timestamp 1688980957
transform 1 0 14444 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1688980957
transform -1 0 10488 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A
timestamp 1688980957
transform 1 0 18768 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__A
timestamp 1688980957
transform 1 0 4968 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_clk_A
timestamp 1688980957
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_clk_A
timestamp 1688980957
transform 1 0 10304 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_clk_A
timestamp 1688980957
transform 1 0 14812 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_clk_A
timestamp 1688980957
transform 1 0 14444 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_clk_A
timestamp 1688980957
transform 1 0 11316 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_clk_A
timestamp 1688980957
transform 1 0 10948 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_clk_A
timestamp 1688980957
transform 1 0 12788 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_clk_A
timestamp 1688980957
transform 1 0 12236 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_clk_A
timestamp 1688980957
transform 1 0 20608 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_clk_A
timestamp 1688980957
transform 1 0 20608 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_clk_A
timestamp 1688980957
transform 1 0 24196 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_clk_A
timestamp 1688980957
transform 1 0 27324 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_clk_A
timestamp 1688980957
transform 1 0 21528 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_clk_A
timestamp 1688980957
transform 1 0 21344 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_clk_A
timestamp 1688980957
transform 1 0 26220 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_clk_A
timestamp 1688980957
transform -1 0 28336 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout89_A
timestamp 1688980957
transform 1 0 9016 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout90_A
timestamp 1688980957
transform 1 0 6624 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout91_A
timestamp 1688980957
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout92_A
timestamp 1688980957
transform -1 0 17296 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout100_A
timestamp 1688980957
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout101_A
timestamp 1688980957
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout102_A
timestamp 1688980957
transform 1 0 24380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1688980957
transform 1 0 30636 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1688980957
transform -1 0 31556 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1688980957
transform 1 0 30176 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1688980957
transform -1 0 31924 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp 1688980957
transform 1 0 18216 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 1688980957
transform 1 0 18032 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 1688980957
transform 1 0 16928 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout114_A
timestamp 1688980957
transform -1 0 30084 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold91_A
timestamp 1688980957
transform 1 0 13984 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold161_A
timestamp 1688980957
transform 1 0 12880 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold163_A
timestamp 1688980957
transform -1 0 18032 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold167_A
timestamp 1688980957
transform 1 0 16744 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold172_A
timestamp 1688980957
transform 1 0 24748 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold174_A
timestamp 1688980957
transform 1 0 21068 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold208_A
timestamp 1688980957
transform 1 0 14996 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold228_A
timestamp 1688980957
transform 1 0 12880 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold303_A
timestamp 1688980957
transform 1 0 19136 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1688980957
transform 1 0 28888 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9936 0 1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1688980957
transform -1 0 9660 0 1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1688980957
transform -1 0 14168 0 -1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1688980957
transform 1 0 13432 0 -1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1688980957
transform 1 0 8740 0 -1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1688980957
transform -1 0 10764 0 -1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1688980957
transform 1 0 14260 0 1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1688980957
transform -1 0 14444 0 -1 24480
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1688980957
transform -1 0 22264 0 1 10336
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1688980957
transform 1 0 20884 0 1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1688980957
transform -1 0 27048 0 1 11424
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1688980957
transform -1 0 27140 0 -1 12512
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1688980957
transform 1 0 21712 0 -1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1688980957
transform 1 0 21804 0 1 23392
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1688980957
transform -1 0 26864 0 -1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1688980957
transform 1 0 26036 0 1 22304
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout89 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout90
timestamp 1688980957
transform -1 0 6624 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout91 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10488 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout92
timestamp 1688980957
transform 1 0 17020 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout93
timestamp 1688980957
transform 1 0 17112 0 1 21216
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout96
timestamp 1688980957
transform -1 0 24932 0 1 13600
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout97
timestamp 1688980957
transform -1 0 26588 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout98 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29256 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_8  fanout99
timestamp 1688980957
transform -1 0 14720 0 -1 14688
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout100 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16468 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout101
timestamp 1688980957
transform 1 0 16836 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout102
timestamp 1688980957
transform -1 0 23828 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout103
timestamp 1688980957
transform 1 0 31188 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout104
timestamp 1688980957
transform -1 0 31096 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout105
timestamp 1688980957
transform -1 0 30728 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout106
timestamp 1688980957
transform -1 0 29992 0 1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout107
timestamp 1688980957
transform -1 0 11592 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout108
timestamp 1688980957
transform 1 0 17664 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout109
timestamp 1688980957
transform -1 0 17848 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout110
timestamp 1688980957
transform -1 0 16744 0 1 27744
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout111
timestamp 1688980957
transform -1 0 31556 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout112
timestamp 1688980957
transform -1 0 25208 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout113
timestamp 1688980957
transform 1 0 31188 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout114
timestamp 1688980957
transform -1 0 31740 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_22 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_29 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5428 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_33 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50
timestamp 1688980957
transform 1 0 7360 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9752 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 10580 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_93 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1688980957
transform 1 0 13156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1688980957
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_121
timestamp 1688980957
transform 1 0 13892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_141
timestamp 1688980957
transform 1 0 15732 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1688980957
transform 1 0 16100 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_148 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16376 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_169
timestamp 1688980957
transform 1 0 18308 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_174
timestamp 1688980957
transform 1 0 18768 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_178
timestamp 1688980957
transform 1 0 19136 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_197
timestamp 1688980957
transform 1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_201
timestamp 1688980957
transform 1 0 21252 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_205 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21620 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_217
timestamp 1688980957
transform 1 0 22724 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 23276 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_241
timestamp 1688980957
transform 1 0 24932 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 25668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_272
timestamp 1688980957
transform 1 0 27784 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_281
timestamp 1688980957
transform 1 0 28612 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_289
timestamp 1688980957
transform 1 0 29348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_309
timestamp 1688980957
transform 1 0 31188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_19
timestamp 1688980957
transform 1 0 4508 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_36
timestamp 1688980957
transform 1 0 6072 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_40
timestamp 1688980957
transform 1 0 6440 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 1688980957
transform 1 0 7544 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_81
timestamp 1688980957
transform 1 0 10212 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_99
timestamp 1688980957
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 12972 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_113
timestamp 1688980957
transform 1 0 13156 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_117
timestamp 1688980957
transform 1 0 13524 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_141
timestamp 1688980957
transform 1 0 15732 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_145
timestamp 1688980957
transform 1 0 16100 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_148
timestamp 1688980957
transform 1 0 16376 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_172
timestamp 1688980957
transform 1 0 18584 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_194
timestamp 1688980957
transform 1 0 20608 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_218
timestamp 1688980957
transform 1 0 22816 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 23276 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_225
timestamp 1688980957
transform 1 0 23460 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_230
timestamp 1688980957
transform 1 0 23920 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_236
timestamp 1688980957
transform 1 0 24472 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_253
timestamp 1688980957
transform 1 0 26036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_265
timestamp 1688980957
transform 1 0 27140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 1688980957
transform 1 0 28244 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_281
timestamp 1688980957
transform 1 0 28612 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_316
timestamp 1688980957
transform 1 0 31832 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_9
timestamp 1688980957
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_21
timestamp 1688980957
transform 1 0 4692 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 5244 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_49
timestamp 1688980957
transform 1 0 7268 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_61
timestamp 1688980957
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_73
timestamp 1688980957
transform 1 0 9476 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_81
timestamp 1688980957
transform 1 0 10212 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_97
timestamp 1688980957
transform 1 0 11684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 1688980957
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_225
timestamp 1688980957
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1688980957
transform 1 0 25668 0 1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 26036 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_265
timestamp 1688980957
transform 1 0 27140 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_273
timestamp 1688980957
transform 1 0 27876 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_298
timestamp 1688980957
transform 1 0 30176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_302
timestamp 1688980957
transform 1 0 30544 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_309
timestamp 1688980957
transform 1 0 31188 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_15
timestamp 1688980957
transform 1 0 4140 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_19
timestamp 1688980957
transform 1 0 4508 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_52
timestamp 1688980957
transform 1 0 7544 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1688980957
transform 1 0 9108 0 -1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_78
timestamp 1688980957
transform 1 0 9936 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_90
timestamp 1688980957
transform 1 0 11040 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_104
timestamp 1688980957
transform 1 0 12328 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_108
timestamp 1688980957
transform 1 0 12696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_113
timestamp 1688980957
transform 1 0 13156 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_119
timestamp 1688980957
transform 1 0 13708 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_163
timestamp 1688980957
transform 1 0 17756 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_203
timestamp 1688980957
transform 1 0 21436 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_228
timestamp 1688980957
transform 1 0 23736 0 -1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_247
timestamp 1688980957
transform 1 0 25484 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_259
timestamp 1688980957
transform 1 0 26588 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_271
timestamp 1688980957
transform 1 0 27692 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 28428 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_290
timestamp 1688980957
transform 1 0 29440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_294
timestamp 1688980957
transform 1 0 29808 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_19
timestamp 1688980957
transform 1 0 4508 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 5244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_29
timestamp 1688980957
transform 1 0 5428 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_43
timestamp 1688980957
transform 1 0 6716 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_55
timestamp 1688980957
transform 1 0 7820 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_63
timestamp 1688980957
transform 1 0 8556 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_97
timestamp 1688980957
transform 1 0 11684 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_103
timestamp 1688980957
transform 1 0 12236 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_135
timestamp 1688980957
transform 1 0 15180 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_158
timestamp 1688980957
transform 1 0 17296 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_180
timestamp 1688980957
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_204
timestamp 1688980957
transform 1 0 21528 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_246
timestamp 1688980957
transform 1 0 25392 0 1 4896
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 26036 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 27140 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_277
timestamp 1688980957
transform 1 0 28244 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_281
timestamp 1688980957
transform 1 0 28612 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_289
timestamp 1688980957
transform 1 0 29348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_298
timestamp 1688980957
transform 1 0 30176 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_306
timestamp 1688980957
transform 1 0 30912 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_309
timestamp 1688980957
transform 1 0 31188 0 1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_27
timestamp 1688980957
transform 1 0 5244 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_60
timestamp 1688980957
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_68
timestamp 1688980957
transform 1 0 9016 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 10212 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 11316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_105
timestamp 1688980957
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_108
timestamp 1688980957
transform 1 0 12696 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_113
timestamp 1688980957
transform 1 0 13156 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_159
timestamp 1688980957
transform 1 0 17388 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_164
timestamp 1688980957
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_169
timestamp 1688980957
transform 1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_205
timestamp 1688980957
transform 1 0 21620 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1688980957
transform 1 0 23184 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_250
timestamp 1688980957
transform 1 0 25760 0 -1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_254
timestamp 1688980957
transform 1 0 26128 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_266
timestamp 1688980957
transform 1 0 27232 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_270
timestamp 1688980957
transform 1 0 27600 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_274
timestamp 1688980957
transform 1 0 27968 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_285
timestamp 1688980957
transform 1 0 28980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_289
timestamp 1688980957
transform 1 0 29348 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 29716 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 30820 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_6
timestamp 1688980957
transform 1 0 3312 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_18
timestamp 1688980957
transform 1 0 4416 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1688980957
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_41
timestamp 1688980957
transform 1 0 6532 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_50
timestamp 1688980957
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_60
timestamp 1688980957
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_68
timestamp 1688980957
transform 1 0 9016 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_78
timestamp 1688980957
transform 1 0 9936 0 1 5984
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_97
timestamp 1688980957
transform 1 0 11684 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_105
timestamp 1688980957
transform 1 0 12420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_118
timestamp 1688980957
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_136
timestamp 1688980957
transform 1 0 15272 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_166
timestamp 1688980957
transform 1 0 18032 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_172
timestamp 1688980957
transform 1 0 18584 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_200
timestamp 1688980957
transform 1 0 21160 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_208
timestamp 1688980957
transform 1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_247
timestamp 1688980957
transform 1 0 25484 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 25852 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_253
timestamp 1688980957
transform 1 0 26036 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_259
timestamp 1688980957
transform 1 0 26588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_303
timestamp 1688980957
transform 1 0 30636 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 31004 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_309
timestamp 1688980957
transform 1 0 31188 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_313
timestamp 1688980957
transform 1 0 31556 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 5244 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_39
timestamp 1688980957
transform 1 0 6348 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_52
timestamp 1688980957
transform 1 0 7544 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1688980957
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_61
timestamp 1688980957
transform 1 0 8372 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_73
timestamp 1688980957
transform 1 0 9476 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_85
timestamp 1688980957
transform 1 0 10580 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_97
timestamp 1688980957
transform 1 0 11684 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_105
timestamp 1688980957
transform 1 0 12420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_108
timestamp 1688980957
transform 1 0 12696 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_120
timestamp 1688980957
transform 1 0 13800 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_124
timestamp 1688980957
transform 1 0 14168 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_140
timestamp 1688980957
transform 1 0 15640 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_202
timestamp 1688980957
transform 1 0 21344 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_214
timestamp 1688980957
transform 1 0 22448 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_219
timestamp 1688980957
transform 1 0 22908 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 23276 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_239
timestamp 1688980957
transform 1 0 24748 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_243
timestamp 1688980957
transform 1 0 25116 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_251
timestamp 1688980957
transform 1 0 25852 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_275
timestamp 1688980957
transform 1 0 28060 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_305
timestamp 1688980957
transform 1 0 30820 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_309
timestamp 1688980957
transform 1 0 31188 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_313
timestamp 1688980957
transform 1 0 31556 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 3036 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 4140 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 5244 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_41
timestamp 1688980957
transform 1 0 6532 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_49
timestamp 1688980957
transform 1 0 7268 0 1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_54
timestamp 1688980957
transform 1 0 7728 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_66
timestamp 1688980957
transform 1 0 8832 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 1688980957
transform 1 0 9936 0 1 7072
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_109
timestamp 1688980957
transform 1 0 12788 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_113
timestamp 1688980957
transform 1 0 13156 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_116
timestamp 1688980957
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_168
timestamp 1688980957
transform 1 0 18216 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_172
timestamp 1688980957
transform 1 0 18584 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_184
timestamp 1688980957
transform 1 0 19688 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_192
timestamp 1688980957
transform 1 0 20424 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 1688980957
transform 1 0 20884 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_226
timestamp 1688980957
transform 1 0 23552 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 1688980957
transform 1 0 25668 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_306
timestamp 1688980957
transform 1 0 30912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_309
timestamp 1688980957
transform 1 0 31188 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_6
timestamp 1688980957
transform 1 0 3312 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_14
timestamp 1688980957
transform 1 0 4048 0 -1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 6348 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 7452 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 7820 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 10212 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 11316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 12420 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 12972 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_134
timestamp 1688980957
transform 1 0 15088 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_147
timestamp 1688980957
transform 1 0 16284 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_177
timestamp 1688980957
transform 1 0 19044 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_199
timestamp 1688980957
transform 1 0 21068 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_220
timestamp 1688980957
transform 1 0 23000 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 1688980957
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_238
timestamp 1688980957
transform 1 0 24656 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1688980957
transform 1 0 28336 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_287
timestamp 1688980957
transform 1 0 29164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_308
timestamp 1688980957
transform 1 0 31096 0 -1 8160
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 3036 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 4140 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 5244 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_46
timestamp 1688980957
transform 1 0 6992 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_58
timestamp 1688980957
transform 1 0 8096 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_70
timestamp 1688980957
transform 1 0 9200 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_97
timestamp 1688980957
transform 1 0 11684 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_105
timestamp 1688980957
transform 1 0 12420 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_109
timestamp 1688980957
transform 1 0 12788 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_131
timestamp 1688980957
transform 1 0 14812 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_184
timestamp 1688980957
transform 1 0 19688 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_188
timestamp 1688980957
transform 1 0 20056 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_197
timestamp 1688980957
transform 1 0 20884 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_209
timestamp 1688980957
transform 1 0 21988 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_229
timestamp 1688980957
transform 1 0 23828 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_233
timestamp 1688980957
transform 1 0 24196 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_237
timestamp 1688980957
transform 1 0 24564 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_246
timestamp 1688980957
transform 1 0 25392 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_279
timestamp 1688980957
transform 1 0 28428 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_312
timestamp 1688980957
transform 1 0 31464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_316
timestamp 1688980957
transform 1 0 31832 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_27
timestamp 1688980957
transform 1 0 5244 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_35
timestamp 1688980957
transform 1 0 5980 0 -1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_40
timestamp 1688980957
transform 1 0 6440 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_52
timestamp 1688980957
transform 1 0 7544 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_81
timestamp 1688980957
transform 1 0 10212 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_107
timestamp 1688980957
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 12972 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_113
timestamp 1688980957
transform 1 0 13156 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_118
timestamp 1688980957
transform 1 0 13616 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_172
timestamp 1688980957
transform 1 0 18584 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_201
timestamp 1688980957
transform 1 0 21252 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 23276 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_244
timestamp 1688980957
transform 1 0 25208 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_255
timestamp 1688980957
transform 1 0 26220 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_260
timestamp 1688980957
transform 1 0 26680 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_264
timestamp 1688980957
transform 1 0 27048 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_277
timestamp 1688980957
transform 1 0 28244 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_289
timestamp 1688980957
transform 1 0 29348 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 3036 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 4140 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 5244 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 6532 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_53
timestamp 1688980957
transform 1 0 7636 0 1 9248
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_67
timestamp 1688980957
transform 1 0 8924 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_79
timestamp 1688980957
transform 1 0 10028 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 10396 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 12788 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_121
timestamp 1688980957
transform 1 0 13892 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_131
timestamp 1688980957
transform 1 0 14812 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_159
timestamp 1688980957
transform 1 0 17388 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_173
timestamp 1688980957
transform 1 0 18676 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_177
timestamp 1688980957
transform 1 0 19044 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 20884 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_233
timestamp 1688980957
transform 1 0 24196 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_258
timestamp 1688980957
transform 1 0 26496 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_288
timestamp 1688980957
transform 1 0 29256 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_6
timestamp 1688980957
transform 1 0 3312 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_14
timestamp 1688980957
transform 1 0 4048 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_37
timestamp 1688980957
transform 1 0 6164 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1688980957
transform 1 0 6532 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1688980957
transform 1 0 7636 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 8004 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_69
timestamp 1688980957
transform 1 0 9108 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_75
timestamp 1688980957
transform 1 0 9660 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_82
timestamp 1688980957
transform 1 0 10304 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_86
timestamp 1688980957
transform 1 0 10672 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_98
timestamp 1688980957
transform 1 0 11776 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1688980957
transform 1 0 13156 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_121
timestamp 1688980957
transform 1 0 13892 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_125
timestamp 1688980957
transform 1 0 14260 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_152
timestamp 1688980957
transform 1 0 16744 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_162
timestamp 1688980957
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 18032 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_172
timestamp 1688980957
transform 1 0 18584 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_176
timestamp 1688980957
transform 1 0 18952 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_184
timestamp 1688980957
transform 1 0 19688 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_188
timestamp 1688980957
transform 1 0 20056 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_192
timestamp 1688980957
transform 1 0 20424 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 23184 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_238
timestamp 1688980957
transform 1 0 24656 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_246
timestamp 1688980957
transform 1 0 25392 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_252
timestamp 1688980957
transform 1 0 25944 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_259
timestamp 1688980957
transform 1 0 26588 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_272
timestamp 1688980957
transform 1 0 27784 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_281
timestamp 1688980957
transform 1 0 28612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_315
timestamp 1688980957
transform 1 0 31740 0 -1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 3036 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_15
timestamp 1688980957
transform 1 0 4140 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_19
timestamp 1688980957
transform 1 0 4508 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_46
timestamp 1688980957
transform 1 0 6992 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_54
timestamp 1688980957
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_109
timestamp 1688980957
transform 1 0 12788 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_132
timestamp 1688980957
transform 1 0 14904 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 15548 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_141
timestamp 1688980957
transform 1 0 15732 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_178
timestamp 1688980957
transform 1 0 19136 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_190
timestamp 1688980957
transform 1 0 20240 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_197
timestamp 1688980957
transform 1 0 20884 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_215
timestamp 1688980957
transform 1 0 22540 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_219
timestamp 1688980957
transform 1 0 22908 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_234
timestamp 1688980957
transform 1 0 24288 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_242
timestamp 1688980957
transform 1 0 25024 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_281
timestamp 1688980957
transform 1 0 28612 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_285
timestamp 1688980957
transform 1 0 28980 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 31004 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_315
timestamp 1688980957
transform 1 0 31740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_19
timestamp 1688980957
transform 1 0 4508 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_23
timestamp 1688980957
transform 1 0 4876 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_44
timestamp 1688980957
transform 1 0 6808 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_50
timestamp 1688980957
transform 1 0 7360 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_110
timestamp 1688980957
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1688980957
transform 1 0 13156 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_127
timestamp 1688980957
transform 1 0 14444 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_131
timestamp 1688980957
transform 1 0 14812 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_149
timestamp 1688980957
transform 1 0 16468 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_160
timestamp 1688980957
transform 1 0 17480 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 18124 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_190
timestamp 1688980957
transform 1 0 20240 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_198
timestamp 1688980957
transform 1 0 20976 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_213
timestamp 1688980957
transform 1 0 22356 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_221
timestamp 1688980957
transform 1 0 23092 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 23460 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_237
timestamp 1688980957
transform 1 0 24564 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1688980957
transform 1 0 28336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_291
timestamp 1688980957
transform 1 0 29532 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_295
timestamp 1688980957
transform 1 0 29900 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_300
timestamp 1688980957
transform 1 0 30360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_308
timestamp 1688980957
transform 1 0 31096 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_315
timestamp 1688980957
transform 1 0 31740 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 3036 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_15
timestamp 1688980957
transform 1 0 4140 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_63
timestamp 1688980957
transform 1 0 8556 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_77
timestamp 1688980957
transform 1 0 9844 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_81
timestamp 1688980957
transform 1 0 10212 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_119
timestamp 1688980957
transform 1 0 13708 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_125
timestamp 1688980957
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_129
timestamp 1688980957
transform 1 0 14628 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_133
timestamp 1688980957
transform 1 0 14996 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 15548 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_149
timestamp 1688980957
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_153
timestamp 1688980957
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_183
timestamp 1688980957
transform 1 0 19596 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_192
timestamp 1688980957
transform 1 0 20424 0 1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_208
timestamp 1688980957
transform 1 0 21896 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_220
timestamp 1688980957
transform 1 0 23000 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_232
timestamp 1688980957
transform 1 0 24104 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_239
timestamp 1688980957
transform 1 0 24748 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_289
timestamp 1688980957
transform 1 0 29348 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_306
timestamp 1688980957
transform 1 0 30912 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1688980957
transform 1 0 3036 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_85
timestamp 1688980957
transform 1 0 10580 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_89
timestamp 1688980957
transform 1 0 10948 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_93
timestamp 1688980957
transform 1 0 11316 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_101
timestamp 1688980957
transform 1 0 12052 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_104
timestamp 1688980957
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_108
timestamp 1688980957
transform 1 0 12696 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_124
timestamp 1688980957
transform 1 0 14168 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_148
timestamp 1688980957
transform 1 0 16376 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_169
timestamp 1688980957
transform 1 0 18308 0 -1 12512
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_191
timestamp 1688980957
transform 1 0 20332 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_203
timestamp 1688980957
transform 1 0 21436 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_208
timestamp 1688980957
transform 1 0 21896 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_221
timestamp 1688980957
transform 1 0 23092 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_233
timestamp 1688980957
transform 1 0 24196 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_241
timestamp 1688980957
transform 1 0 24932 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_265
timestamp 1688980957
transform 1 0 27140 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_269
timestamp 1688980957
transform 1 0 27508 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 27876 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 28428 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_281
timestamp 1688980957
transform 1 0 28612 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_299
timestamp 1688980957
transform 1 0 30268 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 3036 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 4140 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 5244 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1688980957
transform 1 0 5428 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_39
timestamp 1688980957
transform 1 0 6348 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_43
timestamp 1688980957
transform 1 0 6716 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_48
timestamp 1688980957
transform 1 0 7176 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_52
timestamp 1688980957
transform 1 0 7544 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_66
timestamp 1688980957
transform 1 0 8832 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_78
timestamp 1688980957
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1688980957
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1688980957
transform 1 0 10580 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_89
timestamp 1688980957
transform 1 0 10948 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_97
timestamp 1688980957
transform 1 0 11684 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_107
timestamp 1688980957
transform 1 0 12604 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_134
timestamp 1688980957
transform 1 0 15088 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 15456 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1688980957
transform 1 0 15732 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_145
timestamp 1688980957
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_149
timestamp 1688980957
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_160
timestamp 1688980957
transform 1 0 17480 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_164
timestamp 1688980957
transform 1 0 17848 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 20148 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 20700 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_206
timestamp 1688980957
transform 1 0 21712 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_235
timestamp 1688980957
transform 1 0 24380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_247
timestamp 1688980957
transform 1 0 25484 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_306
timestamp 1688980957
transform 1 0 30912 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_19
timestamp 1688980957
transform 1 0 4508 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_31
timestamp 1688980957
transform 1 0 5612 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_43
timestamp 1688980957
transform 1 0 6716 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_51
timestamp 1688980957
transform 1 0 7452 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 7820 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_57
timestamp 1688980957
transform 1 0 8004 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_80
timestamp 1688980957
transform 1 0 10120 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_84
timestamp 1688980957
transform 1 0 10488 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 12972 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_113
timestamp 1688980957
transform 1 0 13156 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_139
timestamp 1688980957
transform 1 0 15548 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_149
timestamp 1688980957
transform 1 0 16468 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_165
timestamp 1688980957
transform 1 0 17940 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1688980957
transform 1 0 18308 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_181
timestamp 1688980957
transform 1 0 19412 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_249
timestamp 1688980957
transform 1 0 25668 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_269
timestamp 1688980957
transform 1 0 27508 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_281
timestamp 1688980957
transform 1 0 28612 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_19
timestamp 1688980957
transform 1 0 4508 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 5244 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_29
timestamp 1688980957
transform 1 0 5428 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_33
timestamp 1688980957
transform 1 0 5796 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_37
timestamp 1688980957
transform 1 0 6164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_40
timestamp 1688980957
transform 1 0 6440 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_63
timestamp 1688980957
transform 1 0 8556 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_78
timestamp 1688980957
transform 1 0 9936 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_93
timestamp 1688980957
transform 1 0 11316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_161
timestamp 1688980957
transform 1 0 17572 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_190
timestamp 1688980957
transform 1 0 20240 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_213
timestamp 1688980957
transform 1 0 22356 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_227
timestamp 1688980957
transform 1 0 23644 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_241
timestamp 1688980957
transform 1 0 24932 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_281
timestamp 1688980957
transform 1 0 28612 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_3
timestamp 1688980957
transform 1 0 3036 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_7
timestamp 1688980957
transform 1 0 3404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_31
timestamp 1688980957
transform 1 0 5612 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_35
timestamp 1688980957
transform 1 0 5980 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_45
timestamp 1688980957
transform 1 0 6900 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_51
timestamp 1688980957
transform 1 0 7452 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 7820 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_60
timestamp 1688980957
transform 1 0 8280 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_79
timestamp 1688980957
transform 1 0 10028 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_83
timestamp 1688980957
transform 1 0 10396 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1688980957
transform 1 0 12880 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_151
timestamp 1688980957
transform 1 0 16652 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_169
timestamp 1688980957
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_183
timestamp 1688980957
transform 1 0 19596 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_194
timestamp 1688980957
transform 1 0 20608 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1688980957
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_235
timestamp 1688980957
transform 1 0 24380 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_243
timestamp 1688980957
transform 1 0 25116 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 28428 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_286
timestamp 1688980957
transform 1 0 29072 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_296
timestamp 1688980957
transform 1 0 29992 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_300
timestamp 1688980957
transform 1 0 30360 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_312
timestamp 1688980957
transform 1 0 31464 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_3
timestamp 1688980957
transform 1 0 3036 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_9
timestamp 1688980957
transform 1 0 3588 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 5244 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_66
timestamp 1688980957
transform 1 0 8832 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_70
timestamp 1688980957
transform 1 0 9200 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_73
timestamp 1688980957
transform 1 0 9476 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_81
timestamp 1688980957
transform 1 0 10212 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_85
timestamp 1688980957
transform 1 0 10580 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_108
timestamp 1688980957
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_135
timestamp 1688980957
transform 1 0 15180 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_175
timestamp 1688980957
transform 1 0 18860 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_197
timestamp 1688980957
transform 1 0 20884 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_209
timestamp 1688980957
transform 1 0 21988 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_236
timestamp 1688980957
transform 1 0 24472 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_240
timestamp 1688980957
transform 1 0 24840 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_248
timestamp 1688980957
transform 1 0 25576 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_289
timestamp 1688980957
transform 1 0 29348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_304
timestamp 1688980957
transform 1 0 30728 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_312
timestamp 1688980957
transform 1 0 31464 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_316
timestamp 1688980957
transform 1 0 31832 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_3
timestamp 1688980957
transform 1 0 3036 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 7820 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1688980957
transform 1 0 8004 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_61
timestamp 1688980957
transform 1 0 8372 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_70
timestamp 1688980957
transform 1 0 9200 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_82
timestamp 1688980957
transform 1 0 10304 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_102
timestamp 1688980957
transform 1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 12972 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_116
timestamp 1688980957
transform 1 0 13432 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_161
timestamp 1688980957
transform 1 0 17572 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_165
timestamp 1688980957
transform 1 0 17940 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_169
timestamp 1688980957
transform 1 0 18308 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_177
timestamp 1688980957
transform 1 0 19044 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_196
timestamp 1688980957
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_203
timestamp 1688980957
transform 1 0 21436 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_239
timestamp 1688980957
transform 1 0 24748 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_274
timestamp 1688980957
transform 1 0 27968 0 -1 15776
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 28612 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_293
timestamp 1688980957
transform 1 0 29716 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_300
timestamp 1688980957
transform 1 0 30360 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_19
timestamp 1688980957
transform 1 0 4508 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 1688980957
transform 1 0 5428 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_45
timestamp 1688980957
transform 1 0 6900 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_50
timestamp 1688980957
transform 1 0 7360 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_67
timestamp 1688980957
transform 1 0 8924 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_71
timestamp 1688980957
transform 1 0 9292 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 10396 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_85
timestamp 1688980957
transform 1 0 10580 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_101
timestamp 1688980957
transform 1 0 12052 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_110
timestamp 1688980957
transform 1 0 12880 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_114
timestamp 1688980957
transform 1 0 13248 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_130
timestamp 1688980957
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_165
timestamp 1688980957
transform 1 0 17940 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_188
timestamp 1688980957
transform 1 0 20056 0 1 15776
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 20884 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_209
timestamp 1688980957
transform 1 0 21988 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_222
timestamp 1688980957
transform 1 0 23184 0 1 15776
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_240
timestamp 1688980957
transform 1 0 24840 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_253
timestamp 1688980957
transform 1 0 26036 0 1 15776
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_264
timestamp 1688980957
transform 1 0 27048 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_276
timestamp 1688980957
transform 1 0 28152 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_284
timestamp 1688980957
transform 1 0 28888 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 31004 0 1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 3036 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 4140 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_35
timestamp 1688980957
transform 1 0 5980 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_41
timestamp 1688980957
transform 1 0 6532 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_44
timestamp 1688980957
transform 1 0 6808 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_57
timestamp 1688980957
transform 1 0 8004 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_61
timestamp 1688980957
transform 1 0 8372 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_71
timestamp 1688980957
transform 1 0 9292 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_79
timestamp 1688980957
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_84
timestamp 1688980957
transform 1 0 10488 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_96
timestamp 1688980957
transform 1 0 11592 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_100
timestamp 1688980957
transform 1 0 11960 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_110
timestamp 1688980957
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_120
timestamp 1688980957
transform 1 0 13800 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_124
timestamp 1688980957
transform 1 0 14168 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_158
timestamp 1688980957
transform 1 0 17296 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 1688980957
transform 1 0 17940 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_178
timestamp 1688980957
transform 1 0 19136 0 -1 16864
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_192
timestamp 1688980957
transform 1 0 20424 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_204
timestamp 1688980957
transform 1 0 21528 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_210
timestamp 1688980957
transform 1 0 22080 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_219
timestamp 1688980957
transform 1 0 22908 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 23276 0 -1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 23460 0 -1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 24564 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_249
timestamp 1688980957
transform 1 0 25668 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_265
timestamp 1688980957
transform 1 0 27140 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_269
timestamp 1688980957
transform 1 0 27508 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 1688980957
transform 1 0 28244 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_281
timestamp 1688980957
transform 1 0 28612 0 -1 16864
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 3036 0 1 16864
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 4140 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 5244 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 5428 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_41
timestamp 1688980957
transform 1 0 6532 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_49
timestamp 1688980957
transform 1 0 7268 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_80
timestamp 1688980957
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1688980957
transform 1 0 10580 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_111
timestamp 1688980957
transform 1 0 12972 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_136
timestamp 1688980957
transform 1 0 15272 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_141
timestamp 1688980957
transform 1 0 15732 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 1688980957
transform 1 0 16100 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 20700 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_200
timestamp 1688980957
transform 1 0 21160 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_224
timestamp 1688980957
transform 1 0 23368 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_236
timestamp 1688980957
transform 1 0 24472 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_242
timestamp 1688980957
transform 1 0 25024 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_248
timestamp 1688980957
transform 1 0 25576 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_253
timestamp 1688980957
transform 1 0 26036 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_277
timestamp 1688980957
transform 1 0 28244 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_281
timestamp 1688980957
transform 1 0 28612 0 1 16864
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 3036 0 -1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 4140 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_27
timestamp 1688980957
transform 1 0 5244 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_35
timestamp 1688980957
transform 1 0 5980 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_100
timestamp 1688980957
transform 1 0 11960 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_157
timestamp 1688980957
transform 1 0 17204 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_210
timestamp 1688980957
transform 1 0 22080 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_222
timestamp 1688980957
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_225
timestamp 1688980957
transform 1 0 23460 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_281
timestamp 1688980957
transform 1 0 28612 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_285
timestamp 1688980957
transform 1 0 28980 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_289
timestamp 1688980957
transform 1 0 29348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_300
timestamp 1688980957
transform 1 0 30360 0 -1 17952
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 3036 0 1 17952
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 4140 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 5244 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_41
timestamp 1688980957
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_45
timestamp 1688980957
transform 1 0 6900 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_93
timestamp 1688980957
transform 1 0 11316 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_97
timestamp 1688980957
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_191
timestamp 1688980957
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 20700 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_197
timestamp 1688980957
transform 1 0 20884 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_223
timestamp 1688980957
transform 1 0 23276 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_232
timestamp 1688980957
transform 1 0 24104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_238
timestamp 1688980957
transform 1 0 24656 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_253
timestamp 1688980957
transform 1 0 26036 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_258
timestamp 1688980957
transform 1 0 26496 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_276
timestamp 1688980957
transform 1 0 28152 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_309
timestamp 1688980957
transform 1 0 31188 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_313
timestamp 1688980957
transform 1 0 31556 0 1 17952
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 3036 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_15
timestamp 1688980957
transform 1 0 4140 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_49
timestamp 1688980957
transform 1 0 7268 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_53
timestamp 1688980957
transform 1 0 7636 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1688980957
transform 1 0 8004 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_85
timestamp 1688980957
transform 1 0 10580 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_89
timestamp 1688980957
transform 1 0 10948 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_122
timestamp 1688980957
transform 1 0 13984 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_155
timestamp 1688980957
transform 1 0 17020 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 18124 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_169
timestamp 1688980957
transform 1 0 18308 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_178
timestamp 1688980957
transform 1 0 19136 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_200
timestamp 1688980957
transform 1 0 21160 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_206
timestamp 1688980957
transform 1 0 21712 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_214
timestamp 1688980957
transform 1 0 22448 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_218
timestamp 1688980957
transform 1 0 22816 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_225
timestamp 1688980957
transform 1 0 23460 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_260
timestamp 1688980957
transform 1 0 26680 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_270
timestamp 1688980957
transform 1 0 27600 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_274
timestamp 1688980957
transform 1 0 27968 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 28428 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_281
timestamp 1688980957
transform 1 0 28612 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_287
timestamp 1688980957
transform 1 0 29164 0 -1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_6
timestamp 1688980957
transform 1 0 3312 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1688980957
transform 1 0 4416 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1688980957
transform 1 0 5152 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 5428 0 1 19040
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 6532 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_53
timestamp 1688980957
transform 1 0 7636 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_63
timestamp 1688980957
transform 1 0 8556 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_74
timestamp 1688980957
transform 1 0 9568 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_78
timestamp 1688980957
transform 1 0 9936 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 10212 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_85
timestamp 1688980957
transform 1 0 10580 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_94
timestamp 1688980957
transform 1 0 11408 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_102
timestamp 1688980957
transform 1 0 12144 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_126
timestamp 1688980957
transform 1 0 14352 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_133
timestamp 1688980957
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_141
timestamp 1688980957
transform 1 0 15732 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_197
timestamp 1688980957
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_225
timestamp 1688980957
transform 1 0 23460 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 25852 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_260
timestamp 1688980957
transform 1 0 26680 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_264
timestamp 1688980957
transform 1 0 27048 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_282
timestamp 1688980957
transform 1 0 28704 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_286
timestamp 1688980957
transform 1 0 29072 0 1 19040
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 3036 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_15
timestamp 1688980957
transform 1 0 4140 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_41
timestamp 1688980957
transform 1 0 6532 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_45
timestamp 1688980957
transform 1 0 6900 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_49
timestamp 1688980957
transform 1 0 7268 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 7820 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_64
timestamp 1688980957
transform 1 0 8648 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_82
timestamp 1688980957
transform 1 0 10304 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_86
timestamp 1688980957
transform 1 0 10672 0 -1 20128
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_95
timestamp 1688980957
transform 1 0 11500 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_107
timestamp 1688980957
transform 1 0 12604 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 12972 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_120
timestamp 1688980957
transform 1 0 13800 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_140
timestamp 1688980957
transform 1 0 15640 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_144
timestamp 1688980957
transform 1 0 16008 0 -1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_148
timestamp 1688980957
transform 1 0 16376 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_160
timestamp 1688980957
transform 1 0 17480 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_172
timestamp 1688980957
transform 1 0 18584 0 -1 20128
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_180
timestamp 1688980957
transform 1 0 19320 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_208
timestamp 1688980957
transform 1 0 21896 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_212
timestamp 1688980957
transform 1 0 22264 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_225
timestamp 1688980957
transform 1 0 23460 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_241
timestamp 1688980957
transform 1 0 24932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_254
timestamp 1688980957
transform 1 0 26128 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_259
timestamp 1688980957
transform 1 0 26588 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 1688980957
transform 1 0 28336 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_293
timestamp 1688980957
transform 1 0 29716 0 -1 20128
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 3036 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_15
timestamp 1688980957
transform 1 0 4140 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_21
timestamp 1688980957
transform 1 0 4692 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_24
timestamp 1688980957
transform 1 0 4968 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_94
timestamp 1688980957
transform 1 0 11408 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_98
timestamp 1688980957
transform 1 0 11776 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_108
timestamp 1688980957
transform 1 0 12696 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_116
timestamp 1688980957
transform 1 0 13432 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_126
timestamp 1688980957
transform 1 0 14352 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_130
timestamp 1688980957
transform 1 0 14720 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_135
timestamp 1688980957
transform 1 0 15180 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 15548 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1688980957
transform 1 0 15732 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_145
timestamp 1688980957
transform 1 0 16100 0 1 20128
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_157
timestamp 1688980957
transform 1 0 17204 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_169
timestamp 1688980957
transform 1 0 18308 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1688980957
transform 1 0 20148 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 20700 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_197
timestamp 1688980957
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_219
timestamp 1688980957
transform 1 0 22908 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_242
timestamp 1688980957
transform 1 0 25024 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_256
timestamp 1688980957
transform 1 0 26312 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_300
timestamp 1688980957
transform 1 0 30360 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_304
timestamp 1688980957
transform 1 0 30728 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_309
timestamp 1688980957
transform 1 0 31188 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_313
timestamp 1688980957
transform 1 0 31556 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_13
timestamp 1688980957
transform 1 0 3956 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_24
timestamp 1688980957
transform 1 0 4968 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_35
timestamp 1688980957
transform 1 0 5980 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_45
timestamp 1688980957
transform 1 0 6900 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_53
timestamp 1688980957
transform 1 0 7636 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 8004 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_69
timestamp 1688980957
transform 1 0 9108 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_75
timestamp 1688980957
transform 1 0 9660 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_96
timestamp 1688980957
transform 1 0 11592 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 1688980957
transform 1 0 12880 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_113
timestamp 1688980957
transform 1 0 13156 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_140
timestamp 1688980957
transform 1 0 15640 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_144
timestamp 1688980957
transform 1 0 16008 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_150
timestamp 1688980957
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_154
timestamp 1688980957
transform 1 0 16928 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1688980957
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_200
timestamp 1688980957
transform 1 0 21160 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_215
timestamp 1688980957
transform 1 0 22540 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 23276 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_225
timestamp 1688980957
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 28336 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_305
timestamp 1688980957
transform 1 0 30820 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_313
timestamp 1688980957
transform 1 0 31556 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_3
timestamp 1688980957
transform 1 0 3036 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 5244 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_29
timestamp 1688980957
transform 1 0 5428 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_53
timestamp 1688980957
transform 1 0 7636 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_57
timestamp 1688980957
transform 1 0 8004 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_61
timestamp 1688980957
transform 1 0 8372 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1688980957
transform 1 0 10580 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_96
timestamp 1688980957
transform 1 0 11592 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_120
timestamp 1688980957
transform 1 0 13800 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_137
timestamp 1688980957
transform 1 0 15364 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_152
timestamp 1688980957
transform 1 0 16744 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_170
timestamp 1688980957
transform 1 0 18400 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_182
timestamp 1688980957
transform 1 0 19504 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_192
timestamp 1688980957
transform 1 0 20424 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_253
timestamp 1688980957
transform 1 0 26036 0 1 21216
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_283
timestamp 1688980957
transform 1 0 28796 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_295
timestamp 1688980957
transform 1 0 29900 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 31004 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_309
timestamp 1688980957
transform 1 0 31188 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_3
timestamp 1688980957
transform 1 0 3036 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_7
timestamp 1688980957
transform 1 0 3404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_66
timestamp 1688980957
transform 1 0 8832 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_70
timestamp 1688980957
transform 1 0 9200 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_76
timestamp 1688980957
transform 1 0 9752 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_137
timestamp 1688980957
transform 1 0 15364 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_141
timestamp 1688980957
transform 1 0 15732 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_162
timestamp 1688980957
transform 1 0 17664 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 18124 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_169
timestamp 1688980957
transform 1 0 18308 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_202
timestamp 1688980957
transform 1 0 21344 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_217
timestamp 1688980957
transform 1 0 22724 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_225
timestamp 1688980957
transform 1 0 23460 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_277
timestamp 1688980957
transform 1 0 28244 0 -1 22304
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 28612 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_293
timestamp 1688980957
transform 1 0 29716 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_19
timestamp 1688980957
transform 1 0 4508 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_23
timestamp 1688980957
transform 1 0 4876 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 5244 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_40
timestamp 1688980957
transform 1 0 6440 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 10212 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_85
timestamp 1688980957
transform 1 0 10580 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_89
timestamp 1688980957
transform 1 0 10948 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_98
timestamp 1688980957
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_152
timestamp 1688980957
transform 1 0 16744 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_187
timestamp 1688980957
transform 1 0 19964 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_214
timestamp 1688980957
transform 1 0 22448 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_243
timestamp 1688980957
transform 1 0 25116 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_274
timestamp 1688980957
transform 1 0 27968 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_278
timestamp 1688980957
transform 1 0 28336 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_292
timestamp 1688980957
transform 1 0 29624 0 1 22304
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_296
timestamp 1688980957
transform 1 0 29992 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_309
timestamp 1688980957
transform 1 0 31188 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_3
timestamp 1688980957
transform 1 0 3036 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_11
timestamp 1688980957
transform 1 0 3772 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_42
timestamp 1688980957
transform 1 0 6624 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_87
timestamp 1688980957
transform 1 0 10764 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_91
timestamp 1688980957
transform 1 0 11132 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_95
timestamp 1688980957
transform 1 0 11500 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_101
timestamp 1688980957
transform 1 0 12052 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_104
timestamp 1688980957
transform 1 0 12328 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_108
timestamp 1688980957
transform 1 0 12696 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_120
timestamp 1688980957
transform 1 0 13800 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_124
timestamp 1688980957
transform 1 0 14168 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_141
timestamp 1688980957
transform 1 0 15732 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_169
timestamp 1688980957
transform 1 0 18308 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1688980957
transform 1 0 23184 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_271
timestamp 1688980957
transform 1 0 27692 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 28428 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_313
timestamp 1688980957
transform 1 0 31556 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_3
timestamp 1688980957
transform 1 0 3036 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 5244 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_29
timestamp 1688980957
transform 1 0 5428 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_48
timestamp 1688980957
transform 1 0 7176 0 1 23392
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 10580 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_97
timestamp 1688980957
transform 1 0 11684 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_107
timestamp 1688980957
transform 1 0 12604 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_119
timestamp 1688980957
transform 1 0 13708 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_124
timestamp 1688980957
transform 1 0 14168 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 15548 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_141
timestamp 1688980957
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_152
timestamp 1688980957
transform 1 0 16744 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_162
timestamp 1688980957
transform 1 0 17664 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_166
timestamp 1688980957
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_185
timestamp 1688980957
transform 1 0 19780 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_189
timestamp 1688980957
transform 1 0 20148 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1688980957
transform 1 0 20516 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_197
timestamp 1688980957
transform 1 0 20884 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_206
timestamp 1688980957
transform 1 0 21712 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_218
timestamp 1688980957
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_223
timestamp 1688980957
transform 1 0 23276 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_265
timestamp 1688980957
transform 1 0 27140 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_273
timestamp 1688980957
transform 1 0 27876 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_281
timestamp 1688980957
transform 1 0 28612 0 1 23392
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_290
timestamp 1688980957
transform 1 0 29440 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_302
timestamp 1688980957
transform 1 0 30544 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_309
timestamp 1688980957
transform 1 0 31188 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_3
timestamp 1688980957
transform 1 0 3036 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_36
timestamp 1688980957
transform 1 0 6072 0 -1 24480
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_44
timestamp 1688980957
transform 1 0 6808 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_57
timestamp 1688980957
transform 1 0 8004 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_92
timestamp 1688980957
transform 1 0 11224 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_97
timestamp 1688980957
transform 1 0 11684 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_101
timestamp 1688980957
transform 1 0 12052 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_113
timestamp 1688980957
transform 1 0 13156 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_161
timestamp 1688980957
transform 1 0 17572 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_165
timestamp 1688980957
transform 1 0 17940 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_179
timestamp 1688980957
transform 1 0 19228 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_183
timestamp 1688980957
transform 1 0 19596 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_187
timestamp 1688980957
transform 1 0 19964 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_199
timestamp 1688980957
transform 1 0 21068 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_207
timestamp 1688980957
transform 1 0 21804 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 22724 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 23276 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_225
timestamp 1688980957
transform 1 0 23460 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_244
timestamp 1688980957
transform 1 0 25208 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_251
timestamp 1688980957
transform 1 0 25852 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_264
timestamp 1688980957
transform 1 0 27048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_276
timestamp 1688980957
transform 1 0 28152 0 -1 24480
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_289
timestamp 1688980957
transform 1 0 29348 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_301
timestamp 1688980957
transform 1 0 30452 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_19
timestamp 1688980957
transform 1 0 4508 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_29
timestamp 1688980957
transform 1 0 5428 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_50
timestamp 1688980957
transform 1 0 7360 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_79
timestamp 1688980957
transform 1 0 10028 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_102
timestamp 1688980957
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_135
timestamp 1688980957
transform 1 0 15180 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_150
timestamp 1688980957
transform 1 0 16560 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_154
timestamp 1688980957
transform 1 0 16928 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_158
timestamp 1688980957
transform 1 0 17296 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_191
timestamp 1688980957
transform 1 0 20332 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 20700 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 20884 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_209
timestamp 1688980957
transform 1 0 21988 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_213
timestamp 1688980957
transform 1 0 22356 0 1 24480
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_225
timestamp 1688980957
transform 1 0 23460 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_237
timestamp 1688980957
transform 1 0 24564 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_249
timestamp 1688980957
transform 1 0 25668 0 1 24480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 26036 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_265
timestamp 1688980957
transform 1 0 27140 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_269
timestamp 1688980957
transform 1 0 27508 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_300
timestamp 1688980957
transform 1 0 30360 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_309
timestamp 1688980957
transform 1 0 31188 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_3
timestamp 1688980957
transform 1 0 3036 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_15
timestamp 1688980957
transform 1 0 4140 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_40
timestamp 1688980957
transform 1 0 6440 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_44
timestamp 1688980957
transform 1 0 6808 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_48
timestamp 1688980957
transform 1 0 7176 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_52
timestamp 1688980957
transform 1 0 7544 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_66
timestamp 1688980957
transform 1 0 8832 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_70
timestamp 1688980957
transform 1 0 9200 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_164
timestamp 1688980957
transform 1 0 17848 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_169
timestamp 1688980957
transform 1 0 18308 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_205
timestamp 1688980957
transform 1 0 21620 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_251
timestamp 1688980957
transform 1 0 25852 0 -1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_260
timestamp 1688980957
transform 1 0 26680 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_272
timestamp 1688980957
transform 1 0 27784 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_281
timestamp 1688980957
transform 1 0 28612 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_293
timestamp 1688980957
transform 1 0 29716 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_3
timestamp 1688980957
transform 1 0 3036 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_7
timestamp 1688980957
transform 1 0 3404 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 1688980957
transform 1 0 5428 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_33
timestamp 1688980957
transform 1 0 5796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_39
timestamp 1688980957
transform 1 0 6348 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_79
timestamp 1688980957
transform 1 0 10028 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 10396 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_85
timestamp 1688980957
transform 1 0 10580 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_97
timestamp 1688980957
transform 1 0 11684 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_101
timestamp 1688980957
transform 1 0 12052 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1688980957
transform 1 0 15456 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_164
timestamp 1688980957
transform 1 0 17848 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_168
timestamp 1688980957
transform 1 0 18216 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1688980957
transform 1 0 20608 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_208
timestamp 1688980957
transform 1 0 21896 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_230
timestamp 1688980957
transform 1 0 23920 0 1 25568
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_257
timestamp 1688980957
transform 1 0 26404 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_292
timestamp 1688980957
transform 1 0 29624 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_296
timestamp 1688980957
transform 1 0 29992 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_302
timestamp 1688980957
transform 1 0 30544 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_309
timestamp 1688980957
transform 1 0 31188 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_27
timestamp 1688980957
transform 1 0 5244 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_51
timestamp 1688980957
transform 1 0 7452 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_73
timestamp 1688980957
transform 1 0 9476 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_77
timestamp 1688980957
transform 1 0 9844 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_81
timestamp 1688980957
transform 1 0 10212 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_88
timestamp 1688980957
transform 1 0 10856 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_92
timestamp 1688980957
transform 1 0 11224 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_100
timestamp 1688980957
transform 1 0 11960 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_104
timestamp 1688980957
transform 1 0 12328 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_113
timestamp 1688980957
transform 1 0 13156 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_123
timestamp 1688980957
transform 1 0 14076 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_136
timestamp 1688980957
transform 1 0 15272 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_140
timestamp 1688980957
transform 1 0 15640 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_146
timestamp 1688980957
transform 1 0 16192 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_172
timestamp 1688980957
transform 1 0 18584 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_202
timestamp 1688980957
transform 1 0 21344 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_245
timestamp 1688980957
transform 1 0 25300 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_263
timestamp 1688980957
transform 1 0 26956 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_307
timestamp 1688980957
transform 1 0 31004 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_315
timestamp 1688980957
transform 1 0 31740 0 -1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 3036 0 1 26656
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 4140 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 5244 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 5428 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_41
timestamp 1688980957
transform 1 0 6532 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_45
timestamp 1688980957
transform 1 0 6900 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_81
timestamp 1688980957
transform 1 0 10212 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_85
timestamp 1688980957
transform 1 0 10580 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_94
timestamp 1688980957
transform 1 0 11408 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_98
timestamp 1688980957
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_102
timestamp 1688980957
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_106
timestamp 1688980957
transform 1 0 12512 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_118
timestamp 1688980957
transform 1 0 13616 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_130
timestamp 1688980957
transform 1 0 14720 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 1688980957
transform 1 0 15732 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_145
timestamp 1688980957
transform 1 0 16100 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_149
timestamp 1688980957
transform 1 0 16468 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_159
timestamp 1688980957
transform 1 0 17388 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_167
timestamp 1688980957
transform 1 0 18124 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 20148 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 20700 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_197
timestamp 1688980957
transform 1 0 20884 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_201
timestamp 1688980957
transform 1 0 21252 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_231
timestamp 1688980957
transform 1 0 24012 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_309
timestamp 1688980957
transform 1 0 31188 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_19
timestamp 1688980957
transform 1 0 4508 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_23
timestamp 1688980957
transform 1 0 4876 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_27
timestamp 1688980957
transform 1 0 5244 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_31
timestamp 1688980957
transform 1 0 5612 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_39
timestamp 1688980957
transform 1 0 6348 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 7820 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_57
timestamp 1688980957
transform 1 0 8004 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_77
timestamp 1688980957
transform 1 0 9844 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_107
timestamp 1688980957
transform 1 0 12604 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 12972 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_113
timestamp 1688980957
transform 1 0 13156 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_118
timestamp 1688980957
transform 1 0 13616 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_150
timestamp 1688980957
transform 1 0 16560 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_165
timestamp 1688980957
transform 1 0 17940 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_169
timestamp 1688980957
transform 1 0 18308 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_173
timestamp 1688980957
transform 1 0 18676 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_195
timestamp 1688980957
transform 1 0 20700 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_203
timestamp 1688980957
transform 1 0 21436 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_254
timestamp 1688980957
transform 1 0 26128 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_264
timestamp 1688980957
transform 1 0 27048 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1688980957
transform 1 0 28336 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_284
timestamp 1688980957
transform 1 0 28888 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_294
timestamp 1688980957
transform 1 0 29808 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_315
timestamp 1688980957
transform 1 0 31740 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_3
timestamp 1688980957
transform 1 0 3036 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_38
timestamp 1688980957
transform 1 0 6256 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_42
timestamp 1688980957
transform 1 0 6624 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_46
timestamp 1688980957
transform 1 0 6992 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_69
timestamp 1688980957
transform 1 0 9108 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_79
timestamp 1688980957
transform 1 0 10028 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_85
timestamp 1688980957
transform 1 0 10580 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_116
timestamp 1688980957
transform 1 0 13432 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_152
timestamp 1688980957
transform 1 0 16744 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_156
timestamp 1688980957
transform 1 0 17112 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_185
timestamp 1688980957
transform 1 0 19780 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1688980957
transform 1 0 20516 0 1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 20884 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_209
timestamp 1688980957
transform 1 0 21988 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 1688980957
transform 1 0 25668 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_268
timestamp 1688980957
transform 1 0 27416 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_3
timestamp 1688980957
transform 1 0 3036 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_11
timestamp 1688980957
transform 1 0 3772 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_41
timestamp 1688980957
transform 1 0 6532 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_47
timestamp 1688980957
transform 1 0 7084 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_77
timestamp 1688980957
transform 1 0 9844 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 12972 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_113
timestamp 1688980957
transform 1 0 13156 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_119
timestamp 1688980957
transform 1 0 13708 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_148
timestamp 1688980957
transform 1 0 16376 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_152
timestamp 1688980957
transform 1 0 16744 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_164
timestamp 1688980957
transform 1 0 17848 0 -1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 18308 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_181
timestamp 1688980957
transform 1 0 19412 0 -1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 20516 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_205
timestamp 1688980957
transform 1 0 21620 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_213
timestamp 1688980957
transform 1 0 22356 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_218
timestamp 1688980957
transform 1 0 22816 0 -1 28832
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_239
timestamp 1688980957
transform 1 0 24748 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_251
timestamp 1688980957
transform 1 0 25852 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_259
timestamp 1688980957
transform 1 0 26588 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_276
timestamp 1688980957
transform 1 0 28152 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_316
timestamp 1688980957
transform 1 0 31832 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_3
timestamp 1688980957
transform 1 0 3036 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_7
timestamp 1688980957
transform 1 0 3404 0 1 28832
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_32
timestamp 1688980957
transform 1 0 5704 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_44
timestamp 1688980957
transform 1 0 6808 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_52
timestamp 1688980957
transform 1 0 7544 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_56
timestamp 1688980957
transform 1 0 7912 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_74
timestamp 1688980957
transform 1 0 9568 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_78
timestamp 1688980957
transform 1 0 9936 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_85
timestamp 1688980957
transform 1 0 10580 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_90
timestamp 1688980957
transform 1 0 11040 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_107
timestamp 1688980957
transform 1 0 12604 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 15548 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_144
timestamp 1688980957
transform 1 0 16008 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_154
timestamp 1688980957
transform 1 0 16928 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_176
timestamp 1688980957
transform 1 0 18952 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 1688980957
transform 1 0 20516 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_197
timestamp 1688980957
transform 1 0 20884 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_205
timestamp 1688980957
transform 1 0 21620 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_235
timestamp 1688980957
transform 1 0 24380 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_239
timestamp 1688980957
transform 1 0 24748 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1688980957
transform 1 0 25300 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 25852 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_270
timestamp 1688980957
transform 1 0 27600 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_283
timestamp 1688980957
transform 1 0 28796 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 31004 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_315
timestamp 1688980957
transform 1 0 31740 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_22
timestamp 1688980957
transform 1 0 4784 0 -1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_26
timestamp 1688980957
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_38
timestamp 1688980957
transform 1 0 6256 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_50
timestamp 1688980957
transform 1 0 7360 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_77
timestamp 1688980957
transform 1 0 9844 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_81
timestamp 1688980957
transform 1 0 10212 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_102
timestamp 1688980957
transform 1 0 12144 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_113
timestamp 1688980957
transform 1 0 13156 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_134
timestamp 1688980957
transform 1 0 15088 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_138
timestamp 1688980957
transform 1 0 15456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 18124 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_180
timestamp 1688980957
transform 1 0 19320 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_202
timestamp 1688980957
transform 1 0 21344 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_206
timestamp 1688980957
transform 1 0 21712 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_214
timestamp 1688980957
transform 1 0 22448 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_219
timestamp 1688980957
transform 1 0 22908 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 28428 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_281
timestamp 1688980957
transform 1 0 28612 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_291
timestamp 1688980957
transform 1 0 29532 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_19
timestamp 1688980957
transform 1 0 4508 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 5244 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 5428 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 6532 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_53
timestamp 1688980957
transform 1 0 7636 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_62
timestamp 1688980957
transform 1 0 8464 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_68
timestamp 1688980957
transform 1 0 9016 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 9844 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 10396 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_105
timestamp 1688980957
transform 1 0 12420 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1688980957
transform 1 0 15456 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_141
timestamp 1688980957
transform 1 0 15732 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_156
timestamp 1688980957
transform 1 0 17112 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_180
timestamp 1688980957
transform 1 0 19320 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 20700 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_312
timestamp 1688980957
transform 1 0 31464 0 1 29920
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_29
timestamp 1688980957
transform 1 0 5428 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_41
timestamp 1688980957
transform 1 0 6532 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_53
timestamp 1688980957
transform 1 0 7636 0 -1 31008
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 8004 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 9108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_81
timestamp 1688980957
transform 1 0 10212 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_108
timestamp 1688980957
transform 1 0 12696 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_113
timestamp 1688980957
transform 1 0 13156 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_135
timestamp 1688980957
transform 1 0 15180 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_161
timestamp 1688980957
transform 1 0 17572 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_165
timestamp 1688980957
transform 1 0 17940 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_169
timestamp 1688980957
transform 1 0 18308 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_211
timestamp 1688980957
transform 1 0 22172 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_220
timestamp 1688980957
transform 1 0 23000 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_225
timestamp 1688980957
transform 1 0 23460 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_232
timestamp 1688980957
transform 1 0 24104 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_236
timestamp 1688980957
transform 1 0 24472 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_248
timestamp 1688980957
transform 1 0 25576 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_252
timestamp 1688980957
transform 1 0 25944 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_278
timestamp 1688980957
transform 1 0 28336 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_284
timestamp 1688980957
transform 1 0 28888 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_19
timestamp 1688980957
transform 1 0 4508 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 5244 0 1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 5428 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 6532 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 7636 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 8740 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 9844 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 10396 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_85
timestamp 1688980957
transform 1 0 10580 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_106
timestamp 1688980957
transform 1 0 12512 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_110
timestamp 1688980957
transform 1 0 12880 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 15456 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_141
timestamp 1688980957
transform 1 0 15732 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_152
timestamp 1688980957
transform 1 0 16744 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_168
timestamp 1688980957
transform 1 0 18216 0 1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_172
timestamp 1688980957
transform 1 0 18584 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_184
timestamp 1688980957
transform 1 0 19688 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_197
timestamp 1688980957
transform 1 0 20884 0 1 31008
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_204
timestamp 1688980957
transform 1 0 21528 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_216
timestamp 1688980957
transform 1 0 22632 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_224
timestamp 1688980957
transform 1 0 23368 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_231
timestamp 1688980957
transform 1 0 24012 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_243
timestamp 1688980957
transform 1 0 25116 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_272
timestamp 1688980957
transform 1 0 27784 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_309
timestamp 1688980957
transform 1 0 31188 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_6
timestamp 1688980957
transform 1 0 3312 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_48
timestamp 1688980957
transform 1 0 7176 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_57
timestamp 1688980957
transform 1 0 8004 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_61
timestamp 1688980957
transform 1 0 8372 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_81
timestamp 1688980957
transform 1 0 10212 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_85
timestamp 1688980957
transform 1 0 10580 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_93
timestamp 1688980957
transform 1 0 11316 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_113
timestamp 1688980957
transform 1 0 13156 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_121
timestamp 1688980957
transform 1 0 13892 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_141
timestamp 1688980957
transform 1 0 15732 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_145
timestamp 1688980957
transform 1 0 16100 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_165
timestamp 1688980957
transform 1 0 17940 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_169
timestamp 1688980957
transform 1 0 18308 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_173
timestamp 1688980957
transform 1 0 18676 0 -1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_177
timestamp 1688980957
transform 1 0 19044 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_189
timestamp 1688980957
transform 1 0 20148 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_195
timestamp 1688980957
transform 1 0 20700 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_216
timestamp 1688980957
transform 1 0 22632 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_225
timestamp 1688980957
transform 1 0 23460 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_229
timestamp 1688980957
transform 1 0 23828 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_256
timestamp 1688980957
transform 1 0 26312 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_274
timestamp 1688980957
transform 1 0 27968 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_307
timestamp 1688980957
transform 1 0 31004 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_309
timestamp 1688980957
transform 1 0 31188 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_313
timestamp 1688980957
transform 1 0 31556 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31924 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 9844 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform 1 0 7912 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 8832 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 6348 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 17204 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 16468 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 25760 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 25484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 16652 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 15640 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 16468 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 15272 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform 1 0 24104 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 24196 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 25116 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 22540 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 21896 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 19964 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 17480 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 19412 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 21344 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 20240 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 20976 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 20792 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform 1 0 16652 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 15640 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform -1 0 25024 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 24748 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 21712 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 21712 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 21620 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 21344 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 21344 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 20792 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 22172 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 22540 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 6256 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 7820 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 18308 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 17480 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 17940 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 17020 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 21344 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 19780 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 19780 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 20424 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold48
timestamp 1688980957
transform -1 0 27508 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 24196 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 23460 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 19596 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform -1 0 18860 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform 1 0 17480 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform 1 0 16744 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold55
timestamp 1688980957
transform -1 0 15640 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform 1 0 7176 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold57
timestamp 1688980957
transform -1 0 26588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform 1 0 25116 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 24564 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform 1 0 22540 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 12236 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 13708 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 14536 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 13616 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold65 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20332 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 11316 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 25208 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 26404 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform 1 0 26864 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform 1 0 27416 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform 1 0 22724 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform 1 0 24748 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform -1 0 6716 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 4600 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 9200 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform -1 0 8280 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 19228 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 20700 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform 1 0 24196 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 24196 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform 1 0 4600 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 5980 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 20240 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform -1 0 19320 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 15732 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 16744 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 24472 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 23736 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 20424 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform 1 0 19320 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold91 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13984 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 14260 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 15548 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform -1 0 17020 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 15732 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold96
timestamp 1688980957
transform -1 0 12880 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 15732 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform -1 0 17204 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 16008 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform 1 0 4600 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 6992 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 17664 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 16008 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 7360 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform 1 0 18124 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 17480 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 30820 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform 1 0 29348 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 16192 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold111
timestamp 1688980957
transform 1 0 27048 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 24380 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 22448 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold114
timestamp 1688980957
transform 1 0 18676 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform 1 0 5980 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 6164 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform -1 0 15180 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 13708 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 8740 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform -1 0 7912 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform -1 0 10028 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform -1 0 17204 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 16468 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform -1 0 7176 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 6440 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 22356 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 21620 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 6900 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform -1 0 5980 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform 1 0 9292 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 9292 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform 1 0 5336 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold133
timestamp 1688980957
transform -1 0 17756 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  hold134
timestamp 1688980957
transform 1 0 16376 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 17388 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform 1 0 16192 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 18216 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform 1 0 19688 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 21160 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 11868 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform -1 0 11040 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold142
timestamp 1688980957
transform 1 0 11776 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 13340 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform -1 0 14812 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 6624 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform -1 0 5336 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 8832 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform -1 0 10028 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold149
timestamp 1688980957
transform -1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform 1 0 13984 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform -1 0 15456 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform -1 0 21160 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform -1 0 21160 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 10028 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform 1 0 8096 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform -1 0 9568 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 17112 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform -1 0 19044 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 13340 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform 1 0 12328 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold161 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform -1 0 9936 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold163
timestamp 1688980957
transform -1 0 18676 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform 1 0 4508 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform 1 0 3496 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform 1 0 7912 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold167
timestamp 1688980957
transform -1 0 16468 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform -1 0 19780 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform -1 0 22816 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 9844 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 11316 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold172
timestamp 1688980957
transform -1 0 24748 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform 1 0 18952 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold174
timestamp 1688980957
transform -1 0 21620 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform 1 0 7084 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform 1 0 10948 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold177
timestamp 1688980957
transform -1 0 12512 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform 1 0 12788 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 14720 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform -1 0 8924 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 6992 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform -1 0 7268 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 9568 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform 1 0 7176 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold185
timestamp 1688980957
transform 1 0 14628 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 15180 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 11316 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform -1 0 31924 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform -1 0 31924 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform -1 0 14260 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform 1 0 9844 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform 1 0 7820 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 12604 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform 1 0 10120 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 30820 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 30084 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform -1 0 11776 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform 1 0 3772 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform 1 0 27876 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 28428 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold201
timestamp 1688980957
transform -1 0 27876 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform -1 0 27508 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform -1 0 7360 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform 1 0 3404 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform 1 0 14444 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold206
timestamp 1688980957
transform -1 0 16836 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform 1 0 16560 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform -1 0 14996 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform 1 0 10764 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold210
timestamp 1688980957
transform 1 0 25300 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform -1 0 25300 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 25576 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 25944 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform -1 0 30728 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform -1 0 30452 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform -1 0 12880 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold217 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31004 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 29532 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold219
timestamp 1688980957
transform -1 0 30728 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform 1 0 29256 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform -1 0 21344 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold222
timestamp 1688980957
transform 1 0 29348 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform -1 0 28612 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold224
timestamp 1688980957
transform -1 0 18216 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform -1 0 16928 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform 1 0 24196 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 23368 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform -1 0 14168 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold229
timestamp 1688980957
transform -1 0 27692 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform -1 0 25852 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold231
timestamp 1688980957
transform 1 0 23828 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform -1 0 24196 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold233
timestamp 1688980957
transform 1 0 23460 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform -1 0 23460 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 23000 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform 1 0 23736 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform 1 0 24932 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform 1 0 25944 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 25484 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform -1 0 25116 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 29348 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold242
timestamp 1688980957
transform 1 0 14904 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold243
timestamp 1688980957
transform 1 0 30084 0 -1 32096
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform -1 0 27600 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold245
timestamp 1688980957
transform 1 0 26404 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform 1 0 26036 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform -1 0 31924 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform -1 0 29348 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform -1 0 27048 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform -1 0 23000 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 31924 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold252
timestamp 1688980957
transform 1 0 30820 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold253
timestamp 1688980957
transform -1 0 30820 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold254
timestamp 1688980957
transform 1 0 26680 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold255
timestamp 1688980957
transform -1 0 25944 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform 1 0 3680 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform -1 0 20056 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold258
timestamp 1688980957
transform -1 0 27784 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold259
timestamp 1688980957
transform -1 0 30176 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform -1 0 7820 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold261
timestamp 1688980957
transform -1 0 11316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform -1 0 9936 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold263
timestamp 1688980957
transform -1 0 21436 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform -1 0 20056 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold265
timestamp 1688980957
transform -1 0 16468 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold266
timestamp 1688980957
transform -1 0 28060 0 -1 27744
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold267
timestamp 1688980957
transform -1 0 27048 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold268
timestamp 1688980957
transform 1 0 27692 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform -1 0 28612 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold270
timestamp 1688980957
transform 1 0 23828 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform -1 0 24196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold272
timestamp 1688980957
transform -1 0 17848 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform 1 0 15916 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold274
timestamp 1688980957
transform 1 0 22264 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform -1 0 24196 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold276
timestamp 1688980957
transform -1 0 6532 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform 1 0 27600 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold278
timestamp 1688980957
transform -1 0 27600 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform -1 0 27232 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform -1 0 27876 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold281
timestamp 1688980957
transform -1 0 25944 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold282
timestamp 1688980957
transform -1 0 31556 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold283
timestamp 1688980957
transform 1 0 28612 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold284
timestamp 1688980957
transform -1 0 30820 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform -1 0 24932 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold286
timestamp 1688980957
transform 1 0 31188 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform -1 0 31096 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform -1 0 30084 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold289
timestamp 1688980957
transform -1 0 28612 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform -1 0 31924 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold291
timestamp 1688980957
transform 1 0 29716 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform -1 0 31464 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform -1 0 28336 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold294
timestamp 1688980957
transform 1 0 28612 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform -1 0 28612 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold296
timestamp 1688980957
transform 1 0 24012 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1688980957
transform -1 0 22540 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold298
timestamp 1688980957
transform 1 0 31188 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform -1 0 28244 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform -1 0 25668 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold301
timestamp 1688980957
transform -1 0 29716 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold302
timestamp 1688980957
transform -1 0 24564 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold303
timestamp 1688980957
transform -1 0 19136 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform 1 0 14904 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 25392 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform 1 0 23644 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold307
timestamp 1688980957
transform -1 0 16836 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform 1 0 11408 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold309
timestamp 1688980957
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform 1 0 31188 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform 1 0 18308 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform -1 0 29348 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold313
timestamp 1688980957
transform -1 0 28336 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform 1 0 26772 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold315
timestamp 1688980957
transform -1 0 19044 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform -1 0 19228 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold317
timestamp 1688980957
transform -1 0 24104 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform 1 0 19412 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold319
timestamp 1688980957
transform 1 0 24380 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform 1 0 10672 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold321
timestamp 1688980957
transform 1 0 14168 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform -1 0 28980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold323
timestamp 1688980957
transform 1 0 17480 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform -1 0 18860 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1688980957
transform -1 0 30452 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform -1 0 31924 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1688980957
transform -1 0 31924 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 31924 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1688980957
transform -1 0 31924 0 -1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 6900 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1688980957
transform 1 0 3036 0 -1 21216
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform -1 0 31924 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform -1 0 19044 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 26036 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 4508 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 3036 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 3036 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 17664 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform -1 0 31924 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 3036 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 31188 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 3036 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 27508 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform -1 0 13892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform -1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 31648 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 3312 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 9752 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 29348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform -1 0 31924 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform -1 0 31924 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform -1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1688980957
transform 1 0 4508 0 -1 31008
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform -1 0 31648 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform -1 0 10212 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform -1 0 31924 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  max_cap95
timestamp 1688980957
transform 1 0 26036 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output37 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26036 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 1688980957
transform 1 0 16192 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output39
timestamp 1688980957
transform -1 0 15640 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output40
timestamp 1688980957
transform 1 0 30452 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output41
timestamp 1688980957
transform -1 0 4508 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output42
timestamp 1688980957
transform -1 0 4508 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output43
timestamp 1688980957
transform -1 0 4508 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output44
timestamp 1688980957
transform 1 0 11592 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output45
timestamp 1688980957
transform 1 0 30452 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output46
timestamp 1688980957
transform -1 0 4508 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output47
timestamp 1688980957
transform 1 0 30452 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output48
timestamp 1688980957
transform -1 0 9476 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output49
timestamp 1688980957
transform 1 0 28980 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output50
timestamp 1688980957
transform -1 0 4508 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output51
timestamp 1688980957
transform -1 0 4508 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output52
timestamp 1688980957
transform 1 0 23920 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 1688980957
transform 1 0 30360 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 1688980957
transform 1 0 29624 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 1688980957
transform -1 0 4508 0 1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 1688980957
transform 1 0 26036 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 1688980957
transform -1 0 4508 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 1688980957
transform 1 0 3036 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 1688980957
transform 1 0 12972 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 1688980957
transform 1 0 16744 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 1688980957
transform -1 0 4508 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 1688980957
transform 1 0 19320 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1688980957
transform 1 0 11592 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1688980957
transform 1 0 20884 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1688980957
transform 1 0 30452 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1688980957
transform 1 0 3036 0 1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1688980957
transform -1 0 6072 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1688980957
transform -1 0 4508 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1688980957
transform 1 0 28152 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1688980957
transform 1 0 26496 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1688980957
transform -1 0 15640 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1688980957
transform 1 0 30452 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1688980957
transform 1 0 28888 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1688980957
transform -1 0 6900 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1688980957
transform 1 0 30452 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1688980957
transform -1 0 7360 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1688980957
transform 1 0 10396 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1688980957
transform -1 0 4508 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1688980957
transform 1 0 30452 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1688980957
transform -1 0 18216 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1688980957
transform 1 0 29624 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1688980957
transform 1 0 28612 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1688980957
transform 1 0 3864 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1688980957
transform -1 0 9936 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1688980957
transform 1 0 23460 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1688980957
transform -1 0 4508 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1688980957
transform -1 0 4508 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1688980957
transform 1 0 30452 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 32200 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 2760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 32200 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 2760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 32200 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 2760 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 32200 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 2760 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 32200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 2760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 32200 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 2760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 32200 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 2760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 32200 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 2760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 32200 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 2760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 32200 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 2760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 32200 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 2760 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 32200 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 32200 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 2760 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 32200 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 2760 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 32200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 2760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 32200 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 2760 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 32200 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 2760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 32200 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 32200 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 2760 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 32200 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 32200 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 2760 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 32200 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 2760 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 32200 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 2760 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 32200 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 2760 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 32200 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 2760 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 32200 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 2760 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 32200 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 2760 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 32200 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 2760 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 32200 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 2760 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 32200 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 2760 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 32200 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 2760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 32200 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 2760 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 32200 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 2760 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 32200 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 2760 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 32200 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 2760 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 32200 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 2760 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 32200 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 2760 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 32200 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 2760 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 32200 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 2760 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 32200 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 2760 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 32200 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 2760 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 32200 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 2760 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 32200 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 2760 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 32200 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 2760 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 32200 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 2760 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 32200 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 2760 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 32200 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 2760 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 32200 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 2760 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 32200 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 2760 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 32200 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 2760 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 32200 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 2760 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 32200 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 2760 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 32200 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 2760 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 32200 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108 Downloads/unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 7912 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 10488 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 13064 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 15640 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 23368 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 25944 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 28520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 31096 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 13064 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 18216 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 23368 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 5336 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 10488 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 15640 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 20792 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 25944 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 31096 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 7912 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 13064 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 18216 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 23368 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 5336 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 10488 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 20792 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 25944 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 31096 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 7912 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 13064 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 18216 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 23368 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 5336 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 10488 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 15640 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 25944 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 31096 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 13064 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 18216 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 23368 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 5336 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 20792 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 25944 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 31096 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 13064 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 18216 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 23368 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 5336 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 10488 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 15640 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 25944 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 31096 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 7912 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 13064 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 18216 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 23368 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 5336 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 10488 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 15640 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 25944 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 31096 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13064 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 18216 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 23368 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 5336 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 10488 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 25944 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 31096 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 13064 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 23368 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 5336 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 10488 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 15640 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 25944 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 31096 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 13064 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 18216 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 23368 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 28520 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 5336 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 15640 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 20792 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 25944 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 31096 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 13064 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 23368 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 28520 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 5336 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 15640 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 25944 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 31096 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 7912 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 13064 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 23368 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 28520 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 5336 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 10488 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 15640 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 25944 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 31096 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 13064 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 18216 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 23368 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 28520 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 5336 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 10488 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 15640 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 20792 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 25944 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 31096 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13064 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 18216 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 23368 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 28520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 5336 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 10488 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 15640 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 25944 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 31096 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 13064 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 23368 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 28520 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 5336 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 10488 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 15640 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 25944 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 31096 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 7912 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 13064 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 18216 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 23368 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 28520 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 5336 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 10488 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 15640 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 25944 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 31096 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 7912 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13064 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 23368 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 28520 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 5336 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 10488 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 15640 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 25944 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 31096 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 7912 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 13064 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 18216 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 23368 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 28520 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 5336 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 10488 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 15640 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 20792 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 25944 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 31096 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 7912 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 13064 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 23368 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 28520 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 5336 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 10488 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 15640 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 20792 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 25944 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 31096 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 7912 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 13064 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 18216 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 23368 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 28520 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 5336 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 10488 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 15640 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 20792 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 25944 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 31096 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 7912 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13064 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 18216 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 23368 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 28520 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 5336 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 10488 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 15640 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 20792 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 25944 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 31096 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 7912 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 13064 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 23368 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 28520 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 5336 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 10488 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 15640 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 20792 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 25944 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 31096 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 7912 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 13064 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 18216 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 23368 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 28520 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 5336 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 10488 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 15640 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 20792 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 25944 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 31096 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 7912 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 13064 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 18216 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 23368 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 28520 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 5336 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 10488 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 15640 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 20792 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 25944 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 31096 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 7912 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 13064 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 18216 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 23368 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 28520 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 5336 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 10488 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 15640 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 20792 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 25944 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 31096 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 7912 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 13064 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 18216 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 23368 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 28520 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 5336 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 10488 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 15640 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 20792 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 25944 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 31096 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 7912 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 13064 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 18216 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 23368 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 28520 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 5336 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 10488 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 15640 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 20792 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 25944 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 31096 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 5336 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 7912 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 10488 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 13064 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 15640 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 18216 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 23368 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 25944 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 28520 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 31096 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  wire94
timestamp 1688980957
transform -1 0 16100 0 1 16864
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 34168 28568 34968 28688 0 FreeSans 480 0 0 0 i_start_rx
port 1 nsew signal input
flabel metal3 s 34168 6128 34968 6248 0 FreeSans 480 0 0 0 i_uart_rx
port 2 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 o_uart_tx
port 3 nsew signal tristate
flabel metal3 s 34168 27208 34968 27328 0 FreeSans 480 0 0 0 rst
port 4 nsew signal input
flabel metal4 s 6280 2672 6600 32144 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 13640 2672 13960 32144 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 21000 2672 21320 32144 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 28360 2672 28680 32144 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 6940 2672 7260 32144 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 14300 2672 14620 32144 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 21660 2672 21980 32144 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 29020 2672 29340 32144 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal3 s 34168 20408 34968 20528 0 FreeSans 480 0 0 0 wb_ack_i
port 7 nsew signal input
flabel metal2 s 16118 33544 16174 34344 0 FreeSans 224 90 0 0 wb_adr_o[0]
port 8 nsew signal tristate
flabel metal2 s 14186 33544 14242 34344 0 FreeSans 224 90 0 0 wb_adr_o[10]
port 9 nsew signal tristate
flabel metal3 s 34168 12248 34968 12368 0 FreeSans 480 0 0 0 wb_adr_o[11]
port 10 nsew signal tristate
flabel metal2 s 1950 33544 2006 34344 0 FreeSans 224 90 0 0 wb_adr_o[12]
port 11 nsew signal tristate
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 wb_adr_o[13]
port 12 nsew signal tristate
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 wb_adr_o[14]
port 13 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wb_adr_o[15]
port 14 nsew signal tristate
flabel metal3 s 34168 25168 34968 25288 0 FreeSans 480 0 0 0 wb_adr_o[1]
port 15 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 wb_adr_o[2]
port 16 nsew signal tristate
flabel metal3 s 34168 22448 34968 22568 0 FreeSans 480 0 0 0 wb_adr_o[3]
port 17 nsew signal tristate
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 wb_adr_o[4]
port 18 nsew signal tristate
flabel metal2 s 32862 33544 32918 34344 0 FreeSans 224 90 0 0 wb_adr_o[5]
port 19 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 wb_adr_o[6]
port 20 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 wb_adr_o[7]
port 21 nsew signal tristate
flabel metal2 s 23846 33544 23902 34344 0 FreeSans 224 90 0 0 wb_adr_o[8]
port 22 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 wb_adr_o[9]
port 23 nsew signal tristate
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 wb_cyc_o
port 24 nsew signal tristate
flabel metal2 s 21914 33544 21970 34344 0 FreeSans 224 90 0 0 wb_dat_i[0]
port 25 nsew signal input
flabel metal3 s 34168 23808 34968 23928 0 FreeSans 480 0 0 0 wb_dat_i[10]
port 26 nsew signal input
flabel metal2 s 6458 33544 6514 34344 0 FreeSans 224 90 0 0 wb_dat_i[11]
port 27 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 wb_dat_i[12]
port 28 nsew signal input
flabel metal3 s 34168 14288 34968 14408 0 FreeSans 480 0 0 0 wb_dat_i[13]
port 29 nsew signal input
flabel metal2 s 18694 33544 18750 34344 0 FreeSans 224 90 0 0 wb_dat_i[14]
port 30 nsew signal input
flabel metal3 s 34168 2728 34968 2848 0 FreeSans 480 0 0 0 wb_dat_i[15]
port 31 nsew signal input
flabel metal2 s 25134 33544 25190 34344 0 FreeSans 224 90 0 0 wb_dat_i[16]
port 32 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 wb_dat_i[17]
port 33 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 wb_dat_i[18]
port 34 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 wb_dat_i[19]
port 35 nsew signal input
flabel metal2 s 17406 33544 17462 34344 0 FreeSans 224 90 0 0 wb_dat_i[1]
port 36 nsew signal input
flabel metal3 s 34168 33328 34968 33448 0 FreeSans 480 0 0 0 wb_dat_i[20]
port 37 nsew signal input
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 wb_dat_i[21]
port 38 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 wb_dat_i[22]
port 39 nsew signal input
flabel metal3 s 34168 10888 34968 11008 0 FreeSans 480 0 0 0 wb_dat_i[23]
port 40 nsew signal input
flabel metal2 s 662 33544 718 34344 0 FreeSans 224 90 0 0 wb_dat_i[24]
port 41 nsew signal input
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 wb_dat_i[25]
port 42 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wb_dat_i[26]
port 43 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 wb_dat_i[27]
port 44 nsew signal input
flabel metal3 s 34168 30608 34968 30728 0 FreeSans 480 0 0 0 wb_dat_i[28]
port 45 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 wb_dat_i[29]
port 46 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wb_dat_i[2]
port 47 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wb_dat_i[30]
port 48 nsew signal input
flabel metal2 s 28998 0 29054 800 0 FreeSans 224 90 0 0 wb_dat_i[31]
port 49 nsew signal input
flabel metal3 s 34168 9528 34968 9648 0 FreeSans 480 0 0 0 wb_dat_i[3]
port 50 nsew signal input
flabel metal3 s 34168 4088 34968 4208 0 FreeSans 480 0 0 0 wb_dat_i[4]
port 51 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 wb_dat_i[5]
port 52 nsew signal input
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 wb_dat_i[6]
port 53 nsew signal input
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 wb_dat_i[7]
port 54 nsew signal input
flabel metal2 s 9678 33544 9734 34344 0 FreeSans 224 90 0 0 wb_dat_i[8]
port 55 nsew signal input
flabel metal3 s 34168 7488 34968 7608 0 FreeSans 480 0 0 0 wb_dat_i[9]
port 56 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 wb_dat_o[0]
port 57 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wb_dat_o[10]
port 58 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 wb_dat_o[11]
port 59 nsew signal tristate
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 wb_dat_o[12]
port 60 nsew signal tristate
flabel metal2 s 12898 33544 12954 34344 0 FreeSans 224 90 0 0 wb_dat_o[13]
port 61 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 wb_dat_o[14]
port 62 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 wb_dat_o[15]
port 63 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 wb_dat_o[16]
port 64 nsew signal tristate
flabel metal2 s 11610 33544 11666 34344 0 FreeSans 224 90 0 0 wb_dat_o[17]
port 65 nsew signal tristate
flabel metal2 s 20626 33544 20682 34344 0 FreeSans 224 90 0 0 wb_dat_o[18]
port 66 nsew signal tristate
flabel metal2 s 31574 33544 31630 34344 0 FreeSans 224 90 0 0 wb_dat_o[19]
port 67 nsew signal tristate
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 wb_dat_o[1]
port 68 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wb_dat_o[20]
port 69 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 wb_dat_o[21]
port 70 nsew signal tristate
flabel metal2 s 34150 33544 34206 34344 0 FreeSans 224 90 0 0 wb_dat_o[22]
port 71 nsew signal tristate
flabel metal2 s 26422 33544 26478 34344 0 FreeSans 224 90 0 0 wb_dat_o[23]
port 72 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wb_dat_o[24]
port 73 nsew signal tristate
flabel metal3 s 34168 31968 34968 32088 0 FreeSans 480 0 0 0 wb_dat_o[25]
port 74 nsew signal tristate
flabel metal3 s 34168 1368 34968 1488 0 FreeSans 480 0 0 0 wb_dat_o[26]
port 75 nsew signal tristate
flabel metal2 s 5170 33544 5226 34344 0 FreeSans 224 90 0 0 wb_dat_o[27]
port 76 nsew signal tristate
flabel metal3 s 34168 17008 34968 17128 0 FreeSans 480 0 0 0 wb_dat_o[28]
port 77 nsew signal tristate
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 wb_dat_o[29]
port 78 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 wb_dat_o[2]
port 79 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 wb_dat_o[30]
port 80 nsew signal tristate
flabel metal3 s 34168 19048 34968 19168 0 FreeSans 480 0 0 0 wb_dat_o[31]
port 81 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 wb_dat_o[3]
port 82 nsew signal tristate
flabel metal2 s 29642 33544 29698 34344 0 FreeSans 224 90 0 0 wb_dat_o[4]
port 83 nsew signal tristate
flabel metal2 s 28354 33544 28410 34344 0 FreeSans 224 90 0 0 wb_dat_o[5]
port 84 nsew signal tristate
flabel metal2 s 3882 33544 3938 34344 0 FreeSans 224 90 0 0 wb_dat_o[6]
port 85 nsew signal tristate
flabel metal2 s 8390 33544 8446 34344 0 FreeSans 224 90 0 0 wb_dat_o[7]
port 86 nsew signal tristate
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 wb_dat_o[8]
port 87 nsew signal tristate
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 wb_dat_o[9]
port 88 nsew signal tristate
flabel metal3 s 0 30608 800 30728 0 FreeSans 480 0 0 0 wb_stb_o
port 89 nsew signal tristate
flabel metal3 s 34168 15648 34968 15768 0 FreeSans 480 0 0 0 wb_we_o
port 90 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34968 34344
<< end >>
