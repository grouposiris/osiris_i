* NGSPICE file created from core.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt core clk i_instr_ID[0] i_instr_ID[10] i_instr_ID[11] i_instr_ID[12] i_instr_ID[13]
+ i_instr_ID[14] i_instr_ID[15] i_instr_ID[16] i_instr_ID[17] i_instr_ID[18] i_instr_ID[19]
+ i_instr_ID[1] i_instr_ID[20] i_instr_ID[21] i_instr_ID[22] i_instr_ID[23] i_instr_ID[24]
+ i_instr_ID[25] i_instr_ID[26] i_instr_ID[27] i_instr_ID[28] i_instr_ID[29] i_instr_ID[2]
+ i_instr_ID[30] i_instr_ID[31] i_instr_ID[3] i_instr_ID[4] i_instr_ID[5] i_instr_ID[6]
+ i_instr_ID[7] i_instr_ID[8] i_instr_ID[9] i_read_data_M[0] i_read_data_M[10] i_read_data_M[11]
+ i_read_data_M[12] i_read_data_M[13] i_read_data_M[14] i_read_data_M[15] i_read_data_M[16]
+ i_read_data_M[17] i_read_data_M[18] i_read_data_M[19] i_read_data_M[1] i_read_data_M[20]
+ i_read_data_M[21] i_read_data_M[22] i_read_data_M[23] i_read_data_M[24] i_read_data_M[25]
+ i_read_data_M[26] i_read_data_M[27] i_read_data_M[28] i_read_data_M[29] i_read_data_M[2]
+ i_read_data_M[30] i_read_data_M[31] i_read_data_M[3] i_read_data_M[4] i_read_data_M[5]
+ i_read_data_M[6] i_read_data_M[7] i_read_data_M[8] i_read_data_M[9] o_data_addr_M[0]
+ o_data_addr_M[10] o_data_addr_M[11] o_data_addr_M[12] o_data_addr_M[13] o_data_addr_M[14]
+ o_data_addr_M[15] o_data_addr_M[16] o_data_addr_M[17] o_data_addr_M[18] o_data_addr_M[19]
+ o_data_addr_M[1] o_data_addr_M[20] o_data_addr_M[21] o_data_addr_M[22] o_data_addr_M[23]
+ o_data_addr_M[24] o_data_addr_M[25] o_data_addr_M[26] o_data_addr_M[27] o_data_addr_M[28]
+ o_data_addr_M[29] o_data_addr_M[2] o_data_addr_M[30] o_data_addr_M[31] o_data_addr_M[3]
+ o_data_addr_M[4] o_data_addr_M[5] o_data_addr_M[6] o_data_addr_M[7] o_data_addr_M[8]
+ o_data_addr_M[9] o_mem_write_M o_pc_IF[0] o_pc_IF[10] o_pc_IF[11] o_pc_IF[12] o_pc_IF[13]
+ o_pc_IF[14] o_pc_IF[15] o_pc_IF[16] o_pc_IF[17] o_pc_IF[18] o_pc_IF[19] o_pc_IF[1]
+ o_pc_IF[20] o_pc_IF[21] o_pc_IF[22] o_pc_IF[23] o_pc_IF[24] o_pc_IF[25] o_pc_IF[26]
+ o_pc_IF[27] o_pc_IF[28] o_pc_IF[29] o_pc_IF[2] o_pc_IF[30] o_pc_IF[31] o_pc_IF[3]
+ o_pc_IF[4] o_pc_IF[5] o_pc_IF[6] o_pc_IF[7] o_pc_IF[8] o_pc_IF[9] o_write_data_M[0]
+ o_write_data_M[10] o_write_data_M[11] o_write_data_M[12] o_write_data_M[13] o_write_data_M[14]
+ o_write_data_M[15] o_write_data_M[16] o_write_data_M[17] o_write_data_M[18] o_write_data_M[19]
+ o_write_data_M[1] o_write_data_M[20] o_write_data_M[21] o_write_data_M[22] o_write_data_M[23]
+ o_write_data_M[24] o_write_data_M[25] o_write_data_M[26] o_write_data_M[27] o_write_data_M[28]
+ o_write_data_M[29] o_write_data_M[2] o_write_data_M[30] o_write_data_M[31] o_write_data_M[3]
+ o_write_data_M[4] o_write_data_M[5] o_write_data_M[6] o_write_data_M[7] o_write_data_M[8]
+ o_write_data_M[9] rst vccd1 vssd1
XANTENNA__4563__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7963_ _8091_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 _7963_/Q sky130_fd_sc_hd__dfxtp_1
X_6914_ _7010_/A _6914_/A2 _6943_/B _6913_/X vssd1 vssd1 vccd1 vccd1 _6914_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6090__B1 _6089_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7030__B _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3979__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5469__C _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7894_ _8504_/CLK _7894_/D vssd1 vssd1 vccd1 vccd1 _7894_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout162_A _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6845_ _6845_/A _6845_/B vssd1 vssd1 vccd1 vccd1 _6845_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_77_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5196__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6776_ _6776_/A _6776_/B vssd1 vssd1 vccd1 vccd1 _6776_/X sky130_fd_sc_hd__or2_4
X_3988_ _8072_/Q _3987_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _6787_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_45_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout427_A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5727_ _5738_/A _5730_/A _5727_/C vssd1 vssd1 vccd1 vccd1 _6380_/A sky130_fd_sc_hd__or3_2
X_8515_ _8515_/CLK _8515_/D vssd1 vssd1 vccd1 vccd1 _8515_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6932__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8446_ _8479_/CLK _8446_/D vssd1 vssd1 vccd1 vccd1 _8446_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5658_ _6494_/A _5658_/B vssd1 vssd1 vccd1 vccd1 _5658_/X sky130_fd_sc_hd__and2_1
XFILLER_0_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4609_ _4608_/X _4607_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4609_/X sky130_fd_sc_hd__mux2_1
X_5589_ _6849_/A _5584_/B _5617_/B1 hold999/X vssd1 vssd1 vccd1 vccd1 _5589_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_103_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5705__S _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6696__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8377_ _8378_/CLK _8377_/D _7271_/Y vssd1 vssd1 vccd1 vccd1 _8377_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold362 _7386_/Q vssd1 vssd1 vccd1 vccd1 _5453_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 _7339_/Q vssd1 vssd1 vccd1 vccd1 _5436_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold351 _5438_/X vssd1 vssd1 vccd1 vccd1 _7627_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7328_ _8019_/CLK _7328_/D vssd1 vssd1 vccd1 vccd1 _7328_/Q sky130_fd_sc_hd__dfxtp_1
X_7259_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7259_/Y sky130_fd_sc_hd__inv_2
Xhold373 _5289_/X vssd1 vssd1 vccd1 vccd1 _7493_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _7342_/Q vssd1 vssd1 vccd1 vccd1 _5439_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _5248_/X vssd1 vssd1 vccd1 vccd1 _7456_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5120__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1040 _5345_/X vssd1 vssd1 vccd1 vccd1 _7572_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 _8152_/Q vssd1 vssd1 vccd1 vccd1 _6580_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 _5266_/X vssd1 vssd1 vccd1 vccd1 _7470_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3682__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1073 _7794_/Q vssd1 vssd1 vccd1 vccd1 _5610_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 _5194_/X vssd1 vssd1 vccd1 vccd1 _7408_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _8138_/Q vssd1 vssd1 vccd1 vccd1 _6566_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5676__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5395__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6687__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3952__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4793__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5647__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4755__A _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4960_ _4958_/X _4959_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__mux2_1
X_3911_ _3923_/B _7941_/Q vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_80_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4891_ _8182_/Q _8214_/Q _8278_/Q _7786_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4891_/X sky130_fd_sc_hd__mux4_1
X_6630_ _7029_/A _6630_/A2 _6605_/B _6629_/X vssd1 vssd1 vccd1 vccd1 _6630_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_80_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3842_ _4775_/B _4071_/A2 _4071_/B1 _6971_/A _3841_/X vssd1 vssd1 vccd1 vccd1 _6126_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_58_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5178__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6914__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6561_ _6777_/A _6592_/A2 _6592_/B1 hold647/X vssd1 vssd1 vccd1 vccd1 _6561_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8300_ _8426_/CLK _8300_/D vssd1 vssd1 vccd1 vccd1 _8300_/Q sky130_fd_sc_hd__dfxtp_1
X_5512_ _8231_/Q _5542_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7701_/D sky130_fd_sc_hd__and3_1
X_3773_ _3770_/X _3771_/Y _3772_/X _4014_/A vssd1 vssd1 vccd1 vccd1 _3773_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6492_ _6494_/A hold45/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__and2_1
XFILLER_0_54_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8231_ _8231_/CLK _8231_/D vssd1 vssd1 vccd1 vccd1 _8231_/Q sky130_fd_sc_hd__dfxtp_1
X_5443_ _5443_/A _7030_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _5443_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6678__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5350__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5374_ _5374_/A _6974_/A _5408_/C vssd1 vssd1 vccd1 vccd1 _6981_/A sky130_fd_sc_hd__or3_1
XANTENNA__3834__A _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8162_ _8427_/CLK _8162_/D vssd1 vssd1 vccd1 vccd1 _8162_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4784__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5981__S0 _5716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7113_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7113_/Y sky130_fd_sc_hd__inv_2
X_4325_ _4325_/A _4325_/B vssd1 vssd1 vccd1 vccd1 _4325_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5638__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8093_ _8385_/CLK _8127_/D vssd1 vssd1 vccd1 vccd1 _8093_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5102__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7044_ _7044_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7044_/Y sky130_fd_sc_hd__nand2_1
X_4256_ _8502_/Q _4257_/B vssd1 vssd1 vccd1 vccd1 _4256_/Y sky130_fd_sc_hd__nor2_1
X_4187_ _8512_/Q _4187_/B vssd1 vssd1 vccd1 vccd1 _4187_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout377_A _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7946_ _8500_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _7946_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7877_ _8080_/CLK _7877_/D vssd1 vssd1 vccd1 vccd1 _7877_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6828_ _7029_/A _6828_/A2 _6779_/B _6827_/X vssd1 vssd1 vccd1 vccd1 _6828_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6759_ _6941_/A _6773_/A2 _6773_/B1 hold509/X vssd1 vssd1 vccd1 vccd1 _6759_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_93_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3975__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8429_ _8465_/CLK _8429_/D vssd1 vssd1 vccd1 vccd1 _8429_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5943__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold170 _7852_/Q vssd1 vssd1 vccd1 vccd1 _6473_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5341__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold181 _6470_/X vssd1 vssd1 vccd1 vccd1 _7952_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _7842_/Q vssd1 vssd1 vccd1 vccd1 _6463_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5629__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_31_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4527__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6357__A1 _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6109__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6109__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6949__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_104_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5332__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6965__A _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1809 _7351_/Q vssd1 vssd1 vccd1 vccd1 hold1809/X sky130_fd_sc_hd__dlygate4sd3_1
X_4110_ _6035_/A _6032_/A vssd1 vssd1 vccd1 vccd1 _4110_/Y sky130_fd_sc_hd__nand2b_1
X_5090_ input6/X _5099_/B _5002_/X _5089_/X vssd1 vssd1 vccd1 vccd1 _7357_/D sky130_fd_sc_hd__o211a_1
X_4041_ _5990_/A vssd1 vssd1 vccd1 vccd1 _4041_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6045__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5992_ _5993_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5992_/Y sky130_fd_sc_hd__nand2_1
X_7800_ _8450_/CLK _7800_/D vssd1 vssd1 vccd1 vccd1 _7800_/Q sky130_fd_sc_hd__dfxtp_1
X_7731_ _8487_/CLK _7731_/D vssd1 vssd1 vccd1 vccd1 _7731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4943_ _4942_/X _4939_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8253_/D sky130_fd_sc_hd__mux2_1
X_7662_ _8079_/CLK _7662_/D vssd1 vssd1 vccd1 vccd1 _7662_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4071__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3998__A_N _7283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6613_ _6853_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6613_/X sky130_fd_sc_hd__and2_1
X_4874_ _8340_/Q _7816_/Q _7482_/Q _7450_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4874_/X sky130_fd_sc_hd__mux4_1
X_3825_ _8000_/Q _4068_/A2 _4068_/B1 _8032_/Q _3824_/X vssd1 vssd1 vccd1 vccd1 _3825_/X
+ sky130_fd_sc_hd__a221o_1
X_7593_ _8427_/CLK _7593_/D vssd1 vssd1 vccd1 vccd1 _7593_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6859__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_12_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_12_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_3756_ _3756_/A1 _4073_/A2 _6941_/A _4073_/B2 _3755_/X vssd1 vssd1 vccd1 vccd1 _3757_/B
+ sky130_fd_sc_hd__a221o_2
X_6544_ _7018_/A _6544_/B vssd1 vssd1 vccd1 vccd1 _8026_/D sky130_fd_sc_hd__and2_1
X_6475_ _6524_/A _6475_/B vssd1 vssd1 vccd1 vccd1 _6475_/X sky130_fd_sc_hd__and2_1
X_3687_ _7834_/Q _7660_/Q vssd1 vssd1 vccd1 vccd1 _3687_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__5482__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8214_ _8402_/CLK _8214_/D vssd1 vssd1 vccd1 vccd1 _8214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7036__A _7076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5426_ _5426_/A _5503_/B _5462_/C vssd1 vssd1 vccd1 vccd1 _5426_/X sky130_fd_sc_hd__and3_1
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4379__B _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5323__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8145_ _8338_/CLK _8145_/D vssd1 vssd1 vccd1 vccd1 _8145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3885__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6875__A _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5357_ _6949_/A _5367_/A2 _5367_/B1 hold749/X vssd1 vssd1 vccd1 vccd1 _5357_/X sky130_fd_sc_hd__a22o_1
X_8076_ _8519_/CLK _8110_/D vssd1 vssd1 vccd1 vccd1 _8076_/Q sky130_fd_sc_hd__dfxtp_1
X_5288_ _6891_/A _5294_/A2 _5294_/B1 hold679/X vssd1 vssd1 vccd1 vccd1 _5288_/X sky130_fd_sc_hd__a22o_1
X_4308_ _4308_/A _4308_/B vssd1 vssd1 vccd1 vccd1 _4308_/Y sky130_fd_sc_hd__nand2_1
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4239_/X sky130_fd_sc_hd__xor2_1
XANTENNA__6284__A0 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7027_ _7027_/A _7027_/B vssd1 vssd1 vccd1 vccd1 _7027_/X sky130_fd_sc_hd__and2_1
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6587__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7929_ _8010_/CLK _7929_/D vssd1 vssd1 vccd1 vccd1 _7929_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6115__A _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4996__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5314__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6785__A _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4920__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6578__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3649__A _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4684__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5250__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4590_ _8336_/Q _7812_/Q _7478_/Q _7446_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4590_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6750__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4987__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold928 _5245_/X vssd1 vssd1 vccd1 vccd1 _7453_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold917 _7435_/Q vssd1 vssd1 vccd1 vccd1 hold917/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold906 _6686_/X vssd1 vssd1 vccd1 vccd1 _8213_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6260_ _6262_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6263_/A sky130_fd_sc_hd__and2_1
Xhold939 _8318_/Q vssd1 vssd1 vccd1 vccd1 hold939/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5305__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5856__A3 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5211_ _6951_/A _5221_/A2 _5221_/B1 hold639/X vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__a22o_1
X_6191_ _6191_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6192_/B sky130_fd_sc_hd__nor2_1
X_5142_ _5142_/A1 _5144_/A2 _5146_/B1 _5141_/X vssd1 vssd1 vccd1 vccd1 _7383_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3867__A2 _6441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1606 _5392_/B vssd1 vssd1 vccd1 vccd1 _5408_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__5069__A1 _5408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1617 _3981_/X vssd1 vssd1 vccd1 vccd1 _6428_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1628 _4203_/Y vssd1 vssd1 vccd1 vccd1 _4205_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5073_ _5073_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5073_/Y sky130_fd_sc_hd__nand2_1
Xhold1639 _8513_/Q vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__buf_1
X_4024_ _8078_/Q _4023_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4024_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6569__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5975_ _5975_/A _5975_/B vssd1 vssd1 vccd1 vccd1 _5976_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4675__S0 _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4926_ _8187_/Q _8219_/Q _8283_/Q _7791_/Q _4996_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4926_/X sky130_fd_sc_hd__mux4_1
X_7714_ _8469_/CLK _7714_/D vssd1 vssd1 vccd1 vccd1 _7714_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3993__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4857_ _8467_/Q _8399_/Q _8431_/Q _8305_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4857_/X sky130_fd_sc_hd__mux4_1
X_7645_ _8504_/CLK _7645_/D vssd1 vssd1 vccd1 vccd1 _7645_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7576_ _8143_/CLK _7576_/D vssd1 vssd1 vccd1 vccd1 _7576_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3808_ _3808_/A0 _3807_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6386_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_132_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4788_ _4787_/X _4786_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5493__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6527_ _7019_/A _6527_/B vssd1 vssd1 vccd1 vccd1 _8009_/D sky130_fd_sc_hd__and2_1
XFILLER_0_113_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3739_ _7998_/Q _4068_/A2 _4068_/B1 _8030_/Q _3738_/X vssd1 vssd1 vccd1 vccd1 _3739_/X
+ sky130_fd_sc_hd__a221o_1
X_6458_ _7837_/Q _7940_/Q _6911_/A vssd1 vssd1 vccd1 vccd1 _6458_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5409_ _5409_/A _6554_/C vssd1 vssd1 vccd1 vccd1 _6973_/C sky130_fd_sc_hd__nand2_1
X_6389_ _6387_/X _6389_/B vssd1 vssd1 vccd1 vccd1 _6390_/B sky130_fd_sc_hd__and2b_1
XANTENNA__5713__S _5716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8128_ _8128_/CLK _8128_/D vssd1 vssd1 vccd1 vccd1 _8128_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6257__B1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3741__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8059_ _8059_/CLK _8059_/D vssd1 vssd1 vccd1 vccd1 _8059_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4902__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6024__A3 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5232__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4999__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5684__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3916__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6732__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4969__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6248__A0 _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4763__A _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4026__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4657__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5760_ _6270_/A _5759_/A _5748_/Y vssd1 vssd1 vccd1 vccd1 _5760_/Y sky130_fd_sc_hd__a21oi_1
X_7214__92 _8385_/CLK vssd1 vssd1 vccd1 vccd1 _8127_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5691_ _5723_/B _5727_/C vssd1 vssd1 vccd1 vccd1 _6008_/B sky130_fd_sc_hd__nor2_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4711_ _4709_/X _4710_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4642_ _8183_/Q _8215_/Q _8279_/Q _7787_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4642_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_72_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7430_ _8486_/CLK _7430_/D vssd1 vssd1 vccd1 vccd1 _7430_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6723__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7361_ _8361_/CLK _7361_/D vssd1 vssd1 vccd1 vccd1 _7361_/Q sky130_fd_sc_hd__dfxtp_1
X_4573_ _8463_/Q _8395_/Q _8427_/Q _8301_/Q _4727_/S0 _7050_/A vssd1 vssd1 vccd1 vccd1
+ _4573_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold703 _8277_/Q vssd1 vssd1 vccd1 vccd1 hold703/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7292_ _8510_/CLK _7292_/D _7102_/Y vssd1 vssd1 vccd1 vccd1 _7292_/Q sky130_fd_sc_hd__dfrtp_4
X_6312_ _6391_/A _6301_/X _6306_/X _6311_/Y vssd1 vssd1 vccd1 vccd1 _6312_/X sky130_fd_sc_hd__o211a_1
Xhold736 _5220_/X vssd1 vssd1 vccd1 vccd1 _7434_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _5325_/X vssd1 vssd1 vccd1 vccd1 _7556_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold725 _7536_/Q vssd1 vssd1 vccd1 vccd1 hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 _6676_/X vssd1 vssd1 vccd1 vccd1 _8203_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 _7496_/Q vssd1 vssd1 vccd1 vccd1 hold747/X sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ _6244_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _6246_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold769 _7593_/Q vssd1 vssd1 vccd1 vccd1 hold769/X sky130_fd_sc_hd__dlygate4sd3_1
X_6174_ _6175_/A _6175_/B vssd1 vssd1 vccd1 vccd1 _6174_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout192_A _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5125_ _5442_/A _5442_/C vssd1 vssd1 vccd1 vccd1 _5125_/X sky130_fd_sc_hd__or2_1
Xhold1425 _4336_/Y vssd1 vssd1 vccd1 vccd1 _4337_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1403 _8385_/Q vssd1 vssd1 vccd1 vccd1 _5058_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1414 hold1803/X vssd1 vssd1 vccd1 vccd1 _5040_/A1 sky130_fd_sc_hd__buf_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1447 _7638_/Q vssd1 vssd1 vccd1 vccd1 _4209_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _4379_/A _5069_/S _5182_/B1 _5055_/X vssd1 vssd1 vccd1 vccd1 _7340_/D sky130_fd_sc_hd__o211a_1
Xhold1436 _4257_/Y vssd1 vssd1 vccd1 vccd1 _4258_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1458 _4246_/X vssd1 vssd1 vccd1 vccd1 _5564_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4896__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1469 _7292_/Q vssd1 vssd1 vccd1 vccd1 _5140_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4007_ _6016_/A _6013_/A vssd1 vssd1 vccd1 vccd1 _4008_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3988__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout457_A _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5214__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5958_ _5881_/C _5957_/Y _5954_/Y vssd1 vssd1 vccd1 vccd1 _5958_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6962__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4909_ _8345_/Q _7821_/Q _7487_/Q _7455_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4909_/X sky130_fd_sc_hd__mux4_1
XANTENNA_hold1474_A _7294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5889_ _5889_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _5892_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5708__S _5716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7628_ _8030_/CLK _7628_/D vssd1 vssd1 vccd1 vccd1 _7628_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6714__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6112__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3736__B _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1641_A _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7559_ _8442_/CLK _7559_/D vssd1 vssd1 vccd1 vccd1 _7559_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__8030__D _8030_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5150__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4639__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5205__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3767__A1 _3766_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4522__S _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4811__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_5 _4059_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output86_A _8103_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6957__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4758__A _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6973__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4878__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6930_ _7008_/A _6930_/A2 _6943_/B _6929_/X vssd1 vssd1 vccd1 vccd1 _6930_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_16_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6861_ _6927_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6861_/X sky130_fd_sc_hd__and2_1
XFILLER_0_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5101__B _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5812_ _5955_/A _5804_/A _5926_/B vssd1 vssd1 vccd1 vccd1 _5812_/X sky130_fd_sc_hd__o21a_1
X_6792_ _7026_/A _6792_/A2 _6838_/A3 _6791_/X vssd1 vssd1 vccd1 vccd1 _6792_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_123_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6944__B2 _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6944__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8531_ _8531_/A _7094_/X vssd1 vssd1 vccd1 vccd1 _8531_/Z sky130_fd_sc_hd__ebufn_1
X_5743_ _3935_/A _6011_/A2 _5743_/B1 _6741_/A vssd1 vssd1 vccd1 vccd1 _5743_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8462_ _8462_/CLK _8462_/D vssd1 vssd1 vccd1 vccd1 _8462_/Q sky130_fd_sc_hd__dfxtp_1
X_5674_ _6551_/A _5674_/B vssd1 vssd1 vccd1 vccd1 _5674_/X sky130_fd_sc_hd__and2_1
X_7413_ _8175_/CLK _7413_/D vssd1 vssd1 vccd1 vccd1 _7413_/Q sky130_fd_sc_hd__dfxtp_1
X_8393_ _8425_/CLK _8393_/D vssd1 vssd1 vccd1 vccd1 _8393_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4625_ _8341_/Q _7817_/Q _7483_/Q _7451_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4625_/X sky130_fd_sc_hd__mux4_1
X_7344_ _8011_/CLK _7344_/D vssd1 vssd1 vccd1 vccd1 _7344_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4556_ _8138_/Q _7537_/Q _7409_/Q _7569_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4556_/X sky130_fd_sc_hd__mux4_1
Xhold511 _7547_/Q vssd1 vssd1 vccd1 vccd1 hold511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 _5458_/X vssd1 vssd1 vccd1 vccd1 _7647_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6867__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold533 _7812_/Q vssd1 vssd1 vccd1 vccd1 hold533/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold544 _5190_/X vssd1 vssd1 vccd1 vccd1 _7404_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold522 _5284_/X vssd1 vssd1 vccd1 vccd1 _7488_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _5636_/X vssd1 vssd1 vccd1 vccd1 _7816_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6359__S _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold588 _6690_/X vssd1 vssd1 vccd1 vccd1 _8217_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7044__A _7044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4487_ _5178_/A1 _4487_/A1 _5468_/C vssd1 vssd1 vccd1 vccd1 _7311_/D sky130_fd_sc_hd__mux2_1
Xhold555 _8288_/Q vssd1 vssd1 vccd1 vccd1 hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _7486_/Q vssd1 vssd1 vccd1 vccd1 hold577/X sky130_fd_sc_hd__dlygate4sd3_1
X_7275_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7275_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5132__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5490__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6226_ _6226_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6227_/B sky130_fd_sc_hd__nor2_1
Xhold599 _8317_/Q vssd1 vssd1 vccd1 vccd1 hold599/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1200 _6868_/X vssd1 vssd1 vccd1 vccd1 _8400_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6157_ _6157_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6159_/A sky130_fd_sc_hd__xor2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6883__A _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1222 _6864_/X vssd1 vssd1 vccd1 vccd1 _8398_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 _8175_/Q vssd1 vssd1 vccd1 vccd1 _6622_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 _8451_/Q vssd1 vssd1 vccd1 vccd1 _6972_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ input15/X _5099_/B _5002_/X _5107_/X vssd1 vssd1 vccd1 vccd1 _7366_/D sky130_fd_sc_hd__o211a_1
Xhold1255 _8347_/Q vssd1 vssd1 vccd1 vccd1 _6820_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ _6270_/A _5901_/X _5957_/B vssd1 vssd1 vccd1 vccd1 _6088_/X sky130_fd_sc_hd__o21a_1
Xhold1244 _6634_/X vssd1 vssd1 vccd1 vccd1 _8181_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _6896_/X vssd1 vssd1 vccd1 vccd1 _8414_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 _6610_/X vssd1 vssd1 vccd1 vccd1 _8169_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1288 _8364_/Q vssd1 vssd1 vccd1 vccd1 _4434_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1277 _6852_/X vssd1 vssd1 vccd1 vccd1 _8392_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5039_ _5429_/A _5465_/C vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5199__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5011__B _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6396__C1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3747__A _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6148__C1 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_114_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8476_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6699__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6777__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput64 _8101_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[0] sky130_fd_sc_hd__buf_12
Xoutput75 _8102_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[1] sky130_fd_sc_hd__buf_12
XANTENNA__6793__A _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput86 _8103_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[2] sky130_fd_sc_hd__buf_12
XFILLER_0_37_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput97 _7292_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[10] sky130_fd_sc_hd__buf_12
XANTENNA_output124_A _7289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3988__A1 _3987_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6926__A1 _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3657__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6033__A _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_105_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8160_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4165__A1 _8516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5362__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4410_ _4410_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4410_/Y sky130_fd_sc_hd__nor2_1
X_5390_ _5389_/A _5374_/A _5388_/X vssd1 vssd1 vccd1 vccd1 _7055_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_22_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3912__B2 _8005_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6179__S _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4341_ _4383_/A _4383_/B _4341_/C vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_1_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5114__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout309 _5297_/Y vssd1 vssd1 vccd1 vccd1 _5299_/B sky130_fd_sc_hd__buf_8
X_7060_ _7071_/B _7059_/Y _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8502_/D sky130_fd_sc_hd__a21oi_1
X_4272_ _4270_/Y _4272_/B vssd1 vssd1 vccd1 vccd1 _4272_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_10_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6011_ _6011_/A1 _6011_/A2 _6005_/Y _6010_/X _6911_/A vssd1 vssd1 vccd1 vccd1 _7877_/D
+ sky130_fd_sc_hd__a221oi_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5968__A2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6208__A _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7962_ _8379_/CLK hold74/X vssd1 vssd1 vccd1 vccd1 _7962_/Q sky130_fd_sc_hd__dfxtp_1
X_6913_ _6913_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6913_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6090__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7030__C _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3979__A1 _4751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3979__B2 _3977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7893_ _8419_/CLK _7893_/D vssd1 vssd1 vccd1 vccd1 _7893_/Q sky130_fd_sc_hd__dfxtp_1
X_6844_ _6777_/A _6845_/B _6843_/X vssd1 vssd1 vccd1 vccd1 _6844_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6775_ _6776_/A _6776_/B vssd1 vssd1 vccd1 vccd1 _6775_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_107_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3987_ _7976_/Q _4079_/A2 _4079_/B1 _8008_/Q _3986_/X vssd1 vssd1 vccd1 vccd1 _3987_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5485__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4162__S _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8514_ _8515_/CLK _8514_/D vssd1 vssd1 vccd1 vccd1 _8514_/Q sky130_fd_sc_hd__dfxtp_1
X_5726_ _5727_/C _5732_/D vssd1 vssd1 vccd1 vccd1 _5726_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_45_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8445_ _8445_/CLK _8445_/D vssd1 vssd1 vccd1 vccd1 _8445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5657_ _5667_/A _5657_/B vssd1 vssd1 vccd1 vccd1 _5657_/X sky130_fd_sc_hd__and2_1
X_5588_ _6847_/A _5585_/B _5585_/Y hold260/X vssd1 vssd1 vccd1 vccd1 _5588_/X sky130_fd_sc_hd__o22a_1
X_4608_ _8468_/Q _8400_/Q _8432_/Q _8306_/Q _4611_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4608_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_115_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5353__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8376_ _8378_/CLK _8376_/D _7270_/Y vssd1 vssd1 vccd1 vccd1 _8376_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4539_ _4538_/X _4537_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _4539_/X sky130_fd_sc_hd__mux2_1
Xhold352 _7468_/Q vssd1 vssd1 vccd1 vccd1 hold352/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _7317_/Q vssd1 vssd1 vccd1 vccd1 _5414_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold341 _5436_/X vssd1 vssd1 vccd1 vccd1 _7625_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7327_ _8019_/CLK _7327_/D vssd1 vssd1 vccd1 vccd1 _7327_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold363 _5453_/X vssd1 vssd1 vccd1 vccd1 _7642_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7258_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7258_/Y sky130_fd_sc_hd__inv_2
Xhold396 _7827_/Q vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _5439_/X vssd1 vssd1 vccd1 vccd1 _7628_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _7388_/Q vssd1 vssd1 vccd1 vccd1 _5455_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6209_ _6209_/A _6209_/B vssd1 vssd1 vccd1 vccd1 _6210_/B sky130_fd_sc_hd__or2_1
Xhold1030 _5310_/X vssd1 vssd1 vccd1 vccd1 _7541_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 _7412_/Q vssd1 vssd1 vccd1 vccd1 _5198_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5959__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1052 _6580_/X vssd1 vssd1 vccd1 vccd1 _8152_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 _5610_/X vssd1 vssd1 vccd1 vccd1 _7794_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 _8137_/Q vssd1 vssd1 vccd1 vccd1 _6565_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1085 _7552_/Q vssd1 vssd1 vccd1 vccd1 _5321_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6620__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1096 _6566_/X vssd1 vssd1 vccd1 vccd1 _8138_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5592__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_5_clk_A clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5344__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5647__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4247__S _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5867__A _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3910_ _3910_/A _3910_/B vssd1 vssd1 vccd1 vccd1 _4097_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4890_ _4888_/X _4889_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4771__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3841_ _7731_/Q _3841_/B vssd1 vssd1 vccd1 vccd1 _3841_/X sky130_fd_sc_hd__or2_1
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6560_ _6706_/A _6560_/B vssd1 vssd1 vccd1 vccd1 _6560_/Y sky130_fd_sc_hd__nand2_1
X_3772_ _4083_/B _3939_/B hold1520/X vssd1 vssd1 vccd1 vccd1 _3772_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_104_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5511_ _8230_/Q _7073_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7700_/D sky130_fd_sc_hd__and3_1
XFILLER_0_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6491_ _6498_/A _6491_/B vssd1 vssd1 vccd1 vccd1 _6491_/X sky130_fd_sc_hd__and2_1
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8230_ _8230_/CLK _8230_/D vssd1 vssd1 vccd1 vccd1 _8230_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5442_ _5442_/A _7082_/A _5442_/C vssd1 vssd1 vccd1 vccd1 _5442_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3777__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5373_ _5374_/A _5408_/C vssd1 vssd1 vccd1 vccd1 _5373_/Y sky130_fd_sc_hd__nor2_1
X_8161_ _8419_/CLK _8161_/D vssd1 vssd1 vccd1 vccd1 _8161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5981__S1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8092_ _8419_/CLK _8126_/D vssd1 vssd1 vccd1 vccd1 _8092_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5107__A _7044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7112_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7112_/Y sky130_fd_sc_hd__inv_2
X_4324_ _4322_/Y _4324_/B vssd1 vssd1 vccd1 vccd1 _4324_/X sky130_fd_sc_hd__and2b_1
X_7043_ _7031_/Y _7043_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _7043_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5638__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4255_ _4416_/A _4413_/B vssd1 vssd1 vccd1 vccd1 _4255_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6850__A3 _6842_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4186_ _8512_/Q _4187_/B vssd1 vssd1 vccd1 vccd1 _4186_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout272_A _3841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7945_ _7977_/CLK _7945_/D vssd1 vssd1 vccd1 vccd1 _7945_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7876_ _8517_/CLK _7876_/D vssd1 vssd1 vccd1 vccd1 _7876_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5496__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6827_ _6959_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6827_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7175__53 _8010_/CLK vssd1 vssd1 vccd1 vccd1 _8055_/CLK sky130_fd_sc_hd__inv_2
X_6758_ _6939_/A _6773_/A2 _6773_/B1 hold675/X vssd1 vssd1 vccd1 vccd1 _6758_/X sky130_fd_sc_hd__a22o_1
X_5709_ _6244_/A _6262_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5709_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5716__S _5716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6689_ _6945_/A _6701_/A2 _6701_/B1 hold839/X vssd1 vssd1 vccd1 vccd1 _6689_/X sky130_fd_sc_hd__a22o_1
XANTENNA_hold1554_A _4052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8428_ _8428_/CLK _8428_/D vssd1 vssd1 vccd1 vccd1 _8428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4620__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5326__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8359_ _8361_/CLK _8359_/D _7253_/Y vssd1 vssd1 vccd1 vccd1 _8359_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3888__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold160 _7866_/Q vssd1 vssd1 vccd1 vccd1 _6487_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _6473_/X vssd1 vssd1 vccd1 vccd1 _7955_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 _7738_/Q vssd1 vssd1 vccd1 vccd1 _6489_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _6463_/X vssd1 vssd1 vccd1 vccd1 _7945_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5629__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7234__112 _8154_/CLK vssd1 vssd1 vccd1 vccd1 _8244_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5687__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__A2 _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5317__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3879__B1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6965__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6457__S _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4766__A _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4040_ _4040_/A0 _4039_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _5990_/A sky130_fd_sc_hd__mux2_2
XANTENNA__6293__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5096__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6832__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4056__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5991_ _5993_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5994_/A sky130_fd_sc_hd__and2_1
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7730_ _8354_/CLK _7730_/D vssd1 vssd1 vccd1 vccd1 _7730_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4942_ _4941_/X _4940_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__mux2_1
X_7661_ _8080_/CLK _7661_/D vssd1 vssd1 vccd1 vccd1 _7661_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4873_ _4872_/X _4869_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8243_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6612_ _7024_/A _6612_/A2 _6666_/A3 _6611_/X vssd1 vssd1 vccd1 vccd1 _6612_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_131_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5020__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4006__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7592_ _8354_/CLK _7592_/D vssd1 vssd1 vccd1 vccd1 _7592_/Q sky130_fd_sc_hd__dfxtp_1
X_3824_ _4067_/A_N _7968_/Q vssd1 vssd1 vccd1 vccd1 _3824_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3755_ _4760_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3755_/X sky130_fd_sc_hd__and2_1
XFILLER_0_55_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6543_ _6545_/A _6543_/B vssd1 vssd1 vccd1 vccd1 _8025_/D sky130_fd_sc_hd__and2_1
XANTENNA__5763__C _5971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3686_ _4769_/B _4071_/A2 _4071_/B1 _6959_/A _3685_/X vssd1 vssd1 vccd1 vccd1 _6298_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5308__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6474_ _6550_/A hold15/X vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__and2_1
XANTENNA__7036__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8213_ _8431_/CLK _8213_/D vssd1 vssd1 vccd1 vccd1 _8213_/Q sky130_fd_sc_hd__dfxtp_1
X_5425_ _5425_/A _5503_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _5425_/X sky130_fd_sc_hd__and3_1
XFILLER_0_112_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5356_ _6947_/A _5367_/A2 _5367_/B1 hold699/X vssd1 vssd1 vccd1 vccd1 _5356_/X sky130_fd_sc_hd__a22o_1
X_8144_ _8448_/CLK _8144_/D vssd1 vssd1 vccd1 vccd1 _8144_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6875__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8075_ _8510_/CLK _8109_/D vssd1 vssd1 vccd1 vccd1 _8075_/Q sky130_fd_sc_hd__dfxtp_1
X_5287_ _6955_/A _5294_/A2 _5294_/B1 hold815/X vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__a22o_1
X_4307_ _4307_/A _7652_/Q vssd1 vssd1 vccd1 vccd1 _4307_/Y sky130_fd_sc_hd__nand2_1
X_4238_ _4228_/Y _4231_/X _4230_/B vssd1 vssd1 vccd1 vccd1 _4238_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6284__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7052__A _7052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7026_ _7026_/A _7026_/B vssd1 vssd1 vccd1 vccd1 _7026_/X sky130_fd_sc_hd__and2_1
XFILLER_0_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4169_ _4169_/A _4169_/B vssd1 vssd1 vccd1 vccd1 _4169_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_94_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _8480_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6891__A _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4047__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6587__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5795__A0 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7928_ _8008_/CLK _7928_/D vssd1 vssd1 vccd1 vccd1 _7928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5300__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7859_ _8090_/CLK _7859_/D vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7872__D _7872_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6785__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5078__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6275__B2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6814__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_85_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _8008_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6578__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4525__S _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4684__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5250__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6750__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold907 _7546_/Q vssd1 vssd1 vccd1 vccd1 hold907/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 _5221_/X vssd1 vssd1 vccd1 vccd1 _7435_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold929 _7777_/Q vssd1 vssd1 vccd1 vccd1 hold929/X sky130_fd_sc_hd__dlygate4sd3_1
X_5210_ _6949_/A _5188_/B _5220_/B1 hold673/X vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6190_ _6191_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6190_/Y sky130_fd_sc_hd__nand2_1
X_5141_ _5450_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _5141_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5072_ input27/X _4448_/B _5140_/B1 _5071_/X vssd1 vssd1 vccd1 vccd1 _7348_/D sky130_fd_sc_hd__o211a_1
Xhold1607 _8503_/Q vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__buf_1
X_4023_ _7982_/Q _4079_/A2 _4079_/B1 _8014_/Q _4022_/X vssd1 vssd1 vccd1 vccd1 _4023_/X
+ sky130_fd_sc_hd__a221o_2
Xhold1629 _4205_/X vssd1 vssd1 vccd1 vccd1 _5558_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1618 _7654_/Q vssd1 vssd1 vccd1 vccd1 _4323_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_76_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _8500_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_92_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6569__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5777__A0 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5241__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5974_ _5974_/A _5974_/B vssd1 vssd1 vccd1 vccd1 _5975_/B sky130_fd_sc_hd__or2_1
X_7713_ _8328_/CLK _7713_/D vssd1 vssd1 vccd1 vccd1 _7713_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4675__S1 _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4925_ _4923_/X _4924_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4856_ _8177_/Q _8209_/Q _8273_/Q _7781_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4856_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7644_ _8195_/CLK _7644_/D vssd1 vssd1 vccd1 vccd1 _7644_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout235_A _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3807_ _3807_/A1 _4073_/A2 _3803_/X _4073_/B2 _3806_/X vssd1 vssd1 vccd1 vccd1 _3807_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_51_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7575_ _8475_/CLK _7575_/D vssd1 vssd1 vccd1 vccd1 _7575_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4787_ _8457_/Q _8389_/Q _8421_/Q _8295_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4787_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_105_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5493__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4170__S _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7145__23 _8478_/CLK vssd1 vssd1 vccd1 vccd1 _7522_/CLK sky130_fd_sc_hd__inv_2
XANTENNA_fanout402_A hold1746/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6526_ _6551_/A _6526_/B vssd1 vssd1 vccd1 vccd1 _8008_/D sky130_fd_sc_hd__and2_1
X_3738_ _4067_/A_N _7966_/Q vssd1 vssd1 vccd1 vccd1 _3738_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_42_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6457_ _6457_/A0 _7939_/Q _6911_/A vssd1 vssd1 vccd1 vccd1 _6457_/X sky130_fd_sc_hd__mux2_1
X_3669_ _3669_/A _3669_/B vssd1 vssd1 vccd1 vccd1 _3669_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5408_ _6553_/A _5408_/B _5408_/C vssd1 vssd1 vccd1 vccd1 _6554_/C sky130_fd_sc_hd__or3_1
X_6388_ _6388_/A _6388_/B vssd1 vssd1 vccd1 vccd1 _6389_/B sky130_fd_sc_hd__or2_1
XFILLER_0_2_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5339_ _6847_/A _5336_/B _5336_/Y hold258/X vssd1 vssd1 vccd1 vccd1 _5339_/X sky130_fd_sc_hd__o22a_1
X_8127_ _8127_/CLK _8127_/D vssd1 vssd1 vccd1 vccd1 _8127_/Q sky130_fd_sc_hd__dfxtp_1
X_8058_ _8058_/CLK _8058_/D vssd1 vssd1 vccd1 vccd1 _8058_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__8028__D _8028_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _8362_/CLK sky130_fd_sc_hd__clkbuf_16
X_7009_ _7023_/A _7009_/B vssd1 vssd1 vccd1 vccd1 _7009_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_103_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6126__A _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5232__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4080__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6732__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6248__A1 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_58_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _8028_/CLK sky130_fd_sc_hd__clkbuf_16
Xclkbuf_4_11_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_11_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4657__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5690_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _6128_/A sky130_fd_sc_hd__or2_4
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _8160_/Q _7559_/Q _7431_/Q _7591_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4710_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4641_ _4639_/X _4640_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4641_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6723__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5931__B1 _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4572_ _8173_/Q _8205_/Q _8269_/Q _7777_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4572_/X sky130_fd_sc_hd__mux4_1
X_7360_ _8096_/CLK _7360_/D vssd1 vssd1 vccd1 vccd1 _7360_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold715 _8265_/Q vssd1 vssd1 vccd1 vccd1 hold715/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4003__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold737 _8452_/Q vssd1 vssd1 vccd1 vccd1 _6418_/B sky130_fd_sc_hd__dlygate4sd3_1
X_7291_ _8370_/CLK _7291_/D _7101_/Y vssd1 vssd1 vccd1 vccd1 _7291_/Q sky130_fd_sc_hd__dfrtp_2
X_6311_ _6130_/A _6307_/Y _6310_/X vssd1 vssd1 vccd1 vccd1 _6311_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold726 _5305_/X vssd1 vssd1 vccd1 vccd1 _7536_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 _6722_/X vssd1 vssd1 vccd1 vccd1 _8277_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold759 _7429_/Q vssd1 vssd1 vccd1 vccd1 hold759/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 _5292_/X vssd1 vssd1 vccd1 vccd1 _7496_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6242_ _6242_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6244_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4593__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5115__A _7076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6239__A1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6173_ _6175_/A _6175_/B vssd1 vssd1 vccd1 vccd1 _6176_/A sky130_fd_sc_hd__nand2_1
X_5124_ _5124_/A1 _4448_/B _5140_/B1 _5123_/X vssd1 vssd1 vccd1 vccd1 _7374_/D sky130_fd_sc_hd__o211a_1
Xhold1404 _4377_/B vssd1 vssd1 vccd1 vccd1 _4487_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1415 _4283_/C vssd1 vssd1 vccd1 vccd1 _4496_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_49_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8464_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1448 _4209_/Y vssd1 vssd1 vccd1 vccd1 _4210_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _7290_/Q vssd1 vssd1 vccd1 vccd1 _5136_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _5437_/A _5468_/C vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__or2_1
Xhold1426 _4345_/X vssd1 vssd1 vccd1 vccd1 _4346_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1437 _4258_/Y vssd1 vssd1 vccd1 vccd1 _4260_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4896__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4006_ _6016_/A _6013_/A vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__or2_1
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5488__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5214__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5957_ _5957_/A _5957_/B vssd1 vssd1 vccd1 vccd1 _5957_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4908_ _4907_/X _4904_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8248_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_118_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ _3974_/Y _6011_/A2 _5887_/X _7258_/A vssd1 vssd1 vccd1 vccd1 _7872_/D sky130_fd_sc_hd__a211oi_2
X_7627_ _8385_/CLK _7627_/D vssd1 vssd1 vccd1 vccd1 _7627_/Q sky130_fd_sc_hd__dfxtp_1
X_4839_ _8335_/Q _7811_/Q _7477_/Q _7445_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4839_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6714__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1467_A _7286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7558_ _8442_/CLK _7558_/D vssd1 vssd1 vccd1 vccd1 _7558_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7489_ _8402_/CLK _7489_/D vssd1 vssd1 vccd1 vccd1 _7489_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5009__B _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6509_ _6550_/A _6509_/B vssd1 vssd1 vccd1 vccd1 _6509_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4584__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6650__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7597__D _7597_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5205__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4639__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4803__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4811__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_6 _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output79_A _8124_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4774__A _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4878__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6860_ _7006_/A _6860_/A2 _6845_/B _6859_/X vssd1 vssd1 vccd1 vccd1 _6860_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_123_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5811_ _6129_/B _5811_/B _5815_/B vssd1 vssd1 vccd1 vccd1 _5811_/X sky130_fd_sc_hd__or3_1
X_6791_ _6923_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6791_/X sky130_fd_sc_hd__and2_1
XFILLER_0_29_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6944__A2 _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8530_ _8530_/A _7093_/X vssd1 vssd1 vccd1 vccd1 _8530_/Z sky130_fd_sc_hd__ebufn_1
X_5742_ _4144_/B _5742_/A2 _5786_/B _5721_/Y _5741_/X vssd1 vssd1 vccd1 vccd1 _5742_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8461_ _8461_/CLK _8461_/D vssd1 vssd1 vccd1 vccd1 _8461_/Q sky130_fd_sc_hd__dfxtp_1
X_5673_ _6545_/A _5673_/B vssd1 vssd1 vccd1 vccd1 _5673_/X sky130_fd_sc_hd__and2_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7412_ _8328_/CLK _7412_/D vssd1 vssd1 vccd1 vccd1 _7412_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5904__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4624_ _4623_/X _4620_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7514_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8392_ _8480_/CLK _8392_/D vssd1 vssd1 vccd1 vccd1 _8392_/Q sky130_fd_sc_hd__dfxtp_1
X_4555_ _8331_/Q _7807_/Q _7473_/Q _7441_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4555_/X sky130_fd_sc_hd__mux4_1
X_7343_ _8500_/CLK _7343_/D vssd1 vssd1 vccd1 vccd1 _7343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold501 _7430_/Q vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _5632_/X vssd1 vssd1 vccd1 vccd1 _7812_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold545 _7445_/Q vssd1 vssd1 vccd1 vccd1 hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _7484_/Q vssd1 vssd1 vccd1 vccd1 hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 _5316_/X vssd1 vssd1 vccd1 vccd1 _7547_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4486_ _5180_/A1 _4354_/C _5470_/C vssd1 vssd1 vccd1 vccd1 _7312_/D sky130_fd_sc_hd__mux2_1
XANTENNA__7044__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold556 _6733_/X vssd1 vssd1 vccd1 vccd1 _8288_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold578 _5282_/X vssd1 vssd1 vccd1 vccd1 _7486_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7274_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7274_/Y sky130_fd_sc_hd__inv_2
Xhold567 _7582_/Q vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4566__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6225_ _6226_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6225_/Y sky130_fd_sc_hd__nand2_1
Xhold589 _7806_/Q vssd1 vssd1 vccd1 vccd1 hold589/X sky130_fd_sc_hd__dlygate4sd3_1
X_6156_ _6157_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6156_/Y sky130_fd_sc_hd__nor2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6883__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6880__A1 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1223 _8432_/Q vssd1 vssd1 vccd1 vccd1 _6934_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 _6622_/X vssd1 vssd1 vccd1 vccd1 _8175_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 _6972_/X vssd1 vssd1 vccd1 vccd1 _8451_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _7044_/A _5538_/C vssd1 vssd1 vccd1 vccd1 _5107_/X sky130_fd_sc_hd__or2_1
Xhold1201 _8444_/Q vssd1 vssd1 vccd1 vccd1 _6958_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1245 _8338_/Q vssd1 vssd1 vccd1 vccd1 _6802_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6632__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6087_ _6105_/A2 _6078_/A _6085_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6087_/X sky130_fd_sc_hd__a22o_1
Xhold1267 _8433_/Q vssd1 vssd1 vccd1 vccd1 _6936_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 _6820_/X vssd1 vssd1 vccd1 vccd1 _8347_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5499__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1289 _5016_/X vssd1 vssd1 vccd1 vccd1 _7320_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1278 _8356_/Q vssd1 vssd1 vccd1 vccd1 _6838_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5038_ _4403_/A _4407_/B _5166_/B1 _5037_/X vssd1 vssd1 vccd1 vccd1 _5038_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5199__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4623__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6989_ _5382_/B _6988_/X _6981_/Y vssd1 vssd1 vccd1 vccd1 _6989_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6148__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6699__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput65 _8111_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[10] sky130_fd_sc_hd__buf_12
Xoutput76 _8121_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[20] sky130_fd_sc_hd__buf_12
XANTENNA__6793__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput87 _8131_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[30] sky130_fd_sc_hd__buf_12
Xoutput98 _7293_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[11] sky130_fd_sc_hd__buf_12
Xhold1790 _5787_/X vssd1 vssd1 vccd1 vccd1 _5788_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output117_A _7284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3938__A _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4533__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5362__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4769__A _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3912__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4340_ _4339_/X _4379_/A _5470_/B vssd1 vssd1 vccd1 vccd1 _4341_/C sky130_fd_sc_hd__mux2_1
X_4271_ _8500_/Q _4271_/B vssd1 vssd1 vccd1 vccd1 _4271_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4548__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6862__A1 _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6010_ _5734_/A _5996_/X _6009_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6010_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_118_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6614__A1 _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4708__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7961_ _8020_/CLK _7961_/D vssd1 vssd1 vccd1 vccd1 _7961_/Q sky130_fd_sc_hd__dfxtp_1
X_6912_ _3939_/C _6943_/B _6911_/X vssd1 vssd1 vccd1 vccd1 _6912_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3979__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7892_ _8504_/CLK _7892_/D vssd1 vssd1 vccd1 vccd1 _7892_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4720__S0 _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6843_ _6911_/A _6843_/B _6901_/B vssd1 vssd1 vccd1 vccd1 _6843_/X sky130_fd_sc_hd__or3_1
X_7251__129 _8487_/CLK vssd1 vssd1 vccd1 vccd1 _8261_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6774_ _6971_/A _6741_/B _6774_/B1 hold617/X vssd1 vssd1 vccd1 vccd1 _6774_/X sky130_fd_sc_hd__a22o_1
X_3986_ _3923_/B _7944_/Q vssd1 vssd1 vccd1 vccd1 _3986_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_57_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6224__A _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5050__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8513_ _8513_/CLK _8513_/D vssd1 vssd1 vccd1 vccd1 _8513_/Q sky130_fd_sc_hd__dfxtp_1
X_5725_ _8455_/Q _5730_/A _4153_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _5725_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5656_ _6999_/A _5656_/B vssd1 vssd1 vccd1 vccd1 _7836_/D sky130_fd_sc_hd__and2_1
XANTENNA_fanout315_A _5186_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8444_ _8480_/CLK _8444_/D vssd1 vssd1 vccd1 vccd1 _8444_/Q sky130_fd_sc_hd__dfxtp_1
X_4607_ _8178_/Q _8210_/Q _8274_/Q _7782_/Q _4611_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4607_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_115_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5353__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4787__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5587_ _3939_/C _5585_/B _5585_/Y hold240/X vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__o22a_1
Xhold320 _7314_/Q vssd1 vssd1 vccd1 vccd1 _5411_/A sky130_fd_sc_hd__dlygate4sd3_1
X_8375_ _8378_/CLK _8375_/D _7269_/Y vssd1 vssd1 vccd1 vccd1 _8375_/Q sky130_fd_sc_hd__dfrtp_1
X_4538_ _8458_/Q _8390_/Q _8422_/Q _8296_/Q _4611_/S0 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4538_/X sky130_fd_sc_hd__mux4_1
Xhold342 _8210_/Q vssd1 vssd1 vccd1 vccd1 hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 _5264_/X vssd1 vssd1 vccd1 vccd1 _7468_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7326_ _8034_/CLK _7326_/D vssd1 vssd1 vccd1 vccd1 _7326_/Q sky130_fd_sc_hd__dfxtp_1
Xhold331 _5414_/X vssd1 vssd1 vccd1 vccd1 _7603_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold364 _7321_/Q vssd1 vssd1 vccd1 vccd1 _5418_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7257_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7257_/Y sky130_fd_sc_hd__inv_2
Xhold386 _8158_/Q vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4469_ _7018_/A _7918_/Q vssd1 vssd1 vccd1 vccd1 _8050_/D sky130_fd_sc_hd__and2_1
Xhold375 _5455_/X vssd1 vssd1 vccd1 vccd1 _7644_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 _5647_/X vssd1 vssd1 vccd1 vccd1 _7827_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _6209_/A _6209_/B vssd1 vssd1 vccd1 vccd1 _6208_/Y sky130_fd_sc_hd__nor2_1
Xhold1042 _5198_/X vssd1 vssd1 vccd1 vccd1 _7412_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6139_ _6140_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6139_/Y sky130_fd_sc_hd__nor2_1
Xhold1031 _8476_/Q vssd1 vssd1 vccd1 vccd1 _7018_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1020 _6700_/X vssd1 vssd1 vccd1 vccd1 _8227_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1053 _8228_/Q vssd1 vssd1 vccd1 vccd1 _6701_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 _7799_/Q vssd1 vssd1 vccd1 vccd1 _5615_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 _6565_/X vssd1 vssd1 vccd1 vccd1 _8137_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1097 _8279_/Q vssd1 vssd1 vccd1 vccd1 _6724_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 _5321_/X vssd1 vssd1 vccd1 vccd1 _7552_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3758__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4353__S _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5592__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5973__A _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5344__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6844__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5647__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3940__B _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6309__A _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4702__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5867__B _5971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5280__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3830__A1 _4773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4771__B _4771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3840_ _3840_/A0 _6452_/B _4074_/S vssd1 vssd1 vccd1 vccd1 _4118_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5032__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3771_ _4761_/B _3966_/B vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__nand2_1
X_5510_ _7531_/Q _5542_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7699_/D sky130_fd_sc_hd__and3_1
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6490_ _7006_/A _6490_/B vssd1 vssd1 vccd1 vccd1 _6490_/X sky130_fd_sc_hd__and2_1
XFILLER_0_81_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5441_ _5441_/A _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5441_/X sky130_fd_sc_hd__and3_1
XFILLER_0_30_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5372_ _5404_/A _7344_/Q vssd1 vssd1 vccd1 vccd1 _5392_/B sky130_fd_sc_hd__or2_1
XFILLER_0_1_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8160_ _8160_/CLK _8160_/D vssd1 vssd1 vccd1 vccd1 _8160_/Q sky130_fd_sc_hd__dfxtp_1
X_7111_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7111_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5107__B _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8091_ _8091_/CLK _8125_/D vssd1 vssd1 vccd1 vccd1 _8091_/Q sky130_fd_sc_hd__dfxtp_1
X_4323_ _8493_/Q _4323_/B vssd1 vssd1 vccd1 vccd1 _4323_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7042_ _7079_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7042_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5638__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4254_ _4253_/X _4412_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _4413_/B sky130_fd_sc_hd__mux2_1
X_4185_ _4440_/B vssd1 vssd1 vccd1 vccd1 _4193_/B sky130_fd_sc_hd__inv_2
XANTENNA__4941__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7944_ _8360_/CLK _7944_/D vssd1 vssd1 vccd1 vccd1 _7944_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5271__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4074__A1 _4073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7875_ _8454_/CLK _7875_/D vssd1 vssd1 vccd1 vccd1 _7875_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5496__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout432_A _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6826_ _7025_/A _6826_/A2 _6838_/A3 _6825_/X vssd1 vssd1 vccd1 vccd1 _6826_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_92_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6757_ _6937_/A _6741_/B _6774_/B1 hold485/X vssd1 vssd1 vccd1 vccd1 _6757_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6889__A _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4901__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3969_ _4074_/S _3967_/X _3968_/X vssd1 vssd1 vccd1 vccd1 _6307_/A sky130_fd_sc_hd__a21oi_4
X_5708_ _6209_/A _6226_/A _5716_/S vssd1 vssd1 vccd1 vccd1 _5708_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6771__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6688_ _6877_/A _6669_/B _6702_/B1 hold855/X vssd1 vssd1 vccd1 vccd1 _6688_/X sky130_fd_sc_hd__a22o_1
X_5639_ _6877_/A _5620_/B _5653_/B1 hold961/X vssd1 vssd1 vccd1 vccd1 _5639_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5326__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8427_ _8427_/CLK _8427_/D vssd1 vssd1 vccd1 vccd1 _8427_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7190__68 _8328_/CLK vssd1 vssd1 vccd1 vccd1 _8103_/CLK sky130_fd_sc_hd__inv_2
X_8358_ _8358_/CLK _8358_/D _7252_/Y vssd1 vssd1 vccd1 vccd1 _8358_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5877__A2 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5017__B _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 _6487_/X vssd1 vssd1 vccd1 vccd1 _7969_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7309_ _8385_/CLK _7309_/D _7119_/Y vssd1 vssd1 vccd1 vccd1 _7309_/Q sky130_fd_sc_hd__dfrtp_4
Xhold150 _7625_/Q vssd1 vssd1 vccd1 vccd1 _5683_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _6489_/X vssd1 vssd1 vccd1 vccd1 _7971_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _7839_/Q vssd1 vssd1 vccd1 vccd1 _6460_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5629__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6826__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold172 _7614_/Q vssd1 vssd1 vccd1 vccd1 _5672_/B sky130_fd_sc_hd__dlygate4sd3_1
X_8289_ _8483_/CLK _8289_/D vssd1 vssd1 vccd1 vccd1 _8289_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3760__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6129__A _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5014__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6357__A3 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6762__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6799__A _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5317__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3879__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3951__A _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4923__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6045__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5990_ _5990_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _5993_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5253__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3803__A1 _3802_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4941_ _8479_/Q _8411_/Q _8443_/Q _8317_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4941_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7660_ _8080_/CLK _7660_/D vssd1 vssd1 vccd1 vccd1 _7660_/Q sky130_fd_sc_hd__dfxtp_1
X_4872_ _4871_/X _4870_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4872_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3823_ _3823_/A _3823_/B vssd1 vssd1 vccd1 vccd1 _3848_/B sky130_fd_sc_hd__and2_1
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6611_ _6917_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6611_/X sky130_fd_sc_hd__and2_1
XANTENNA__6753__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7591_ _8442_/CLK _7591_/D vssd1 vssd1 vccd1 vccd1 _7591_/Q sky130_fd_sc_hd__dfxtp_1
X_6542_ _6706_/A _6542_/B vssd1 vssd1 vccd1 vccd1 _8024_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3754_ _8083_/Q _3753_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3754_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4721__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3845__B _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3685_ _3685_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3685_/X sky130_fd_sc_hd__or2_1
XANTENNA__5308__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6473_ _7022_/A _6473_/B vssd1 vssd1 vccd1 vccd1 _6473_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8212_ _8402_/CLK _8212_/D vssd1 vssd1 vccd1 vccd1 _8212_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5424_ _5424_/A _5503_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _5424_/X sky130_fd_sc_hd__and3_1
XFILLER_0_30_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8143_ _8143_/CLK _8143_/D vssd1 vssd1 vccd1 vccd1 _8143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6808__A1 _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5355_ _6945_/A _5367_/A2 _5367_/B1 hold567/X vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__a22o_1
X_8074_ _8500_/CLK _8108_/D vssd1 vssd1 vccd1 vccd1 _8074_/Q sky130_fd_sc_hd__dfxtp_1
X_5286_ _6953_/A _5294_/A2 _5294_/B1 hold791/X vssd1 vssd1 vccd1 vccd1 _5286_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4306_ _4307_/A _7652_/Q vssd1 vssd1 vccd1 vccd1 _4308_/A sky130_fd_sc_hd__or2_1
XANTENNA_fanout382_A _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4237_ _4235_/Y _4237_/B vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__6284__A2 _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7052__B _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7025_ _7025_/A _7025_/B vssd1 vssd1 vccd1 vccd1 _7025_/X sky130_fd_sc_hd__and2_1
XANTENNA__5389__C_N _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5788__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4168_ _4166_/Y _4168_/B vssd1 vssd1 vccd1 vccd1 _4169_/B sky130_fd_sc_hd__and2b_1
XANTENNA__6891__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_4_clk_A clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4099_ _5946_/A _5943_/A vssd1 vssd1 vccd1 vccd1 _4099_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_78_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5244__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7927_ _8368_/CLK _7927_/D vssd1 vssd1 vccd1 vccd1 _7927_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5795__A1 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7858_ _8020_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 _7858_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6809_ _6941_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6809_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7789_ _8475_/CLK _7789_/D vssd1 vssd1 vccd1 vccd1 _7789_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4631__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3755__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3771__A _4761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6275__A2 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4905__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 _3646_/Y vssd1 vssd1 vccd1 vccd1 _6660_/A1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3710__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4806__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6735__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold919 _7569_/Q vssd1 vssd1 vccd1 vccd1 hold919/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold908 _5315_/X vssd1 vssd1 vccd1 vccd1 _7546_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5140_ _5140_/A1 _4448_/B _5140_/B1 _5139_/X vssd1 vssd1 vccd1 vccd1 _7382_/D sky130_fd_sc_hd__o211a_1
XANTENNA__3721__B1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5071_ _6553_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5071_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1608 _4250_/Y vssd1 vssd1 vccd1 vccd1 _4251_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4022_ _7283_/Q _7950_/Q vssd1 vssd1 vccd1 vccd1 _4022_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_36_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1619 _4323_/Y vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_126_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4029__A1 _4028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5973_ _5974_/A _5974_/B vssd1 vssd1 vccd1 vccd1 _5973_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5777__A1 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7712_ _8143_/CLK _7712_/D vssd1 vssd1 vccd1 vccd1 _7712_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4924_ _8154_/Q _7553_/Q _7425_/Q _7585_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4924_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_35_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4855_ _4853_/X _4854_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4855_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6726__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7643_ _8373_/CLK _7643_/D vssd1 vssd1 vccd1 vccd1 _7643_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4786_ _8167_/Q _8199_/Q _8263_/Q _7771_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4786_/X sky130_fd_sc_hd__mux4_1
X_7574_ _8343_/CLK _7574_/D vssd1 vssd1 vccd1 vccd1 _7574_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout228_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3806_ _4774_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3806_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3737_ _6279_/A _6281_/A vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__or2_1
X_6525_ _6550_/A _6525_/B vssd1 vssd1 vccd1 vccd1 _8007_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6456_ _7835_/Q _7938_/Q _6911_/A vssd1 vssd1 vccd1 vccd1 _6456_/X sky130_fd_sc_hd__mux2_1
X_3668_ _7835_/Q _3658_/Y _3665_/X _3666_/Y _3667_/X vssd1 vssd1 vccd1 vccd1 _3669_/B
+ sky130_fd_sc_hd__o2111a_1
X_7160__38 _8029_/CLK vssd1 vssd1 vccd1 vccd1 _8040_/CLK sky130_fd_sc_hd__inv_2
X_5407_ _7079_/C _5548_/B vssd1 vssd1 vccd1 vccd1 _7069_/B sky130_fd_sc_hd__nand2_4
XANTENNA__5701__A1 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6387_ _6388_/A _6388_/B vssd1 vssd1 vccd1 vccd1 _6387_/X sky130_fd_sc_hd__and2_1
X_5338_ _3939_/C _5336_/B _5336_/Y hold246/X vssd1 vssd1 vccd1 vccd1 _5338_/X sky130_fd_sc_hd__o22a_1
X_8126_ _8126_/CLK _8126_/D vssd1 vssd1 vccd1 vccd1 _8126_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__7063__A _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8057_ _8057_/CLK _8057_/D vssd1 vssd1 vccd1 vccd1 _8057_/Q sky130_fd_sc_hd__dfxtp_1
X_7008_ _7008_/A _7008_/B vssd1 vssd1 vccd1 vccd1 _7008_/X sky130_fd_sc_hd__and2_1
X_5269_ _6853_/A _5262_/B _5295_/B1 hold541/X vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5217__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5768__A1 _5971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6126__B _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6717__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6248__A2 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout290 _6703_/Y vssd1 vssd1 vccd1 vccd1 _6705_/B sky130_fd_sc_hd__buf_8
XANTENNA__4536__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6317__A _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5208__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3676__A _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ _8150_/Q _7549_/Q _7421_/Q _7581_/Q _4640_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4640_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_84_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6184__B2 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5891__A _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6310_ _6414_/A2 _6301_/A _6309_/Y _5759_/Y _6308_/X vssd1 vssd1 vccd1 vccd1 _6310_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4571_ _4569_/X _4570_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4571_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold716 _6710_/X vssd1 vssd1 vccd1 vccd1 _8265_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3942__B1 _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7290_ _7977_/CLK _7290_/D _7100_/Y vssd1 vssd1 vccd1 vccd1 _7290_/Q sky130_fd_sc_hd__dfrtp_1
Xhold705 _7403_/Q vssd1 vssd1 vccd1 vccd1 _5470_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold727 _7774_/Q vssd1 vssd1 vccd1 vccd1 hold727/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold738 _6418_/X vssd1 vssd1 vccd1 vccd1 _7900_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6198__S _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6241_ _6225_/Y _6229_/B _6227_/B vssd1 vssd1 vccd1 vccd1 _6247_/A sky130_fd_sc_hd__a21o_1
Xhold749 _7584_/Q vssd1 vssd1 vccd1 vccd1 hold749/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6172_ _6172_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6175_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4593__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5115__B _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5123_ _5441_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5123_/X sky130_fd_sc_hd__or2_1
Xhold1405 _7885_/Q vssd1 vssd1 vccd1 vccd1 hold1405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 _4397_/X vssd1 vssd1 vccd1 vccd1 _4399_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1449 _4218_/X vssd1 vssd1 vccd1 vccd1 _4219_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5054_ _4382_/A _5069_/S _5182_/B1 _5053_/X vssd1 vssd1 vccd1 vccd1 _5054_/X sky130_fd_sc_hd__o211a_1
Xhold1427 _4346_/X vssd1 vssd1 vccd1 vccd1 _5578_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 _4260_/X vssd1 vssd1 vccd1 vccd1 _5566_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4005_ _4208_/A _4004_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _6013_/A sky130_fd_sc_hd__mux2_2
XANTENNA_fanout178_A _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7205__83 _8510_/CLK vssd1 vssd1 vccd1 vccd1 _8118_/CLK sky130_fd_sc_hd__inv_2
XANTENNA_fanout345_A _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5956_ _6126_/A _6270_/A vssd1 vssd1 vccd1 vccd1 _5957_/B sky130_fd_sc_hd__nand2_1
X_5887_ _5734_/A _5872_/Y _5886_/X vssd1 vssd1 vccd1 vccd1 _5887_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_48_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6962__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4907_ _4906_/X _4905_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4838_ _4837_/X _4834_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8238_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7626_ _8494_/CLK _7626_/D vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7557_ _8413_/CLK _7557_/D vssd1 vssd1 vccd1 vccd1 _7557_/Q sky130_fd_sc_hd__dfxtp_1
X_4769_ _7026_/A _4769_/B vssd1 vssd1 vccd1 vccd1 _8126_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6897__A _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7488_ _8440_/CLK _7488_/D vssd1 vssd1 vccd1 vccd1 _7488_/Q sky130_fd_sc_hd__dfxtp_1
X_6508_ _7027_/A hold19/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__and2_1
X_6439_ _6999_/A _6439_/B vssd1 vssd1 vccd1 vccd1 _7921_/D sky130_fd_sc_hd__and2_1
XFILLER_0_30_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4584__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8109_ _8109_/CLK _8109_/D vssd1 vssd1 vccd1 vccd1 _8109_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5150__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5610__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6166__B2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5913__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5913__A1 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_91_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3924__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 _6453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6790_ _7008_/A _6790_/A2 _6779_/B _6789_/X vssd1 vssd1 vccd1 vccd1 _6790_/X sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_44_clk_A _7871_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5810_ _6270_/A _5810_/B vssd1 vssd1 vccd1 vccd1 _5815_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_123_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5741_ _6028_/S _5879_/S _4095_/A _5740_/Y _5736_/Y vssd1 vssd1 vccd1 vccd1 _5741_/X
+ sky130_fd_sc_hd__o41a_1
XANTENNA__5601__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7129__7 _8343_/CLK vssd1 vssd1 vccd1 vccd1 _7506_/CLK sky130_fd_sc_hd__inv_2
X_8460_ _8460_/CLK _8460_/D vssd1 vssd1 vccd1 vccd1 _8460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7411_ _8354_/CLK _7411_/D vssd1 vssd1 vccd1 vccd1 _7411_/Q sky130_fd_sc_hd__dfxtp_1
X_5672_ _7022_/A _5672_/B vssd1 vssd1 vccd1 vccd1 _5672_/X sky130_fd_sc_hd__and2_1
XFILLER_0_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8391_ _8468_/CLK _8391_/D vssd1 vssd1 vccd1 vccd1 _8391_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_59_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4623_ _4622_/X _4621_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3915__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7342_ _8030_/CLK _7342_/D vssd1 vssd1 vccd1 vccd1 _7342_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6510__A _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4554_ _4553_/X _4550_/X _7365_/Q vssd1 vssd1 vccd1 vccd1 _7504_/D sky130_fd_sc_hd__mux2_1
Xhold502 _5216_/X vssd1 vssd1 vccd1 vccd1 _7430_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_102_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold513 _7779_/Q vssd1 vssd1 vccd1 vccd1 hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 _5280_/X vssd1 vssd1 vccd1 vccd1 _7484_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7273_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7273_/Y sky130_fd_sc_hd__inv_2
Xhold535 _7459_/Q vssd1 vssd1 vccd1 vccd1 hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _8458_/Q vssd1 vssd1 vccd1 vccd1 _7000_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _5237_/X vssd1 vssd1 vccd1 vccd1 _7445_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4030__A _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4485_ _5182_/A1 _4372_/B _5470_/C vssd1 vssd1 vccd1 vccd1 _7313_/D sky130_fd_sc_hd__mux2_1
Xhold557 _7575_/Q vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
X_6224_ _6226_/A _6226_/B vssd1 vssd1 vccd1 vccd1 _6227_/A sky130_fd_sc_hd__and2_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold568 _5355_/X vssd1 vssd1 vccd1 vccd1 _7582_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4566__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5132__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4110__A_N _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout295_A _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6155_ _6157_/A _6157_/B vssd1 vssd1 vccd1 vccd1 _6155_/Y sky130_fd_sc_hd__nand2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1224 _6934_/X vssd1 vssd1 vccd1 vccd1 _8432_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1213 _8423_/Q vssd1 vssd1 vccd1 vccd1 _6916_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5106_ input14/X _5099_/B _5148_/B1 _5105_/X vssd1 vssd1 vccd1 vccd1 _7365_/D sky130_fd_sc_hd__o211a_1
X_6086_ _4089_/A _6398_/A2 _5732_/X _6072_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _6086_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1202 _6958_/X vssd1 vssd1 vccd1 vccd1 _8444_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 _6802_/X vssd1 vssd1 vccd1 vccd1 _8338_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 _8419_/Q vssd1 vssd1 vccd1 vccd1 _6906_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _8177_/Q vssd1 vssd1 vccd1 vccd1 _6626_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5037_ _5428_/A _5540_/C vssd1 vssd1 vccd1 vccd1 _5037_/X sky130_fd_sc_hd__or2_1
Xhold1268 _6936_/X vssd1 vssd1 vccd1 vccd1 _8433_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout462_A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1279 _6838_/X vssd1 vssd1 vccd1 vccd1 _8356_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5499__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5199__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6396__A1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4904__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6988_ _7067_/A _5386_/B _6597_/B _6987_/X _6595_/Y vssd1 vssd1 vccd1 vccd1 _6988_/X
+ sky130_fd_sc_hd__a221o_1
X_5939_ _5937_/X _5938_/X _6028_/S vssd1 vssd1 vccd1 vccd1 _5939_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6404__B _6406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7609_ _7907_/CLK _7609_/D vssd1 vssd1 vccd1 vccd1 _7609_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6699__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_10_0_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__6420__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1744_A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput66 _8112_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[11] sky130_fd_sc_hd__buf_12
Xoutput88 _8132_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[31] sky130_fd_sc_hd__buf_12
Xoutput99 _7294_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[12] sky130_fd_sc_hd__buf_12
Xoutput77 _8122_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[21] sky130_fd_sc_hd__buf_12
XANTENNA__5831__A0 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1780 _6115_/A vssd1 vssd1 vccd1 vccd1 _4076_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1791 _7704_/Q vssd1 vssd1 vccd1 vccd1 _3971_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6926__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7196__74 _8510_/CLK vssd1 vssd1 vccd1 vccd1 _8109_/CLK sky130_fd_sc_hd__inv_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output91_A _8106_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5362__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4133__A_N _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5114__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5745__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6311__A1 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4270_ _8500_/Q _4271_/B vssd1 vssd1 vccd1 vccd1 _4270_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4548__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7960_ _8503_/CLK _7960_/D vssd1 vssd1 vccd1 vccd1 _7960_/Q sky130_fd_sc_hd__dfxtp_1
X_6911_ _6911_/A _6911_/B _6963_/B vssd1 vssd1 vccd1 vccd1 _6911_/X sky130_fd_sc_hd__or3_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7891_ _8463_/CLK _7891_/D vssd1 vssd1 vccd1 vccd1 _7891_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4720__S1 _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6842_ _7939_/Q _7940_/Q _6842_/C vssd1 vssd1 vccd1 vccd1 _6842_/X sky130_fd_sc_hd__or3_4
XFILLER_0_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6378__A1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3985_ _3985_/A _3985_/B vssd1 vssd1 vccd1 vccd1 _3985_/X sky130_fd_sc_hd__and2_1
XFILLER_0_57_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6773_ _6969_/A _6773_/A2 _6773_/B1 _6773_/B2 vssd1 vssd1 vccd1 vccd1 _6773_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_134_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8512_ _8515_/CLK _8512_/D vssd1 vssd1 vccd1 vccd1 _8512_/Q sky130_fd_sc_hd__dfxtp_1
X_5724_ _5738_/A _5730_/A vssd1 vssd1 vccd1 vccd1 _5732_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_45_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5655_ _6999_/A _5655_/B vssd1 vssd1 vccd1 vccd1 _7835_/D sky130_fd_sc_hd__and2_1
XFILLER_0_45_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8443_ _8476_/CLK _8443_/D vssd1 vssd1 vccd1 vccd1 _8443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4606_ _4604_/X _4605_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4606_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8374_ _8378_/CLK _8374_/D _7268_/Y vssd1 vssd1 vccd1 vccd1 _8374_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4787__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5586_ _6777_/A _5585_/B _5585_/Y hold312/X vssd1 vssd1 vccd1 vccd1 _5586_/X sky130_fd_sc_hd__o22a_1
X_7325_ _8034_/CLK _7325_/D vssd1 vssd1 vccd1 vccd1 _7325_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout308_A _5333_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7055__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5353__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold310 _7392_/Q vssd1 vssd1 vccd1 vccd1 _5459_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ _8168_/Q _8200_/Q _8264_/Q _7772_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4537_/X sky130_fd_sc_hd__mux4_1
Xhold343 _6683_/X vssd1 vssd1 vccd1 vccd1 _8210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _7384_/Q vssd1 vssd1 vccd1 vccd1 _5451_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _5411_/X vssd1 vssd1 vccd1 vccd1 _7600_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold365 _5418_/X vssd1 vssd1 vccd1 vccd1 _7607_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7256_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7256_/Y sky130_fd_sc_hd__inv_2
Xhold387 _6586_/X vssd1 vssd1 vccd1 vccd1 _8158_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _7461_/Q vssd1 vssd1 vccd1 vccd1 hold376/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4468_ _7023_/A _7919_/Q vssd1 vssd1 vccd1 vccd1 _8051_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold354 _7828_/Q vssd1 vssd1 vccd1 vccd1 hold354/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold398 _7543_/Q vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _6209_/A _6209_/B vssd1 vssd1 vccd1 vccd1 _6210_/A sky130_fd_sc_hd__nand2_1
X_6138_ _6140_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6141_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3803__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4399_ _5042_/A1 _4407_/B _4399_/B1 _4398_/Y vssd1 vssd1 vccd1 vccd1 _8377_/D sky130_fd_sc_hd__a22o_1
Xhold1010 _6998_/X vssd1 vssd1 vccd1 vccd1 _8456_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1032 _7018_/X vssd1 vssd1 vccd1 vccd1 _8476_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 _8266_/Q vssd1 vssd1 vccd1 vccd1 _6711_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1065 _8142_/Q vssd1 vssd1 vccd1 vccd1 _6570_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 _8473_/Q vssd1 vssd1 vccd1 vccd1 _7015_/B sky130_fd_sc_hd__dlygate4sd3_1
X_6069_ _5694_/Y _6068_/X _6067_/X vssd1 vssd1 vccd1 vccd1 _6069_/Y sky130_fd_sc_hd__a21oi_1
Xhold1054 _6701_/X vssd1 vssd1 vccd1 vccd1 _8228_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 _5615_/X vssd1 vssd1 vccd1 vccd1 _7799_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 _6724_/X vssd1 vssd1 vccd1 vccd1 _8279_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 _8480_/Q vssd1 vssd1 vccd1 vccd1 _7022_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4634__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5592__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5344__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6844__A2 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4809__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5280__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4702__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3830__A2 _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6780__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3770_ _4083_/B _3941_/B _6877_/A vssd1 vssd1 vccd1 vccd1 _3770_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5440_ _5440_/A _7030_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _5440_/X sky130_fd_sc_hd__and3_1
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5371_ _7065_/A _7067_/A _7069_/A vssd1 vssd1 vccd1 vccd1 _6974_/A sky130_fd_sc_hd__or3_2
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7110_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7110_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8090_ _8090_/CLK _8124_/D vssd1 vssd1 vccd1 vccd1 _8090_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4322_ _8493_/Q _4323_/B vssd1 vssd1 vccd1 vccd1 _4322_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7041_ _7031_/Y _7041_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8493_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4253_ _4253_/A _4253_/B vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__xor2_1
XANTENNA__5404__A _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4184_ _4183_/Y hold212/X _7082_/A vssd1 vssd1 vccd1 vccd1 _4440_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4941__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6143__S0 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7943_ _8030_/CLK _7943_/D vssd1 vssd1 vccd1 vccd1 _7943_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5271__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7874_ _8339_/CLK _7874_/D vssd1 vssd1 vccd1 vccd1 _7874_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout258_A _5335_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6235__A _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6825_ _6891_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6825_/X sky130_fd_sc_hd__and2_1
XFILLER_0_108_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6756_ _6935_/A _6741_/B _6774_/B1 hold845/X vssd1 vssd1 vccd1 vccd1 _6756_/X sky130_fd_sc_hd__a22o_1
X_3968_ _3968_/A _3968_/B vssd1 vssd1 vccd1 vccd1 _3968_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout425_A _7283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6771__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5707_ _5705_/X _5706_/X _5838_/A vssd1 vssd1 vccd1 vccd1 _5707_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6889__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3899_ _7974_/Q _4079_/A2 _4079_/B1 _8006_/Q _3898_/X vssd1 vssd1 vccd1 vccd1 _3899_/X
+ sky130_fd_sc_hd__a221o_2
X_6687_ _6941_/A _6669_/B _6702_/B1 hold707/X vssd1 vssd1 vccd1 vccd1 _6687_/X sky130_fd_sc_hd__a22o_1
X_8426_ _8426_/CLK _8426_/D vssd1 vssd1 vccd1 vccd1 _8426_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5326__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5638_ _6941_/A _5652_/A2 _5652_/B1 hold829/X vssd1 vssd1 vccd1 vccd1 _5638_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8357_ _8487_/CLK _8357_/D vssd1 vssd1 vccd1 vccd1 _8357_/Q sky130_fd_sc_hd__dfxtp_1
X_5569_ _6550_/A _5569_/B vssd1 vssd1 vccd1 vccd1 _7758_/D sky130_fd_sc_hd__and2_1
XANTENNA__3888__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold140 _7742_/Q vssd1 vssd1 vccd1 vccd1 _6493_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 _7768_/Q vssd1 vssd1 vccd1 vccd1 _6519_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _5683_/X vssd1 vssd1 vccd1 vccd1 _7863_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7308_ _8382_/CLK _7308_/D _7118_/Y vssd1 vssd1 vccd1 vccd1 _7308_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA_hold1442_A _7303_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold195 _6460_/X vssd1 vssd1 vccd1 vccd1 _7942_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _7840_/Q vssd1 vssd1 vccd1 vccd1 _6461_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _5672_/X vssd1 vssd1 vccd1 vccd1 _7852_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8288_ _8479_/CLK _8288_/D vssd1 vssd1 vccd1 vccd1 _8288_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6039__A0 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4696__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6762__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7166__44 _8465_/CLK vssd1 vssd1 vccd1 vccd1 _8046_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6799__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5317__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3879__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4539__S _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4923__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4056__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5253__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3679__A _7282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6055__A _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4940_ _8189_/Q _8221_/Q _8285_/Q _7793_/Q _4990_/S0 _4990_/S1 vssd1 vssd1 vccd1
+ vccd1 _4940_/X sky130_fd_sc_hd__mux4_1
X_4871_ _8469_/Q _8401_/Q _8433_/Q _8307_/Q _4997_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4871_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_47_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6610_ _7010_/A _6610_/A2 _6602_/X _6609_/X vssd1 vssd1 vccd1 vccd1 _6610_/X sky130_fd_sc_hd__a31o_1
X_3822_ _6350_/A _6352_/A vssd1 vssd1 vccd1 vccd1 _3823_/B sky130_fd_sc_hd__nand2_1
X_7590_ _8486_/CLK _7590_/D vssd1 vssd1 vccd1 vccd1 _7590_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6753__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6541_ _6550_/A _6541_/B vssd1 vssd1 vccd1 vccd1 _8023_/D sky130_fd_sc_hd__and2_1
XFILLER_0_82_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3753_ _7987_/Q _4068_/A2 _4068_/B1 _8019_/Q _3752_/X vssd1 vssd1 vccd1 vccd1 _3753_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_131_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3684_ _3669_/A _3669_/B _3676_/B vssd1 vssd1 vccd1 vccd1 _3841_/B sky130_fd_sc_hd__a21o_2
XANTENNA__5308__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6472_ _6545_/A hold39/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__and2_1
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5423_ _5423_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5423_/X sky130_fd_sc_hd__and3_1
X_8211_ _8469_/CLK _8211_/D vssd1 vssd1 vccd1 vccd1 _8211_/Q sky130_fd_sc_hd__dfxtp_1
X_8142_ _8343_/CLK _8142_/D vssd1 vssd1 vccd1 vccd1 _8142_/Q sky130_fd_sc_hd__dfxtp_1
X_5354_ _6877_/A _5335_/B _5368_/B1 hold807/X vssd1 vssd1 vccd1 vccd1 _5354_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4611__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4305_ _4398_/A _4395_/B _4392_/B vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__and3_1
X_8073_ _8143_/CLK _8073_/D vssd1 vssd1 vccd1 vccd1 _8073_/Q sky130_fd_sc_hd__dfxtp_1
X_5285_ _6951_/A _5262_/B _5295_/B1 hold811/X vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__a22o_1
X_4236_ _8505_/Q _7642_/Q vssd1 vssd1 vccd1 vccd1 _4237_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6284__A3 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7024_ _7024_/A _7024_/B vssd1 vssd1 vccd1 vccd1 _7024_/X sky130_fd_sc_hd__and2_1
X_4167_ _8515_/Q _7632_/Q vssd1 vssd1 vccd1 vccd1 _4168_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout375_A hold1637/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4047__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4098_ _5846_/A _6342_/S _5820_/A _4097_/Y _4096_/Y vssd1 vssd1 vccd1 vccd1 _4098_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5244__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4678__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4184__S _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5795__A2 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7926_ _8480_/CLK _7926_/D vssd1 vssd1 vccd1 vccd1 _7926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7857_ _8504_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _7857_/Q sky130_fd_sc_hd__dfxtp_1
X_6808_ _6434_/A _6808_/A2 _6838_/A3 _6807_/X vssd1 vssd1 vccd1 vccd1 _6808_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_135_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6744__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7788_ _8346_/CLK _7788_/D vssd1 vssd1 vccd1 vccd1 _7788_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6739_ _7939_/Q _7940_/Q _6740_/C vssd1 vssd1 vccd1 vccd1 _6739_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__4850__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8409_ _8477_/CLK _8409_/D vssd1 vssd1 vccd1 vccd1 _8409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5180__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3771__B _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout450 _4775_/A vssd1 vssd1 vccd1 vccd1 _6706_/A sky130_fd_sc_hd__buf_4
XANTENNA__6680__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout461 input63/X vssd1 vssd1 vccd1 vccd1 _7267_/A sky130_fd_sc_hd__buf_8
XFILLER_0_45_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4905__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6603__A _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6735__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold909 _8478_/Q vssd1 vssd1 vccd1 vccd1 _7020_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3681__B _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3721__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5070_ _7279_/A _5070_/B _5470_/B vssd1 vssd1 vccd1 vccd1 _7347_/D sky130_fd_sc_hd__or3b_1
X_4021_ _4021_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _4045_/B sky130_fd_sc_hd__and2_1
Xhold1609 _4251_/Y vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ _5974_/A _5974_/B vssd1 vssd1 vccd1 vccd1 _5975_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5777__A2 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4923_ _8347_/Q _7823_/Q _7489_/Q _7457_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4923_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7711_ _8448_/CLK _7711_/D vssd1 vssd1 vccd1 vccd1 _7711_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4017__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4732__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7642_ _8369_/CLK _7642_/D vssd1 vssd1 vccd1 vccd1 _7642_/Q sky130_fd_sc_hd__dfxtp_1
X_4854_ _8144_/Q _7543_/Q _7415_/Q _7575_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4854_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6187__C1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6513__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6726__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4785_ _4783_/X _4784_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__mux2_1
X_7573_ _8175_/CLK _7573_/D vssd1 vssd1 vccd1 vccd1 _7573_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3805_ _4774_/B _4071_/A2 _4071_/B1 _6969_/A _3804_/X vssd1 vssd1 vccd1 vccd1 _6388_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_132_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4832__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3736_ _6279_/A _6281_/A vssd1 vssd1 vccd1 vccd1 _3736_/Y sky130_fd_sc_hd__nand2_1
X_6524_ _6524_/A _6524_/B vssd1 vssd1 vccd1 vccd1 _8006_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3667_ _7834_/Q _3659_/Y _3663_/X _7902_/Q vssd1 vssd1 vccd1 vccd1 _3667_/X sky130_fd_sc_hd__o211a_1
X_6455_ _7834_/Q _7937_/Q _6911_/A vssd1 vssd1 vccd1 vccd1 _6455_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7224__102 _8195_/CLK vssd1 vssd1 vccd1 vccd1 _8234_/CLK sky130_fd_sc_hd__inv_2
X_5406_ _5373_/Y _6973_/B _5548_/B _7079_/B vssd1 vssd1 vccd1 vccd1 _7598_/D sky130_fd_sc_hd__and4bb_1
X_6386_ _6386_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6388_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5162__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5337_ _6777_/A _5336_/B _5336_/Y hold228/X vssd1 vssd1 vccd1 vccd1 _5337_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_100_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7063__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8125_ _8125_/CLK _8125_/D vssd1 vssd1 vccd1 vccd1 _8125_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6111__C1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_595 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5268_ _6917_/A _5294_/A2 _5294_/B1 _5268_/B2 vssd1 vssd1 vccd1 vccd1 _5268_/X sky130_fd_sc_hd__a22o_1
X_8056_ _8056_/CLK _8056_/D vssd1 vssd1 vccd1 vccd1 _8056_/Q sky130_fd_sc_hd__dfxtp_1
X_4219_ _4219_/A _4219_/B vssd1 vssd1 vccd1 vccd1 _4219_/X sky130_fd_sc_hd__xor2_1
X_7007_ _7007_/A _7007_/B vssd1 vssd1 vccd1 vccd1 _7007_/X sky130_fd_sc_hd__and2_1
XANTENNA__4899__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5199_ _6927_/A _5221_/A2 _5221_/B1 hold821/X vssd1 vssd1 vccd1 vccd1 _5199_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4907__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5217__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6414__B1 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7909_ _8466_/CLK _7909_/D vssd1 vssd1 vccd1 vccd1 _7909_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3779__A1 _3778_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6717__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6423__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7136__14 _8328_/CLK vssd1 vssd1 vccd1 vccd1 _7513_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7254__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6248__A3 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _6842_/X vssd1 vssd1 vccd1 vccd1 _6845_/B sky130_fd_sc_hd__buf_12
XANTENNA__4817__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout291 _6667_/Y vssd1 vssd1 vccd1 vccd1 _6701_/A2 sky130_fd_sc_hd__buf_6
XANTENNA__5208__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3884__A_N _7283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6956__A1 _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6708__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6333__A _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5916__C1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6184__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4814__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4570_ _8140_/Q _7539_/Q _7411_/Q _7571_/Q _7362_/Q _4727_/S1 vssd1 vssd1 vccd1 vccd1
+ _4570_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_21_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold706 _5470_/X vssd1 vssd1 vccd1 vccd1 _7659_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold728 _5590_/X vssd1 vssd1 vccd1 vccd1 _7774_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold717 _7331_/Q vssd1 vssd1 vccd1 vccd1 _5428_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5144__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6240_ _3895_/B _6417_/A2 _6230_/Y _6239_/X _6347_/B1 vssd1 vssd1 vccd1 vccd1 _6240_/Y
+ sky130_fd_sc_hd__a221oi_2
Xhold739 _7789_/Q vssd1 vssd1 vccd1 vccd1 hold739/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6171_ _6155_/Y _6159_/B _6156_/Y vssd1 vssd1 vccd1 vccd1 _6177_/A sky130_fd_sc_hd__a21o_1
X_5122_ input23/X _5144_/A2 _5146_/B1 _5121_/X vssd1 vssd1 vccd1 vccd1 _7373_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1406 _8384_/Q vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1417 _8367_/Q vssd1 vssd1 vccd1 vccd1 _5022_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1428 hold1807/X vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__buf_1
Xhold1439 _7289_/Q vssd1 vssd1 vccd1 vccd1 _5134_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5053_ _7339_/Q _5468_/C vssd1 vssd1 vccd1 vccd1 _5053_/X sky130_fd_sc_hd__or2_1
XANTENNA__6508__A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ _4004_/A1 _4084_/A2 _4000_/X _4084_/B2 _4003_/X vssd1 vssd1 vccd1 vccd1 _4004_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_79_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5955_ _5955_/A _6008_/A vssd1 vssd1 vccd1 vccd1 _5955_/Y sky130_fd_sc_hd__nor2_2
XANTENNA_fanout240_A _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5886_ _5694_/Y _5881_/X _5882_/X _5885_/X vssd1 vssd1 vccd1 vccd1 _5886_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_48_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6243__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4906_ _8474_/Q _8406_/Q _8438_/Q _8312_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4906_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_118_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4837_ _4836_/X _4835_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7625_ _8030_/CLK _7625_/D vssd1 vssd1 vccd1 vccd1 _7625_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7220__98 _8388_/CLK vssd1 vssd1 vccd1 vccd1 _8230_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4805__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6897__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4768_ _6551_/A _4768_/B vssd1 vssd1 vccd1 vccd1 _8125_/D sky130_fd_sc_hd__and2_1
X_7556_ _8160_/CLK _7556_/D vssd1 vssd1 vccd1 vccd1 _7556_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7074__A _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4699_ _8481_/Q _8413_/Q _8445_/Q _8319_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4699_/X sky130_fd_sc_hd__mux4_1
X_7487_ _8475_/CLK _7487_/D vssd1 vssd1 vccd1 vccd1 _7487_/Q sky130_fd_sc_hd__dfxtp_1
X_3719_ _4770_/B _4071_/A2 _4071_/B1 _3717_/X _3718_/X vssd1 vssd1 vccd1 vccd1 _6318_/A
+ sky130_fd_sc_hd__o221a_4
X_6507_ _6524_/A _6507_/B vssd1 vssd1 vccd1 vccd1 _6507_/X sky130_fd_sc_hd__and2_1
X_6438_ _3770_/X _3771_/Y _3772_/X _6911_/A vssd1 vssd1 vccd1 vccd1 _6438_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1522_A _7354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8108_ _8108_/CLK _8108_/D vssd1 vssd1 vccd1 vccd1 _8108_/Q sky130_fd_sc_hd__dfxtp_2
X_6369_ _6370_/A _6370_/B vssd1 vssd1 vccd1 vccd1 _6369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3770__C_N _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
X_8039_ _8039_/CLK _8039_/D vssd1 vssd1 vccd1 vccd1 _8039_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6418__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__buf_1
XANTENNA__4637__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6650__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6137__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5041__B _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6938__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7060__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5610__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5992__A _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 _6442_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5126__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4547__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7051__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5601__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6063__A _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5740_ _6307_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5740_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_57_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_108_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8460_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4282__S _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6998__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7410_ _8175_/CLK _7410_/D vssd1 vssd1 vccd1 vccd1 _7410_/Q sky130_fd_sc_hd__dfxtp_1
X_5671_ _7022_/A hold77/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__and2_1
X_8390_ _8468_/CLK _8390_/D vssd1 vssd1 vccd1 vccd1 _8390_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5904__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4622_ _8470_/Q _8402_/Q _8434_/Q _8308_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4622_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_72_568 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5365__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3915__B2 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7341_ _8385_/CLK _7341_/D vssd1 vssd1 vccd1 vccd1 _7341_/Q sky130_fd_sc_hd__dfxtp_1
X_4553_ _4552_/X _4551_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4553_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold514 _5595_/X vssd1 vssd1 vccd1 vccd1 _7779_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5407__A _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold503 _7775_/Q vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold525 _7378_/Q vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _6550_/A _7903_/Q vssd1 vssd1 vccd1 vccd1 _8035_/D sky130_fd_sc_hd__and2_1
X_7272_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7272_/Y sky130_fd_sc_hd__inv_2
Xhold536 _5251_/X vssd1 vssd1 vccd1 vccd1 _7459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _8226_/Q vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 _5348_/X vssd1 vssd1 vccd1 vccd1 _7575_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ _6223_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6226_/B sky130_fd_sc_hd__xnor2_1
Xhold547 _7327_/Q vssd1 vssd1 vccd1 vccd1 _5424_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5841__S _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6154_ _6154_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6157_/B sky130_fd_sc_hd__xnor2_2
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6880__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1214 _6916_/X vssd1 vssd1 vccd1 vccd1 _8423_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1203 _8334_/Q vssd1 vssd1 vccd1 vccd1 _6794_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout190_A _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5105_ _5474_/A _5542_/C vssd1 vssd1 vccd1 vccd1 _5105_/X sky130_fd_sc_hd__or2_1
X_6085_ _5694_/Y _6084_/X _6083_/X vssd1 vssd1 vccd1 vccd1 _6085_/X sky130_fd_sc_hd__a21bo_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1225 _8406_/Q vssd1 vssd1 vccd1 vccd1 _6880_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6632__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1236 _6906_/X vssd1 vssd1 vccd1 vccd1 _8419_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 _8436_/Q vssd1 vssd1 vccd1 vccd1 _6942_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1258 _6626_/X vssd1 vssd1 vccd1 vccd1 _8177_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5036_ _5036_/A1 _5067_/S _5172_/B1 _5035_/X vssd1 vssd1 vccd1 vccd1 _7330_/D sky130_fd_sc_hd__o211a_1
Xhold1269 _8346_/Q vssd1 vssd1 vccd1 vccd1 _6818_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout455_A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6987_ _8528_/Z _6976_/Y _6986_/Y _5399_/A vssd1 vssd1 vccd1 vccd1 _6987_/X sky130_fd_sc_hd__a22o_1
XANTENNA__7069__A _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5938_ _5798_/X _5807_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5938_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5869_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5869_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6148__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7608_ _8369_/CLK _7608_/D vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5356__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3906__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7539_ _8419_/CLK _7539_/D vssd1 vssd1 vccd1 vccd1 _7539_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4221__A _4221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5108__B1 _5002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput67 _8113_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[12] sky130_fd_sc_hd__buf_12
XANTENNA__5751__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput89 _8104_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[3] sky130_fd_sc_hd__buf_12
Xoutput78 _8123_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[22] sky130_fd_sc_hd__buf_12
XFILLER_0_98_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1770 _6111_/X vssd1 vssd1 vccd1 vccd1 _7882_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5831__A1 _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1792 _8508_/Q vssd1 vssd1 vccd1 vccd1 _4029_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3842__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1781 _8489_/Q vssd1 vssd1 vccd1 vccd1 _3808_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7033__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5595__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5347__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4830__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6611__A _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5227__A _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output84_A _8129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5745__S1 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6862__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6614__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7131__9 _8464_/CLK vssd1 vssd1 vccd1 vccd1 _7508_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_89_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5897__A _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6910_ _6999_/A _6910_/A2 _6943_/B _6909_/X vssd1 vssd1 vccd1 vccd1 _6910_/X sky130_fd_sc_hd__a31o_1
X_7890_ _8503_/CLK _7890_/D vssd1 vssd1 vccd1 vccd1 _7890_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6841_ _7939_/Q _7940_/Q _6842_/C vssd1 vssd1 vccd1 vccd1 _6841_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8511_ _8513_/CLK _8511_/D vssd1 vssd1 vccd1 vccd1 _8511_/Q sky130_fd_sc_hd__dfxtp_1
X_3984_ _5946_/A _5943_/A vssd1 vssd1 vccd1 vccd1 _3985_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6772_ _6967_/A _6741_/B _6773_/B1 _6772_/B2 vssd1 vssd1 vccd1 vccd1 _6772_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5050__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5723_ _7596_/Q _5723_/B _5723_/C vssd1 vssd1 vccd1 vccd1 _5723_/X sky130_fd_sc_hd__or3_2
XANTENNA__4025__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6521__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5654_ _5667_/A _5654_/B vssd1 vssd1 vccd1 vccd1 _7834_/D sky130_fd_sc_hd__and2_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8442_ _8442_/CLK _8442_/D vssd1 vssd1 vccd1 vccd1 _8442_/Q sky130_fd_sc_hd__dfxtp_1
X_4605_ _8145_/Q _7544_/Q _7416_/Q _7576_/Q _4611_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4605_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_5_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8373_ _8373_/CLK _8373_/D _7267_/Y vssd1 vssd1 vccd1 vccd1 _8373_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5585_ _7010_/A _5585_/B vssd1 vssd1 vccd1 vccd1 _5585_/Y sky130_fd_sc_hd__nand2_1
Xhold300 _7469_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
X_7324_ _8368_/CLK _7324_/D vssd1 vssd1 vccd1 vccd1 _7324_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4010__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold311 _5459_/X vssd1 vssd1 vccd1 vccd1 _7648_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _5451_/X vssd1 vssd1 vccd1 vccd1 _7640_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _7405_/Q vssd1 vssd1 vccd1 vccd1 hold344/X sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ _4534_/X _4535_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4536_/X sky130_fd_sc_hd__mux2_1
Xhold322 _8518_/Q vssd1 vssd1 vccd1 vccd1 _5550_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4467_ _7010_/A _7920_/Q vssd1 vssd1 vccd1 vccd1 _8052_/D sky130_fd_sc_hd__and2_1
Xhold366 _8206_/Q vssd1 vssd1 vccd1 vccd1 hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _5253_/X vssd1 vssd1 vccd1 vccd1 _7461_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7255_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7255_/Y sky130_fd_sc_hd__inv_2
Xhold355 _5648_/X vssd1 vssd1 vccd1 vccd1 _7828_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 _5312_/X vssd1 vssd1 vccd1 vccd1 _7543_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6206_ _6206_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6209_/B sky130_fd_sc_hd__xnor2_1
Xhold388 _7389_/Q vssd1 vssd1 vccd1 vccd1 _5456_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4398_ _4398_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _4398_/Y sky130_fd_sc_hd__nor2_1
Xhold1000 _5589_/X vssd1 vssd1 vccd1 vccd1 _7773_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7071__B _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6137_ _6137_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6140_/B sky130_fd_sc_hd__xnor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 _8287_/Q vssd1 vssd1 vccd1 vccd1 _6732_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 _7411_/Q vssd1 vssd1 vccd1 vccd1 _5197_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1022 _6711_/X vssd1 vssd1 vccd1 vccd1 _8266_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1066 _6570_/X vssd1 vssd1 vccd1 vccd1 _8142_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _7015_/X vssd1 vssd1 vccd1 vccd1 _8473_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6068_ _5873_/X _5880_/X _6250_/S vssd1 vssd1 vccd1 vccd1 _6068_/X sky130_fd_sc_hd__mux2_1
Xhold1055 _7568_/Q vssd1 vssd1 vccd1 vccd1 _5341_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 _8420_/Q vssd1 vssd1 vccd1 vccd1 _6910_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 _7544_/Q vssd1 vssd1 vccd1 vccd1 _5313_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ _5419_/A _5453_/C vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1088 _7022_/X vssd1 vssd1 vccd1 vccd1 _8480_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4915__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_90_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6431__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5329__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7262__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_clk_A _7871_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4068__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output122_A _7287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_101_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5280__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5032__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4100__A_N _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_116_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4560__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5370_ _5470_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _5370_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4321_ _4315_/Y _4317_/B _4314_/Y vssd1 vssd1 vccd1 vccd1 _4325_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_120_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7040_ _7078_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7040_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4252_ _4242_/Y _4246_/B _4244_/B vssd1 vssd1 vccd1 vccd1 _4253_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_129_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5404__B _5404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4183_ _4183_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__6143__S1 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7942_ _8361_/CLK _7942_/D vssd1 vssd1 vccd1 vccd1 _7942_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6516__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4735__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5271__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7873_ _8469_/CLK _7873_/D vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6824_ _7028_/A _6824_/A2 _6838_/A3 _6823_/X vssd1 vssd1 vccd1 vccd1 _6824_/X sky130_fd_sc_hd__a31o_1
X_6755_ _6933_/A _6741_/B _6774_/B1 hold406/X vssd1 vssd1 vccd1 vccd1 _6755_/X sky130_fd_sc_hd__a22o_1
X_3967_ _3967_/A1 _4073_/A2 _6917_/A _4073_/B2 _3966_/X vssd1 vssd1 vccd1 vccd1 _3967_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6251__A _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5706_ _6175_/A _6191_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5706_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6771__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8029_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8425_ _8425_/CLK _8425_/D vssd1 vssd1 vccd1 vccd1 _8425_/Q sky130_fd_sc_hd__dfxtp_1
X_3898_ _3923_/B _7942_/Q vssd1 vssd1 vccd1 vccd1 _3898_/X sky130_fd_sc_hd__and2b_1
X_6686_ _6939_/A _6701_/A2 _6701_/B1 hold905/X vssd1 vssd1 vccd1 vccd1 _6686_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout418_A _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5637_ _6939_/A _5652_/A2 _5652_/B1 hold819/X vssd1 vssd1 vccd1 vccd1 _5637_/X sky130_fd_sc_hd__a22o_1
X_8356_ _8450_/CLK _8356_/D vssd1 vssd1 vccd1 vccd1 _8356_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5568_ _7027_/A _5568_/B vssd1 vssd1 vccd1 vccd1 _7757_/D sky130_fd_sc_hd__and2_1
XFILLER_0_130_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold130 _7609_/Q vssd1 vssd1 vccd1 vccd1 _5667_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _7611_/Q vssd1 vssd1 vccd1 vccd1 _5669_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4519_ _5389_/A _5374_/A _5409_/A vssd1 vssd1 vccd1 vccd1 _4519_/X sky130_fd_sc_hd__o21a_1
X_8287_ _8319_/CLK _8287_/D vssd1 vssd1 vccd1 vccd1 _8287_/Q sky130_fd_sc_hd__dfxtp_1
Xhold141 _6493_/X vssd1 vssd1 vccd1 vccd1 _7975_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7307_ _8091_/CLK _7307_/D _7117_/Y vssd1 vssd1 vccd1 vccd1 _7307_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_111_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6287__B2 _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7082__A _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3814__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 _6519_/X vssd1 vssd1 vccd1 vccd1 _8001_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _6461_/X vssd1 vssd1 vccd1 vccd1 _7943_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _7767_/Q vssd1 vssd1 vccd1 vccd1 _6518_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _7520_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7688_/D sky130_fd_sc_hd__and3_1
Xhold196 _7900_/Q vssd1 vssd1 vccd1 vccd1 _5000_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6826__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6039__A1 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_97_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _8373_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4645__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6426__A _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4696__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4123__A_N _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5014__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7257__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3785__A _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6762__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_21_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8402_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_64_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7181__59 _8010_/CLK vssd1 vssd1 vccd1 vccd1 _8061_/CLK sky130_fd_sc_hd__inv_2
X_7241__119 _8154_/CLK vssd1 vssd1 vccd1 vccd1 _8251_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6100__S _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _8020_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5253__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3679__B _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _8179_/Q _8211_/Q _8275_/Q _7783_/Q _4997_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4870_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3821_ _6350_/A _6352_/A vssd1 vssd1 vccd1 vccd1 _3823_/A sky130_fd_sc_hd__or2_1
XANTENNA__6202__A1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6753__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5961__A0 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6540_ _7018_/A _6540_/B vssd1 vssd1 vccd1 vccd1 _8022_/D sky130_fd_sc_hd__and2_1
XFILLER_0_70_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _8086_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3752_ _4067_/A_N _7955_/Q vssd1 vssd1 vccd1 vccd1 _3752_/X sky130_fd_sc_hd__and2b_1
X_6471_ _6534_/A hold11/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__and2_1
XFILLER_0_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _8092_/Q _3682_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3683_/X sky130_fd_sc_hd__mux2_1
X_8210_ _8466_/CLK _8210_/D vssd1 vssd1 vccd1 vccd1 _8210_/Q sky130_fd_sc_hd__dfxtp_1
X_5422_ _5422_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5422_/X sky130_fd_sc_hd__and3_1
XFILLER_0_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5713__A0 _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4611__S1 _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8141_ _8270_/CLK _8141_/D vssd1 vssd1 vccd1 vccd1 _8141_/Q sky130_fd_sc_hd__dfxtp_1
X_5353_ _6941_/A _5367_/A2 _5367_/B1 hold402/X vssd1 vssd1 vccd1 vccd1 _5353_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4304_ _4303_/Y _5046_/A1 _5503_/B vssd1 vssd1 vccd1 vccd1 _4392_/B sky130_fd_sc_hd__mux2_1
X_8072_ _8473_/CLK hold56/X vssd1 vssd1 vccd1 vccd1 _8072_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6808__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5284_ _6949_/A _5294_/A2 _5294_/B1 hold521/X vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__a22o_1
X_4235_ _8505_/Q _7642_/Q vssd1 vssd1 vccd1 vccd1 _4235_/Y sky130_fd_sc_hd__nor2_1
X_7023_ _7023_/A _7023_/B vssd1 vssd1 vccd1 vccd1 _7023_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_79_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _8030_/CLK sky130_fd_sc_hd__clkbuf_16
X_4166_ _8515_/Q _7632_/Q vssd1 vssd1 vccd1 vccd1 _4166_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4097_ _4097_/A _5963_/S vssd1 vssd1 vccd1 vccd1 _4097_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout368_A _7083_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5244__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4678__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7925_ _8457_/CLK _7925_/D vssd1 vssd1 vccd1 vccd1 _7925_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5795__A3 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7856_ _8020_/CLK _7856_/D vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
X_6807_ _6939_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6807_/X sky130_fd_sc_hd__and2_1
X_7787_ _8343_/CLK _7787_/D vssd1 vssd1 vccd1 vccd1 _7787_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7077__A _7077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4999_ _4998_/X _4995_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8261_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_135_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6738_ _6971_/A _6705_/B _6738_/B1 hold635/X vssd1 vssd1 vccd1 vccd1 _6738_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4850__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6669_ _6741_/A _6669_/B vssd1 vssd1 vccd1 vccd1 _6669_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_61_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8408_ _8476_/CLK _8408_/D vssd1 vssd1 vccd1 vccd1 _8408_/Q sky130_fd_sc_hd__dfxtp_1
X_8339_ _8339_/CLK _8339_/D vssd1 vssd1 vccd1 vccd1 _8339_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3730__A2 _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout440 _6539_/A vssd1 vssd1 vccd1 vccd1 _6524_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6680__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout451 _6494_/A vssd1 vssd1 vccd1 vccd1 _6498_/A sky130_fd_sc_hd__clkbuf_4
Xfanout462 input63/X vssd1 vssd1 vccd1 vccd1 _6347_/B1 sky130_fd_sc_hd__clkbuf_4
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6156__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6603__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6735__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3721__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6120__B1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6671__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4020_ _4020_/A _5974_/A vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5889__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8218_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5971_ _5971_/A _5971_/B vssd1 vssd1 vccd1 vccd1 _5974_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5857__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7710_ _8428_/CLK _7710_/D vssd1 vssd1 vccd1 vccd1 _7710_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5777__A3 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4922_ _4921_/X _4918_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8250_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_129_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7641_ _8370_/CLK _7641_/D vssd1 vssd1 vccd1 vccd1 _7641_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4853_ _8337_/Q _7813_/Q _7479_/Q _7447_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4853_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6726__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4784_ _8134_/Q _7533_/Q _7405_/Q _7565_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4784_/X sky130_fd_sc_hd__mux4_1
X_7572_ _8328_/CLK _7572_/D vssd1 vssd1 vccd1 vccd1 _7572_/Q sky130_fd_sc_hd__dfxtp_1
X_3804_ _7730_/Q _4070_/B vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__or2_1
X_6523_ _6706_/A _6523_/B vssd1 vssd1 vccd1 vccd1 _8005_/D sky130_fd_sc_hd__and2_1
XANTENNA__4832__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3735_ _4768_/B _4071_/A2 _4071_/B1 _6891_/A _3734_/X vssd1 vssd1 vccd1 vccd1 _6281_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_132_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6454_ _7006_/A _6454_/B vssd1 vssd1 vccd1 vccd1 _6454_/X sky130_fd_sc_hd__and2_1
X_3666_ _7834_/Q _3659_/Y _3660_/Y _7837_/Q vssd1 vssd1 vccd1 vccd1 _3666_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_113_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5405_ _7055_/A vssd1 vssd1 vccd1 vccd1 _5548_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6385_ _6371_/A _6373_/B _6369_/Y vssd1 vssd1 vccd1 vccd1 _6390_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5336_ _6706_/A _5336_/B vssd1 vssd1 vccd1 vccd1 _5336_/Y sky130_fd_sc_hd__nand2_2
X_8124_ _8124_/CLK _8124_/D vssd1 vssd1 vccd1 vccd1 _8124_/Q sky130_fd_sc_hd__dfxtp_1
X_5267_ _6849_/A _5263_/B _5263_/Y hold230/X vssd1 vssd1 vccd1 vccd1 _5267_/X sky130_fd_sc_hd__o22a_1
X_8055_ _8055_/CLK _8055_/D vssd1 vssd1 vccd1 vccd1 _8055_/Q sky130_fd_sc_hd__dfxtp_1
X_7006_ _7006_/A _7006_/B vssd1 vssd1 vccd1 vccd1 _7006_/X sky130_fd_sc_hd__and2_1
X_4218_ _4208_/Y _4212_/B _4210_/B vssd1 vssd1 vccd1 vccd1 _4218_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4899__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6662__A1 _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5198_ _6925_/A _5221_/A2 _5221_/B1 _5198_/B2 vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__a22o_1
X_4149_ _5732_/C _5690_/A _5723_/C _4153_/A _5723_/B vssd1 vssd1 vccd1 vccd1 _4149_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__5217__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7908_ _8029_/CLK _7908_/D vssd1 vssd1 vccd1 vccd1 _7908_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4520__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6178__A0 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6717__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7839_ _8361_/CLK _7839_/D vssd1 vssd1 vccd1 vccd1 _7839_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6423__B _6423_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5039__B _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3782__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4587__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7151__29 _8354_/CLK vssd1 vssd1 vccd1 vccd1 _7528_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_100_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7270__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout292 _6667_/Y vssd1 vssd1 vccd1 vccd1 _6669_/B sky130_fd_sc_hd__buf_8
Xfanout270 _3706_/Y vssd1 vssd1 vccd1 vccd1 _4084_/B2 sky130_fd_sc_hd__buf_8
Xfanout281 _6901_/B vssd1 vssd1 vccd1 vccd1 _6905_/B sky130_fd_sc_hd__buf_6
XFILLER_0_88_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5502__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5208__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3957__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4814__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3973__A _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7247__125 _8355_/CLK vssd1 vssd1 vccd1 vccd1 _8257_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold707 _8214_/Q vssd1 vssd1 vccd1 vccd1 hold707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold718 _5428_/X vssd1 vssd1 vccd1 vccd1 _7617_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 _8140_/Q vssd1 vssd1 vccd1 vccd1 hold729/X sky130_fd_sc_hd__dlygate4sd3_1
X_6170_ _6164_/X _6166_/X _6168_/Y _6169_/X _7026_/A vssd1 vssd1 vccd1 vccd1 _7885_/D
+ sky130_fd_sc_hd__o311a_1
X_5121_ _7031_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5121_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1407 _7646_/Q vssd1 vssd1 vccd1 vccd1 _4264_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6644__A1 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1418 _4227_/B vssd1 vssd1 vccd1 vccd1 _4505_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1429 _7304_/Q vssd1 vssd1 vccd1 vccd1 _5164_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5052_ _5052_/A1 _5067_/S _5166_/B1 _5051_/X vssd1 vssd1 vccd1 vccd1 _7338_/D sky130_fd_sc_hd__o211a_1
X_4003_ _4754_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _4003_/X sky130_fd_sc_hd__and2_1
XANTENNA__5412__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4743__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5080__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5954_ _5957_/A _5953_/Y _6129_/B vssd1 vssd1 vccd1 vccd1 _5954_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6524__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5885_ _6250_/S _5739_/Y _5878_/X _5884_/X vssd1 vssd1 vccd1 vccd1 _5885_/X sky130_fd_sc_hd__a31o_1
X_4905_ _8184_/Q _8216_/Q _8280_/Q _7788_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4905_/X sky130_fd_sc_hd__mux4_1
X_4836_ _8464_/Q _8396_/Q _8428_/Q _8302_/Q _5475_/A _7358_/Q vssd1 vssd1 vccd1 vccd1
+ _4836_/X sky130_fd_sc_hd__mux4_1
XANTENNA_fanout233_A _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7624_ _8033_/CLK _7624_/D vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4805__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7555_ _8486_/CLK _7555_/D vssd1 vssd1 vccd1 vccd1 _7555_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6580__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4767_ _6545_/A _4767_/B vssd1 vssd1 vccd1 vccd1 _8124_/D sky130_fd_sc_hd__and2_1
X_6506_ _6550_/A hold23/X vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__and2_1
XFILLER_0_31_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4698_ _8191_/Q _8223_/Q _8287_/Q _7795_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4698_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout400_A _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3718_ _3718_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3718_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7486_ _8346_/CLK _7486_/D vssd1 vssd1 vccd1 vccd1 _7486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3649_ _3649_/A vssd1 vssd1 vccd1 vccd1 _7052_/A sky130_fd_sc_hd__clkinv_4
X_6437_ _7017_/A _6437_/B vssd1 vssd1 vccd1 vccd1 _7919_/D sky130_fd_sc_hd__and2_1
XANTENNA__4569__S0 _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6368_ _6370_/A _6370_/B vssd1 vssd1 vccd1 vccd1 _6371_/A sky130_fd_sc_hd__nand2_1
X_8107_ _8107_/CLK _8107_/D vssd1 vssd1 vccd1 vccd1 _8107_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4918__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5319_ _6945_/A _5299_/B _5331_/B1 hold627/X vssd1 vssd1 vccd1 vccd1 _5319_/X sky130_fd_sc_hd__a22o_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7090__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6299_ _6299_/A _6299_/B vssd1 vssd1 vccd1 vccd1 _6301_/A sky130_fd_sc_hd__nor2_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
X_8038_ _8038_/CLK _8038_/D vssd1 vssd1 vccd1 vccd1 _8038_/Q sky130_fd_sc_hd__dfxtp_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__buf_1
XANTENNA__4741__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7060__A1 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6434__A _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5610__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6571__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7265__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_9 _6449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6874__A1 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6609__A _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output152_A _8038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6626__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4980__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3968__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5062__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5601__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5670_ _6534_/A hold49/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__and2_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6011__C1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4621_ _8180_/Q _8212_/Q _8276_/Q _7784_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4621_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_57_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5365__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6562__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3915__A2 _3669_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7340_ _8494_/CLK _7340_/D vssd1 vssd1 vccd1 vccd1 _7340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4552_ _8460_/Q _8392_/Q _8424_/Q _8298_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4552_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_123_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold504 _5591_/X vssd1 vssd1 vccd1 vccd1 _7775_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold526 _5445_/X vssd1 vssd1 vccd1 vccd1 _7634_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _7023_/A _7904_/Q vssd1 vssd1 vccd1 vccd1 _8036_/D sky130_fd_sc_hd__and2_1
XFILLER_0_13_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold515 _7587_/Q vssd1 vssd1 vccd1 vccd1 hold515/X sky130_fd_sc_hd__dlygate4sd3_1
X_7271_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7271_/Y sky130_fd_sc_hd__inv_2
X_6222_ _6212_/Y _6218_/X _6219_/X _6220_/X _6221_/Y vssd1 vssd1 vccd1 vccd1 _7888_/D
+ sky130_fd_sc_hd__o41a_1
Xhold548 _5424_/X vssd1 vssd1 vccd1 vccd1 _7613_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold537 _8285_/Q vssd1 vssd1 vccd1 vccd1 hold537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _7590_/Q vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_9_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6153_ _6147_/X _6149_/X _6151_/Y _6152_/Y vssd1 vssd1 vccd1 vccd1 _6153_/X sky130_fd_sc_hd__o31a_1
XANTENNA__6519__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _6794_/X vssd1 vssd1 vccd1 vccd1 _8334_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6084_ _5897_/B _5909_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6084_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ input13/X _5099_/B _5002_/X _5103_/X vssd1 vssd1 vccd1 vccd1 _7364_/D sky130_fd_sc_hd__o211a_1
Xhold1215 _8378_/Q vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 _6942_/X vssd1 vssd1 vccd1 vccd1 _8436_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 _6880_/X vssd1 vssd1 vccd1 vccd1 _8406_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _8412_/Q vssd1 vssd1 vccd1 vccd1 _6892_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4723__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5035_ _5427_/A _5463_/C vssd1 vssd1 vccd1 vccd1 _5035_/X sky130_fd_sc_hd__or2_1
Xhold1259 _8409_/Q vssd1 vssd1 vccd1 vccd1 _6886_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3878__A _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout448_A _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6986_ _7354_/Q _6986_/B vssd1 vssd1 vccd1 vccd1 _6986_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout350_A _5732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7069__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5937_ _5795_/X _5797_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5937_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7607_ _8365_/CLK _7607_/D vssd1 vssd1 vccd1 vccd1 _7607_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5868_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5871_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4819_ _8139_/Q _7538_/Q _7410_/Q _7570_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4819_/X sky130_fd_sc_hd__mux4_1
X_5799_ _5797_/X _5798_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5799_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3817__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5356__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7538_ _8175_/CLK _7538_/D vssd1 vssd1 vccd1 vccd1 _7538_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3906__A2 _3904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1465_A _7312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7469_ _7805_/CLK _7469_/D vssd1 vssd1 vccd1 vccd1 _7469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_120_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1632_A _4039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6856__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput68 _8114_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[13] sky130_fd_sc_hd__buf_12
XANTENNA__6429__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4648__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput79 _8124_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[23] sky130_fd_sc_hd__buf_12
XANTENNA__4962__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6608__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1771 _7721_/Q vssd1 vssd1 vccd1 vccd1 _3887_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1760 _7725_/Q vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5831__A2 _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5292__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1793 _4032_/B vssd1 vssd1 vccd1 vccd1 _6050_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3842__A1 _4775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3842__B2 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1782 _3811_/B vssd1 vssd1 vccd1 vccd1 _6400_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_2_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5044__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5595__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5347__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6611__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output77_A _8122_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4705__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5283__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6840_ _7029_/A _6840_/A2 _6779_/B _6839_/X vssd1 vssd1 vccd1 vccd1 _6840_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_77_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5586__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6771_ _6965_/A _6773_/A2 _6773_/B1 hold799/X vssd1 vssd1 vccd1 vccd1 _6771_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_119_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8510_ _8510_/CLK _8510_/D vssd1 vssd1 vccd1 vccd1 _8510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3983_ _5946_/A _5943_/A vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__or2_1
X_5722_ _5732_/C _5723_/B _5723_/C vssd1 vssd1 vccd1 vccd1 _6406_/B sky130_fd_sc_hd__nor3_4
XFILLER_0_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7187__65 _8010_/CLK vssd1 vssd1 vccd1 vccd1 _8099_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5338__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8441_ _8477_/CLK _8441_/D vssd1 vssd1 vccd1 vccd1 _8441_/Q sky130_fd_sc_hd__dfxtp_1
X_5653_ _6971_/A _5620_/B _5653_/B1 hold671/X vssd1 vssd1 vccd1 vccd1 _5653_/X sky130_fd_sc_hd__a22o_1
X_4604_ _8338_/Q _7814_/Q _7480_/Q _7448_/Q _4611_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4604_/X sky130_fd_sc_hd__mux4_1
X_5584_ _6741_/A _5584_/B vssd1 vssd1 vccd1 vccd1 _5584_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8372_ _8485_/CLK _8372_/D _7266_/Y vssd1 vssd1 vccd1 vccd1 _8372_/Q sky130_fd_sc_hd__dfrtp_1
Xhold301 _5265_/X vssd1 vssd1 vccd1 vccd1 _7469_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7323_ _8368_/CLK _7323_/D vssd1 vssd1 vccd1 vccd1 _7323_/Q sky130_fd_sc_hd__dfxtp_1
X_4535_ _8135_/Q _7534_/Q _7406_/Q _7566_/Q _4611_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4535_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold312 _7770_/Q vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _7436_/Q vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _5550_/X vssd1 vssd1 vccd1 vccd1 _7739_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6838__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4466_ _6999_/A _7921_/Q vssd1 vssd1 vccd1 vccd1 _8053_/D sky130_fd_sc_hd__and2_1
Xhold345 _5191_/X vssd1 vssd1 vccd1 vccd1 _7405_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _6679_/X vssd1 vssd1 vccd1 vccd1 _8206_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 _7382_/Q vssd1 vssd1 vccd1 vccd1 _5449_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7254_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7254_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_41_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold378 _8314_/Q vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
X_6205_ _6190_/Y _6194_/B _6192_/B vssd1 vssd1 vccd1 vccd1 _6211_/A sky130_fd_sc_hd__a21o_1
Xhold389 _5456_/X vssd1 vssd1 vccd1 vccd1 _7645_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4944__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4397_ _4401_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout398_A _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6136_ _6114_/Y _6119_/B _6116_/B vssd1 vssd1 vccd1 vccd1 _6142_/A sky130_fd_sc_hd__a21o_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1001 _8275_/Q vssd1 vssd1 vccd1 vccd1 _6720_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1023 _8477_/Q vssd1 vssd1 vccd1 vccd1 _7019_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1012 _6732_/X vssd1 vssd1 vccd1 vccd1 _8287_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5274__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6067_ _6250_/S _5878_/X _6066_/X _5740_/B vssd1 vssd1 vccd1 vccd1 _6067_/X sky130_fd_sc_hd__o211a_1
Xhold1034 _5197_/X vssd1 vssd1 vccd1 vccd1 _7411_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 _7465_/Q vssd1 vssd1 vccd1 vccd1 _5257_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 _5341_/X vssd1 vssd1 vccd1 vccd1 _7568_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 _8324_/Q vssd1 vssd1 vccd1 vccd1 _6773_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 _8390_/Q vssd1 vssd1 vccd1 vccd1 _6848_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1078 _5313_/X vssd1 vssd1 vccd1 vccd1 _7544_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5018_ _5018_/A1 _4425_/B _5146_/B1 _5017_/X vssd1 vssd1 vccd1 vccd1 _7321_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5026__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6774__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6969_ _6969_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6969_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5329__A1 _3814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5047__B _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold890 _5641_/X vssd1 vssd1 vccd1 vccd1 _7821_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5063__A _5404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5510__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1590 _4329_/Y vssd1 vssd1 vccd1 vccd1 _4330_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output115_A _7310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6765__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4841__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6780__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4320_ _4390_/A _4390_/B _4327_/C vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__and3_1
XFILLER_0_120_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4926__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4251_ _4249_/Y _4251_/B vssd1 vssd1 vccd1 vccd1 _4251_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_129_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4182_ _4180_/Y _4182_/B vssd1 vssd1 vccd1 vccd1 _4183_/B sky130_fd_sc_hd__and2b_1
XANTENNA__4059__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5256__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7941_ _8364_/CLK hold76/X vssd1 vssd1 vccd1 vccd1 _7941_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5420__B _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7872_ _8504_/CLK _7872_/D vssd1 vssd1 vccd1 vccd1 _7872_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5008__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4036__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6756__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6823_ _6955_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6823_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6532__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6220__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6754_ _6931_/A _6773_/A2 _6773_/B1 hold575/X vssd1 vssd1 vccd1 vccd1 _6754_/X sky130_fd_sc_hd__a22o_1
X_3966_ _4748_/B _3966_/B vssd1 vssd1 vccd1 vccd1 _3966_/X sky130_fd_sc_hd__and2_1
XFILLER_0_128_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6685_ _6937_/A _6669_/B _6702_/B1 hold459/X vssd1 vssd1 vccd1 vccd1 _6685_/X sky130_fd_sc_hd__a22o_1
X_5705_ _6140_/A _6157_/A _5744_/S vssd1 vssd1 vccd1 vccd1 _5705_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_18_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3990__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5636_ _6937_/A _5620_/B _5653_/B1 hold565/X vssd1 vssd1 vccd1 vccd1 _5636_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3897_ _3897_/A _3897_/B _3897_/C _3897_/D vssd1 vssd1 vccd1 vccd1 _4092_/A sky130_fd_sc_hd__or4_2
X_8424_ _8483_/CLK _8424_/D vssd1 vssd1 vccd1 vccd1 _8424_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout313_A _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5567_ _6524_/A _5567_/B vssd1 vssd1 vccd1 vccd1 _7756_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8355_ _8355_/CLK _8355_/D vssd1 vssd1 vccd1 vccd1 _8355_/Q sky130_fd_sc_hd__dfxtp_1
Xhold131 _5667_/X vssd1 vssd1 vccd1 vccd1 _7847_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _5669_/X vssd1 vssd1 vccd1 vccd1 _7849_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _7746_/Q vssd1 vssd1 vccd1 vccd1 _6497_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _6553_/A _5408_/B _5391_/A vssd1 vssd1 vccd1 vccd1 _5374_/A sky130_fd_sc_hd__or3b_4
X_5498_ _7519_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7687_/D sky130_fd_sc_hd__and3_1
Xhold142 _7627_/Q vssd1 vssd1 vccd1 vccd1 _5685_/B sky130_fd_sc_hd__dlygate4sd3_1
X_8286_ _8460_/CLK _8286_/D vssd1 vssd1 vccd1 vccd1 _8286_/Q sky130_fd_sc_hd__dfxtp_1
X_7306_ _8382_/CLK _7306_/D _7116_/Y vssd1 vssd1 vccd1 vccd1 _7306_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3742__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold164 _7749_/Q vssd1 vssd1 vccd1 vccd1 _6500_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4449_/A _4449_/B vssd1 vssd1 vccd1 vccd1 _4449_/X sky130_fd_sc_hd__or2_1
Xhold186 _7629_/Q vssd1 vssd1 vccd1 vccd1 _5687_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 _6518_/X vssd1 vssd1 vccd1 vccd1 _8000_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4917__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 _5000_/X vssd1 vssd1 vccd1 vccd1 _7282_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6039__A2 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7099_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7099_/Y sky130_fd_sc_hd__inv_2
X_6119_ _6119_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6119_/X sky130_fd_sc_hd__or2_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6426__B _6426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6747__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6442__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3981__B1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__7273__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5505__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5238__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6617__A _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3740__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6738__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3820_ _4772_/B _4071_/A2 _4071_/B1 _6965_/A _3819_/X vssd1 vssd1 vccd1 vccd1 _6352_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6352__A _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4571__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3751_ _3736_/Y _3737_/X _3750_/X vssd1 vssd1 vccd1 vccd1 _3897_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_40_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7157__35 _8480_/CLK vssd1 vssd1 vccd1 vccd1 _8037_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5961__A1 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3972__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6470_ _6548_/A _6470_/B vssd1 vssd1 vccd1 vccd1 _6470_/X sky130_fd_sc_hd__and2_1
X_3682_ _7996_/Q _4068_/A2 _4068_/B1 _8028_/Q _3680_/X vssd1 vssd1 vccd1 vccd1 _3682_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5421_ _5421_/A _5453_/B _5451_/C vssd1 vssd1 vccd1 vccd1 _5421_/X sky130_fd_sc_hd__and3_1
XANTENNA__5713__A1 _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8140_ _8173_/CLK _8140_/D vssd1 vssd1 vccd1 vccd1 _8140_/Q sky130_fd_sc_hd__dfxtp_1
X_5352_ _6939_/A _5367_/A2 _5367_/B1 hold561/X vssd1 vssd1 vccd1 vccd1 _5352_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5415__B _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8071_ _8071_/CLK _8105_/D vssd1 vssd1 vccd1 vccd1 _8071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4303_ _5572_/B vssd1 vssd1 vccd1 vccd1 _4303_/Y sky130_fd_sc_hd__inv_2
X_5283_ _6947_/A _5294_/A2 _5294_/B1 hold641/X vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__a22o_1
X_7022_ _7022_/A _7022_/B vssd1 vssd1 vccd1 vccd1 _7022_/X sky130_fd_sc_hd__and2_1
X_4234_ _4425_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4234_/Y sky130_fd_sc_hd__nand2_1
X_4165_ _8516_/Q _4156_/B _4159_/B vssd1 vssd1 vccd1 vccd1 _4165_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6527__A _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4096_ _3949_/Y _4093_/Y _4095_/A _3922_/B _4097_/A vssd1 vssd1 vccd1 vccd1 _4096_/Y
+ sky130_fd_sc_hd__o2111ai_1
XANTENNA_fanout263_A _5226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7924_ _8471_/CLK _7924_/D vssd1 vssd1 vccd1 vccd1 _7924_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6729__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7855_ _8504_/CLK _7855_/D vssd1 vssd1 vccd1 vccd1 _7855_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_42_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6806_ _7019_/A _6806_/A2 _6779_/B _6805_/X vssd1 vssd1 vccd1 vccd1 _6806_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6262__A _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout430_A _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4998_ _4997_/X _4996_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4998_/X sky130_fd_sc_hd__mux2_1
X_7786_ _8477_/CLK _7786_/D vssd1 vssd1 vccd1 vccd1 _7786_/Q sky130_fd_sc_hd__dfxtp_1
X_3949_ _5765_/A vssd1 vssd1 vccd1 vccd1 _3949_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6737_ _6969_/A _6737_/A2 _6737_/B1 hold755/X vssd1 vssd1 vccd1 vccd1 _6737_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6668_ _6842_/C _6704_/B vssd1 vssd1 vccd1 vccd1 _6670_/B sky130_fd_sc_hd__or2_1
XFILLER_0_116_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_57_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5619_ _6776_/A _6842_/C vssd1 vssd1 vccd1 vccd1 _5621_/B sky130_fd_sc_hd__or2_1
XFILLER_0_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6599_ _6595_/Y _6598_/X _5382_/X vssd1 vssd1 vccd1 vccd1 _6600_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8407_ _8475_/CLK _8407_/D vssd1 vssd1 vccd1 vccd1 _8407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8338_ _8338_/CLK _8338_/D vssd1 vssd1 vccd1 vccd1 _8338_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5180__A2 _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_100_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8269_ _8478_/CLK _8269_/D vssd1 vssd1 vccd1 vccd1 _8269_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout441 _6539_/A vssd1 vssd1 vccd1 vccd1 _6520_/A sky130_fd_sc_hd__clkbuf_4
Xfanout430 _6434_/A vssd1 vssd1 vccd1 vccd1 _7025_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6680__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout452 _4775_/A vssd1 vssd1 vccd1 vccd1 _6494_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_115_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6437__A _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout463 _7281_/A vssd1 vssd1 vccd1 vccd1 _7273_/A sky130_fd_sc_hd__buf_8
XANTENNA__6417__C1 _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7268__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6408__C1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5857__S1 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5970_ _5945_/Y _5949_/B _5947_/B vssd1 vssd1 vccd1 vccd1 _5976_/A sky130_fd_sc_hd__a21o_1
XANTENNA__5631__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4921_ _4920_/X _4919_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__mux2_1
X_7640_ _8368_/CLK _7640_/D vssd1 vssd1 vccd1 vccd1 _7640_/Q sky130_fd_sc_hd__dfxtp_1
X_4852_ _4851_/X _4848_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8240_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3803_ _8097_/Q _3802_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3803_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4783_ _8327_/Q _7803_/Q _7469_/Q _7437_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4783_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5934__A1 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7571_ _8354_/CLK _7571_/D vssd1 vssd1 vccd1 vccd1 _7571_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6522_ _7008_/A _6522_/B vssd1 vssd1 vccd1 vccd1 _8004_/D sky130_fd_sc_hd__and2_1
XFILLER_0_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3734_ _7724_/Q _4070_/B vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__or2_1
X_3665_ _7837_/Q _3660_/Y _3661_/Y _7836_/Q vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__o22a_1
X_6453_ _7018_/A _6453_/B vssd1 vssd1 vccd1 vccd1 _7935_/D sky130_fd_sc_hd__and2_1
X_5404_ _5404_/A _5404_/B _5404_/C vssd1 vssd1 vccd1 vccd1 _7055_/A sky130_fd_sc_hd__and3_2
XANTENNA__5698__A0 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6384_ _6378_/Y _6381_/X _6382_/Y _6383_/Y vssd1 vssd1 vccd1 vccd1 _7897_/D sky130_fd_sc_hd__o31a_1
X_8123_ _8123_/CLK _8123_/D vssd1 vssd1 vccd1 vccd1 _8123_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_3_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5162__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5335_ _6741_/A _5335_/B vssd1 vssd1 vccd1 vccd1 _5335_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__5860__S _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5266_ _6847_/A _5262_/B _5295_/B1 _5266_/B2 vssd1 vssd1 vccd1 vccd1 _5266_/X sky130_fd_sc_hd__a22o_1
X_8054_ _8054_/CLK _8054_/D vssd1 vssd1 vccd1 vccd1 _8054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4217_ _4215_/Y _4217_/B vssd1 vssd1 vccd1 vccd1 _4219_/A sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout380_A _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7005_ _7005_/A _7005_/B vssd1 vssd1 vccd1 vccd1 _7005_/X sky130_fd_sc_hd__and2_1
X_5197_ _6923_/A _5188_/B _5220_/B1 _5197_/B2 vssd1 vssd1 vccd1 vccd1 _5197_/X sky130_fd_sc_hd__a22o_1
X_4148_ _8453_/Q _4148_/B vssd1 vssd1 vccd1 vccd1 _5723_/C sky130_fd_sc_hd__or2_2
X_4079_ _7984_/Q _4079_/A2 _4079_/B1 _8016_/Q _4078_/X vssd1 vssd1 vccd1 vccd1 _4079_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6414__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7907_ _7907_/CLK _7907_/D vssd1 vssd1 vccd1 vccd1 _7907_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4520__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7088__A _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6178__A1 _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7838_ _8364_/CLK _7838_/D vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7769_ _8500_/CLK _7769_/D vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5336__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4587__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4386__S _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 _6841_/Y vssd1 vssd1 vccd1 vccd1 _6901_/B sky130_fd_sc_hd__buf_8
Xfanout260 _5299_/Y vssd1 vssd1 vccd1 vccd1 _5332_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout271 _4081_/B vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__buf_4
XFILLER_0_88_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout293 _6605_/B vssd1 vssd1 vccd1 vccd1 _6666_/A3 sky130_fd_sc_hd__buf_8
XANTENNA__5502__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6956__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5613__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6169__A1 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4415__A _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3973__B _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold719 _8466_/Q vssd1 vssd1 vccd1 vccd1 _7008_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold708 _6687_/X vssd1 vssd1 vccd1 vccd1 _8214_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5144__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5120_ input22/X _5144_/A2 _5146_/B1 _5119_/X vssd1 vssd1 vccd1 vccd1 _7372_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4296__S _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5051_ _5435_/A _5463_/C vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__or2_1
X_4002_ _4754_/B _3676_/A _4082_/B1 _6929_/A _4001_/X vssd1 vssd1 vccd1 vccd1 _6016_/A
+ sky130_fd_sc_hd__o221a_4
Xhold1419 _8359_/Q vssd1 vssd1 vccd1 vccd1 _4448_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1408 _4264_/Y vssd1 vssd1 vccd1 vccd1 _4265_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6805__A _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5604__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5080__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ _6270_/A _5953_/B vssd1 vssd1 vccd1 vccd1 _5953_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5884_ _3973_/X _3974_/Y _6105_/A2 _5883_/X vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_5_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4904_ _4902_/X _4903_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__mux2_1
X_4835_ _8174_/Q _8206_/Q _8270_/Q _7778_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4835_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_90_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7623_ _8385_/CLK hold99/X vssd1 vssd1 vccd1 vccd1 _7623_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4766_ _7005_/A _4766_/B vssd1 vssd1 vccd1 vccd1 _8123_/D sky130_fd_sc_hd__and2_1
X_7554_ _8354_/CLK _7554_/D vssd1 vssd1 vccd1 vccd1 _7554_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6540__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6580__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout226_A _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3717_ _8093_/Q _3716_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3717_/X sky130_fd_sc_hd__mux2_2
X_6505_ _6545_/A hold57/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__and2_1
XFILLER_0_132_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7485_ _8461_/CLK _7485_/D vssd1 vssd1 vccd1 vccd1 _7485_/Q sky130_fd_sc_hd__dfxtp_1
X_4697_ _4695_/X _4696_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3648_ _5473_/A vssd1 vssd1 vccd1 vccd1 _3648_/Y sky130_fd_sc_hd__inv_2
XANTENNA__7074__C _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4569__S1 _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6436_ _7018_/A _6436_/B vssd1 vssd1 vccd1 vccd1 _7918_/D sky130_fd_sc_hd__and2_1
XFILLER_0_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6367_ _6367_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6370_/B sky130_fd_sc_hd__xnor2_1
X_5318_ _6877_/A _5332_/A2 _5332_/B1 hold995/X vssd1 vssd1 vccd1 vccd1 _5318_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_101_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8106_ _8106_/CLK hold56/A vssd1 vssd1 vccd1 vccd1 _8106_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_87_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
X_6298_ _6298_/A _6298_/B vssd1 vssd1 vccd1 vccd1 _6299_/B sky130_fd_sc_hd__nor2_1
X_5249_ _6951_/A _5226_/B _5259_/B1 hold429/X vssd1 vssd1 vccd1 vccd1 _5249_/X sky130_fd_sc_hd__a22o_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
X_8037_ _8037_/CLK _8037_/D vssd1 vssd1 vccd1 vccd1 _8037_/Q sky130_fd_sc_hd__dfxtp_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4741__S1 _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6938__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4009__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6434__B _6434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4235__A _8505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6450__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7211__89 _8090_/CLK vssd1 vssd1 vccd1 vccd1 _8124_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6571__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5126__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7281__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6609__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5513__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4980__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4844__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6625__A _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7284__RESET_B _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3984__A _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4620_ _4618_/X _4619_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4620_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6562__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5365__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4551_ _8170_/Q _8202_/Q _8266_/Q _7774_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4551_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_123_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold505 _7419_/Q vssd1 vssd1 vccd1 vccd1 hold505/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4482_ _7022_/A _7905_/Q vssd1 vssd1 vccd1 vccd1 _8037_/D sky130_fd_sc_hd__and2_1
Xhold527 _8221_/Q vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _5360_/X vssd1 vssd1 vccd1 vccd1 _7587_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7270_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7270_/Y sky130_fd_sc_hd__inv_2
X_6221_ _3872_/B _6417_/A2 _6347_/B1 vssd1 vssd1 vccd1 vccd1 _6221_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold538 _6730_/X vssd1 vssd1 vccd1 vccd1 _8285_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 _7462_/Q vssd1 vssd1 vccd1 vccd1 hold549/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6152_ _3764_/B _6417_/A2 _7267_/A vssd1 vssd1 vccd1 vccd1 _6152_/Y sky130_fd_sc_hd__a21oi_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5103_ _5103_/A _5538_/C vssd1 vssd1 vccd1 vccd1 _5103_/X sky130_fd_sc_hd__or2_1
XANTENNA__5423__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6083_ _6083_/A _6083_/B vssd1 vssd1 vccd1 vccd1 _6083_/X sky130_fd_sc_hd__or2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1205 _8424_/Q vssd1 vssd1 vccd1 vccd1 _6918_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 _5044_/X vssd1 vssd1 vccd1 vccd1 _7334_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _8396_/Q vssd1 vssd1 vccd1 vccd1 _6860_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5825__B1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5034_/A1 _4416_/B _5166_/B1 _5033_/X vssd1 vssd1 vccd1 vccd1 _7329_/D sky130_fd_sc_hd__o211a_1
Xhold1238 _6892_/X vssd1 vssd1 vccd1 vccd1 _8412_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4723__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1227 _8442_/Q vssd1 vssd1 vccd1 vccd1 _6954_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout176_A _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3878__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6985_ _7090_/A _6985_/B vssd1 vssd1 vccd1 vccd1 _8453_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_73_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5936_ _6250_/S _5936_/B vssd1 vssd1 vccd1 vccd1 _5936_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7606_ _8365_/CLK _7606_/D vssd1 vssd1 vccd1 vccd1 _7606_/Q sky130_fd_sc_hd__dfxtp_1
X_5867_ _6198_/S _5971_/B vssd1 vssd1 vccd1 vccd1 _5870_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__6270__A _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4818_ _8332_/Q _7808_/Q _7474_/Q _7442_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4818_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5798_ _5701_/X _5705_/X _5859_/S vssd1 vssd1 vccd1 vccd1 _5798_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5356__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7537_ _8461_/CLK _7537_/D vssd1 vssd1 vccd1 vccd1 _7537_/Q sky130_fd_sc_hd__dfxtp_1
X_4749_ _7015_/A hold55/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__and2_1
XFILLER_0_7_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7468_ _7805_/CLK _7468_/D vssd1 vssd1 vccd1 vccd1 _7468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5108__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4929__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6419_ _6534_/A _6419_/B vssd1 vssd1 vccd1 vccd1 _6419_/X sky130_fd_sc_hd__and2_1
XFILLER_0_98_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7399_ _8501_/CLK _7399_/D vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
Xoutput69 _8115_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[14] sky130_fd_sc_hd__buf_12
XANTENNA__4962__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6608__A2 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5816__B1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1750 _6417_/Y vssd1 vssd1 vccd1 vccd1 _7899_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1761 _8500_/Q vssd1 vssd1 vccd1 vccd1 _3796_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5292__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6445__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1794 _7902_/Q vssd1 vssd1 vccd1 vccd1 _6454_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1783 _8514_/Q vssd1 vssd1 vccd1 vccd1 _3993_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3842__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1772 _6226_/A vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5831__A3 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5595__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6792__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7276__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5347__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4412__B _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4650__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5283__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4705__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3982_ _3982_/A0 _3981_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _5943_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_69_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6770_ _6963_/A _6773_/A2 _6774_/B1 hold795/X vssd1 vssd1 vccd1 vccd1 _6770_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_134_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5721_ _5721_/A vssd1 vssd1 vccd1 vccd1 _5721_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5652_ _6969_/A _5652_/A2 _5652_/B1 hold709/X vssd1 vssd1 vccd1 vccd1 _5652_/X sky130_fd_sc_hd__a22o_1
X_8440_ _8440_/CLK _8440_/D vssd1 vssd1 vccd1 vccd1 _8440_/Q sky130_fd_sc_hd__dfxtp_1
X_5583_ _6740_/C _6704_/B vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__or2_2
XFILLER_0_115_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5418__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5743__C1 _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4603_ _4602_/X _4599_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7511_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_4_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8371_ _8485_/CLK _8371_/D _7265_/Y vssd1 vssd1 vccd1 vccd1 _8371_/Q sky130_fd_sc_hd__dfrtp_1
X_4534_ _8328_/Q _7804_/Q _7470_/Q _7438_/Q _4611_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4534_/X sky130_fd_sc_hd__mux4_1
X_7322_ _8369_/CLK _7322_/D vssd1 vssd1 vccd1 vccd1 _7322_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4010__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold302 _7397_/Q vssd1 vssd1 vccd1 vccd1 _5464_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _5586_/X vssd1 vssd1 vccd1 vccd1 _7770_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _5228_/X vssd1 vssd1 vccd1 vccd1 _7436_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold324 _7395_/Q vssd1 vssd1 vccd1 vccd1 _5462_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold368 _7326_/Q vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _5449_/X vssd1 vssd1 vccd1 vccd1 _7638_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7253_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7253_/Y sky130_fd_sc_hd__inv_2
X_4465_ _7017_/A _7922_/Q vssd1 vssd1 vccd1 vccd1 _8054_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold346 _7329_/Q vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ _6204_/A1 _6417_/A2 _6203_/X _6347_/B1 vssd1 vssd1 vccd1 vccd1 _6204_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_7_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4944__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold379 _6763_/X vssd1 vssd1 vccd1 vccd1 _8314_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4396_ _4392_/A _5462_/C _4395_/X _4394_/X vssd1 vssd1 vccd1 vccd1 _8378_/D sky130_fd_sc_hd__a31o_1
XANTENNA_fanout293_A _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6135_ _6120_/Y _6125_/X _6133_/X _6134_/Y vssd1 vssd1 vccd1 vccd1 _7883_/D sky130_fd_sc_hd__o31a_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _6720_/X vssd1 vssd1 vccd1 vccd1 _8275_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1024 _7019_/X vssd1 vssd1 vccd1 vccd1 _8477_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6066_ _6302_/A _6066_/B vssd1 vssd1 vccd1 vccd1 _6066_/X sky130_fd_sc_hd__or2_1
Xhold1013 _8483_/Q vssd1 vssd1 vccd1 vccd1 _7025_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5274__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1035 _7811_/Q vssd1 vssd1 vccd1 vccd1 _5631_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _5418_/A _5451_/C vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__or2_1
Xhold1046 _5257_/X vssd1 vssd1 vccd1 vccd1 _7465_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 _7497_/Q vssd1 vssd1 vccd1 vccd1 _5293_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 _8174_/Q vssd1 vssd1 vccd1 vccd1 _6620_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 _6773_/X vssd1 vssd1 vccd1 vccd1 _8324_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6774__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6968_ _7027_/A _6968_/A2 _6970_/A3 _6967_/X vssd1 vssd1 vccd1 vccd1 _6968_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5919_ _5921_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5922_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7096__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6899_ _6965_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6899_/X sky130_fd_sc_hd__and2_1
XFILLER_0_134_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5329__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4632__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4659__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold891 _8297_/Q vssd1 vssd1 vccd1 vccd1 hold891/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold880 _5611_/X vssd1 vssd1 vccd1 vccd1 _7795_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5063__B _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5265__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4699__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4068__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1580 _4222_/Y vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6175__A _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5510__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1591 _4330_/Y vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6214__B1 _5739_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output108_A _7303_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6903__A _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6765__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4871__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4926__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4250_ _4250_/A _7644_/Q vssd1 vssd1 vccd1 vccd1 _4250_/Y sky130_fd_sc_hd__nand2_1
X_4181_ _8513_/Q _4181_/B vssd1 vssd1 vccd1 vccd1 _4181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_129_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4059__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5256__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7940_ _8079_/CLK _7940_/D vssd1 vssd1 vccd1 vccd1 _7940_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__5420__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7871_ _7871_/CLK _7871_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6822_ _7026_/A _6822_/A2 _6838_/A3 _6821_/X vssd1 vssd1 vccd1 vccd1 _6822_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6813__A _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6753_ _6929_/A _6741_/B _6774_/B1 hold619/X vssd1 vssd1 vccd1 vccd1 _6753_/X sky130_fd_sc_hd__a22o_1
X_3965_ _8071_/Q _3964_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3965_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6684_ _6935_/A _6669_/B _6702_/B1 hold451/X vssd1 vssd1 vccd1 vccd1 _6684_/X sky130_fd_sc_hd__a22o_1
X_5704_ _5697_/X _5703_/X _6028_/S vssd1 vssd1 vccd1 vccd1 _5704_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3896_ _3896_/A _3896_/B _4132_/A _3896_/D vssd1 vssd1 vccd1 vccd1 _3897_/D sky130_fd_sc_hd__or4_1
XFILLER_0_18_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8423_ _8468_/CLK _8423_/D vssd1 vssd1 vccd1 vccd1 _8423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5635_ _6935_/A _5620_/B _5653_/B1 hold835/X vssd1 vssd1 vccd1 vccd1 _5635_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3990__B2 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4614__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout306_A _5582_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8354_ _8354_/CLK _8354_/D vssd1 vssd1 vccd1 vccd1 _8354_/Q sky130_fd_sc_hd__dfxtp_1
Xhold110 _7756_/Q vssd1 vssd1 vccd1 vccd1 _6507_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5566_ _6545_/A _5566_/B vssd1 vssd1 vccd1 vccd1 _7755_/D sky130_fd_sc_hd__and2_1
XFILLER_0_130_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold121 _6497_/X vssd1 vssd1 vccd1 vccd1 _7979_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _5389_/A _5404_/C vssd1 vssd1 vccd1 vccd1 _5409_/A sky130_fd_sc_hd__nand2b_2
Xhold132 _7745_/Q vssd1 vssd1 vccd1 vccd1 _6496_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 _5685_/X vssd1 vssd1 vccd1 vccd1 _7865_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8285_ _8346_/CLK _8285_/D vssd1 vssd1 vccd1 vccd1 _8285_/Q sky130_fd_sc_hd__dfxtp_1
X_7305_ _8379_/CLK _7305_/D _7115_/Y vssd1 vssd1 vccd1 vccd1 _7305_/Q sky130_fd_sc_hd__dfrtp_4
X_5497_ _7518_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7686_/D sky130_fd_sc_hd__and3_1
XANTENNA__3742__B2 _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3742__A1 _4771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 _6500_/X vssd1 vssd1 vccd1 vccd1 _7982_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _4448_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4448_/X sky130_fd_sc_hd__and2_1
Xhold176 _7628_/Q vssd1 vssd1 vccd1 vccd1 _5686_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _7623_/Q vssd1 vssd1 vccd1 vccd1 _5681_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6692__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold187 _5687_/X vssd1 vssd1 vccd1 vccd1 _7867_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4917__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold198 _7334_/Q vssd1 vssd1 vccd1 vccd1 _5431_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4379_ _4379_/A _5069_/S vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__and2_1
X_7098_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7098_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6039__A3 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6118_ _6119_/A _6119_/B vssd1 vssd1 vccd1 vccd1 _6118_/Y sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6049_ _5734_/A _6038_/X _6048_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6049_/Y sky130_fd_sc_hd__o22ai_1
XFILLER_0_96_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4942__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6747__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4853__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4605__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3981__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5505__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6683__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5238__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6617__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4852__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6738__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6199__C1 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6633__A _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3750_ _3750_/A _3750_/B _4138_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__or3_1
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5961__A2 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3681_ _7282_/Q _3923_/B vssd1 vssd1 vccd1 vccd1 _3681_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_55_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6910__A1 _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5420_ _5420_/A _7073_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _5420_/X sky130_fd_sc_hd__and3_1
XANTENNA__5174__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5351_ _6937_/A _5335_/B _5368_/B1 hold875/X vssd1 vssd1 vccd1 vccd1 _5351_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5415__C _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8070_ _8469_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 _8070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5282_ _6945_/A _5294_/A2 _5294_/B1 hold577/X vssd1 vssd1 vccd1 vccd1 _5282_/X sky130_fd_sc_hd__a22o_1
X_4302_ _4302_/A _4302_/B vssd1 vssd1 vccd1 vccd1 _4302_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__6674__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4233_ _4232_/X _4421_/A _5453_/B vssd1 vssd1 vccd1 vccd1 _4422_/B sky130_fd_sc_hd__mux2_1
X_7021_ _7024_/A _7021_/B vssd1 vssd1 vccd1 vccd1 _7021_/X sky130_fd_sc_hd__and2_1
XFILLER_0_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5229__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4164_ _4449_/A _4449_/B vssd1 vssd1 vccd1 vccd1 _4164_/Y sky130_fd_sc_hd__nand2_1
X_4095_ _4095_/A vssd1 vssd1 vccd1 vccd1 _4095_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_4_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5431__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7923_ _8010_/CLK _7923_/D vssd1 vssd1 vccd1 vccd1 _7923_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout256_A _5584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7854_ _8071_/CLK _7854_/D vssd1 vssd1 vccd1 vccd1 _7854_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6729__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6805_ _6937_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6805_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7785_ _8431_/CLK _7785_/D vssd1 vssd1 vccd1 vccd1 _7785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout423_A _7357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4835__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7077__C _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4997_ _8487_/Q _8419_/Q _8451_/Q _8325_/Q _4997_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4997_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6736_ _6967_/A _6737_/A2 _6737_/B1 hold653/X vssd1 vssd1 vccd1 vccd1 _6736_/X sky130_fd_sc_hd__a22o_1
X_3948_ _4745_/B _3676_/A _4082_/B1 _3939_/C _3947_/X vssd1 vssd1 vccd1 vccd1 _5765_/A
+ sky130_fd_sc_hd__o221a_4
X_6667_ _6842_/C _6704_/B vssd1 vssd1 vccd1 vccd1 _6667_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_46_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3879_ _3879_/A1 _4073_/A2 _6955_/A _4073_/B2 _3878_/X vssd1 vssd1 vccd1 vccd1 _6444_/B
+ sky130_fd_sc_hd__a221o_1
X_5618_ _6776_/A _6842_/C vssd1 vssd1 vccd1 vccd1 _5618_/Y sky130_fd_sc_hd__nor2_2
X_6598_ _6596_/Y _6597_/Y _6593_/X vssd1 vssd1 vccd1 vccd1 _6598_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_61_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8406_ _8476_/CLK _8406_/D vssd1 vssd1 vccd1 vccd1 _8406_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5549_ _5667_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _5549_/X sky130_fd_sc_hd__and2_1
X_8337_ _8467_/CLK _8337_/D vssd1 vssd1 vccd1 vccd1 _8337_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8268_ _8462_/CLK _8268_/D vssd1 vssd1 vccd1 vccd1 _8268_/Q sky130_fd_sc_hd__dfxtp_1
X_8199_ _8326_/CLK _8199_/D vssd1 vssd1 vccd1 vccd1 _8199_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout420 _7357_/Q vssd1 vssd1 vccd1 vccd1 _4996_/S0 sky130_fd_sc_hd__buf_8
Xfanout431 _6660_/A1 vssd1 vssd1 vccd1 vccd1 _6434_/A sky130_fd_sc_hd__clkbuf_4
Xfanout453 _5667_/A vssd1 vssd1 vccd1 vccd1 _7006_/A sky130_fd_sc_hd__clkbuf_4
Xfanout464 _7281_/A vssd1 vssd1 vccd1 vccd1 _7279_/A sky130_fd_sc_hd__buf_8
Xfanout442 _7005_/A vssd1 vssd1 vccd1 vccd1 _6539_/A sky130_fd_sc_hd__clkbuf_4
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6968__A1 _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5768__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5640__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4672__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6453__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6172__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4826__S0 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3954__A1 _3953_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5156__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5516__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3890__B1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5631__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4582__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7217__95 _8096_/CLK vssd1 vssd1 vccd1 vccd1 _8130_/CLK sky130_fd_sc_hd__inv_2
X_4920_ _8476_/Q _8408_/Q _8440_/Q _8314_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4920_/X sky130_fd_sc_hd__mux4_1
X_4851_ _4850_/X _4849_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3802_ _8001_/Q _4068_/A2 _4068_/B1 _8033_/Q _3801_/X vssd1 vssd1 vccd1 vccd1 _3802_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6187__A2 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4782_ _4781_/X _4778_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8230_/D sky130_fd_sc_hd__mux2_1
X_7570_ _8175_/CLK _7570_/D vssd1 vssd1 vccd1 vccd1 _7570_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5934__A2 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6521_ _6552_/A _6521_/B vssd1 vssd1 vccd1 vccd1 _8003_/D sky130_fd_sc_hd__and2_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3733_ _6279_/A vssd1 vssd1 vccd1 vccd1 _3733_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3664_ _3661_/Y _7836_/Q _3653_/Y _7665_/Q vssd1 vssd1 vccd1 vccd1 _3669_/A sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_113_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6452_ _7022_/A _6452_/B vssd1 vssd1 vccd1 vccd1 _7934_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5403_ _7090_/A _6554_/B vssd1 vssd1 vccd1 vccd1 _7597_/D sky130_fd_sc_hd__nor2_2
XANTENNA__5698__A1 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5426__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8122_ _8122_/CLK _8122_/D vssd1 vssd1 vccd1 vccd1 _8122_/Q sky130_fd_sc_hd__dfxtp_2
X_6383_ _3836_/B _6292_/A _7279_/A vssd1 vssd1 vccd1 vccd1 _6383_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5334_ _6558_/A _6740_/C vssd1 vssd1 vccd1 vccd1 _5336_/B sky130_fd_sc_hd__or2_2
XFILLER_0_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8053_ _8053_/CLK _8053_/D vssd1 vssd1 vccd1 vccd1 _8053_/Q sky130_fd_sc_hd__dfxtp_1
X_5265_ _3939_/C _5263_/B _5263_/Y hold300/X vssd1 vssd1 vccd1 vccd1 _5265_/X sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6538__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7004_ _7008_/A _7004_/B vssd1 vssd1 vccd1 vccd1 _7004_/X sky130_fd_sc_hd__and2_1
X_4216_ _8508_/Q _4216_/B vssd1 vssd1 vccd1 vccd1 _4217_/B sky130_fd_sc_hd__nand2_1
X_5196_ _6921_/A _5221_/A2 _5221_/B1 hold667/X vssd1 vssd1 vccd1 vccd1 _5196_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6662__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4147_ _8455_/Q _5730_/A vssd1 vssd1 vccd1 vccd1 _5690_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__4058__A _4756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_A _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5622__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4078_ _3923_/B _7952_/Q vssd1 vssd1 vccd1 vccd1 _4078_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_92_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7906_ _8477_/CLK _7906_/D vssd1 vssd1 vccd1 vccd1 _7906_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4492__S _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7837_ _8079_/CLK _7837_/D vssd1 vssd1 vccd1 vccd1 _7837_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7088__B _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7231__109 _8448_/CLK vssd1 vssd1 vccd1 vccd1 _8241_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6178__A2 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4808__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7768_ _8030_/CLK _7768_/D vssd1 vssd1 vccd1 vccd1 _7768_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold1488_A _7311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6719_ _6933_/A _6705_/B _6738_/B1 hold439/X vssd1 vssd1 vccd1 vccd1 _6719_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7699_ _8419_/CLK _7699_/D vssd1 vssd1 vccd1 vccd1 _7699_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5138__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4361__A1 _7052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6448__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5310__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout250 _6669_/Y vssd1 vssd1 vccd1 vccd1 _6702_/B1 sky130_fd_sc_hd__buf_6
XFILLER_0_100_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout283 _6776_/X vssd1 vssd1 vccd1 vccd1 _6779_/B sky130_fd_sc_hd__buf_6
Xfanout272 _3841_/B vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__clkbuf_8
Xfanout261 _5262_/Y vssd1 vssd1 vccd1 vccd1 _5294_/B1 sky130_fd_sc_hd__buf_6
Xfanout294 _6602_/X vssd1 vssd1 vccd1 vccd1 _6605_/B sky130_fd_sc_hd__clkbuf_16
XANTENNA__7279__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5613__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6911__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold709 _7832_/Q vssd1 vssd1 vccd1 vccd1 hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6892__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5262__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5050_ _5050_/A1 _5067_/S _5172_/B1 _5049_/X vssd1 vssd1 vccd1 vccd1 _7337_/D sky130_fd_sc_hd__o211a_1
X_4001_ _7710_/Q _4081_/B vssd1 vssd1 vccd1 vccd1 _4001_/X sky130_fd_sc_hd__or2_1
Xhold1409 _4265_/Y vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6644__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3863__B1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_56_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6805__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5952_ _5952_/A _5952_/B vssd1 vssd1 vccd1 vccd1 _5953_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5604__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5080__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4903_ _8151_/Q _7550_/Q _7422_/Q _7582_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4903_/X sky130_fd_sc_hd__mux4_1
X_5883_ _3973_/X _6398_/A2 _6413_/B1 _6251_/A _6011_/A2 vssd1 vssd1 vccd1 vccd1 _5883_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4834_ _4832_/X _4833_/X _7359_/Q vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5368__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6821__A _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7622_ _8032_/CLK _7622_/D vssd1 vssd1 vccd1 vccd1 _7622_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7553_ _8154_/CLK _7553_/D vssd1 vssd1 vccd1 vccd1 _7553_/Q sky130_fd_sc_hd__dfxtp_1
X_4765_ _7019_/A _4765_/B vssd1 vssd1 vccd1 vccd1 _8122_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_114_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3716_ _7997_/Q _4068_/A2 _4068_/B1 _8029_/Q _3715_/X vssd1 vssd1 vccd1 vccd1 _3716_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6504_ _6545_/A hold37/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__and2_1
XFILLER_0_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6580__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4696_ _8158_/Q _7557_/Q _7429_/Q _7589_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4696_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7484_ _8472_/CLK _7484_/D vssd1 vssd1 vccd1 vccd1 _7484_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout219_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3647_ _7365_/Q vssd1 vssd1 vccd1 vccd1 _3647_/Y sky130_fd_sc_hd__inv_2
X_6435_ _7018_/A _6435_/B vssd1 vssd1 vccd1 vccd1 _7917_/D sky130_fd_sc_hd__and2_1
XFILLER_0_113_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6366_ _6356_/X _6360_/X _6363_/X _6364_/X _6365_/Y vssd1 vssd1 vccd1 vccd1 _7896_/D
+ sky130_fd_sc_hd__o41a_1
X_5317_ _6941_/A _5332_/A2 _5331_/B1 hold593/X vssd1 vssd1 vccd1 vccd1 _5317_/X sky130_fd_sc_hd__a22o_1
X_8105_ _8105_/CLK _8105_/D vssd1 vssd1 vccd1 vccd1 _8105_/Q sky130_fd_sc_hd__dfxtp_1
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_6297_ _6298_/A _6298_/B vssd1 vssd1 vccd1 vccd1 _6297_/Y sky130_fd_sc_hd__nand2_1
X_8036_ _8036_/CLK _8036_/D vssd1 vssd1 vccd1 vccd1 _8036_/Q sky130_fd_sc_hd__dfxtp_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _6949_/A _5258_/A2 _5258_/B1 hold394/X vssd1 vssd1 vccd1 vccd1 _5248_/X sky130_fd_sc_hd__a22o_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5179_ _5469_/A _5470_/C vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__or2_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6399__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7045__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7099__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1772_A _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5359__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4950__S _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6571__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5781__S _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6874__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6087__A1 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6087__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5513__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6626__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5810__A _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6625__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5598__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5062__A2 _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6641__A _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6562__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4161__A _4161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5770__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4550_ _4548_/X _4549_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold517 _7446_/Q vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
X_4481_ _7017_/A _7906_/Q vssd1 vssd1 vccd1 vccd1 _8038_/D sky130_fd_sc_hd__and2_1
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold506 _5205_/X vssd1 vssd1 vccd1 vccd1 _7419_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6220_ _3896_/B _6414_/A2 _6130_/X _6213_/X vssd1 vssd1 vccd1 vccd1 _6220_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold539 _7793_/Q vssd1 vssd1 vccd1 vccd1 hold539/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 _6694_/X vssd1 vssd1 vccd1 vccd1 _8221_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5392__C_N _5408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6151_ _6391_/A _6142_/Y _6150_/Y vssd1 vssd1 vccd1 vccd1 _6151_/Y sky130_fd_sc_hd__o21ai_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5102_ input12/X _5099_/B _5148_/B1 _5101_/X vssd1 vssd1 vccd1 vccd1 _7363_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6082_ _5907_/X _6081_/Y _6342_/S vssd1 vssd1 vccd1 vccd1 _6083_/B sky130_fd_sc_hd__mux2_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _6918_/X vssd1 vssd1 vccd1 vccd1 _8424_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1217 _8416_/Q vssd1 vssd1 vccd1 vccd1 _6900_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 _6954_/X vssd1 vssd1 vccd1 vccd1 _8442_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5033_ _5426_/A _5462_/C vssd1 vssd1 vccd1 vccd1 _5033_/X sky130_fd_sc_hd__or2_1
Xhold1239 _8403_/Q vssd1 vssd1 vccd1 vccd1 _6874_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5589__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6984_ _7074_/A _6983_/X _6990_/S vssd1 vssd1 vccd1 vccd1 _6985_/B sky130_fd_sc_hd__mux2_1
XANTENNA_fanout169_A _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5935_ _5791_/Y _5934_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _5936_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_75_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5866_ _5845_/Y _5850_/B _5847_/B vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout336_A _3814_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6551__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _8034_/CLK sky130_fd_sc_hd__clkbuf_16
X_4817_ _4816_/X _4813_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8235_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7605_ _8363_/CLK _7605_/D vssd1 vssd1 vccd1 vccd1 _7605_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5797_ _5698_/X _5700_/X _5797_/S vssd1 vssd1 vccd1 vccd1 _5797_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _6551_/A _4748_/B vssd1 vssd1 vccd1 vccd1 _8105_/D sky130_fd_sc_hd__and2_1
X_7536_ _8355_/CLK _7536_/D vssd1 vssd1 vccd1 vccd1 _7536_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7467_ _8451_/CLK _7467_/D vssd1 vssd1 vccd1 vccd1 _7467_/Q sky130_fd_sc_hd__dfxtp_1
X_4679_ _4678_/X _4677_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4679_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6856__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6418_ _6534_/A _6418_/B vssd1 vssd1 vccd1 vccd1 _6418_/X sky130_fd_sc_hd__and2_1
XFILLER_0_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7398_ _8008_/CLK _7398_/D vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_6349_ _6333_/Y _6338_/B _6335_/B vssd1 vssd1 vccd1 vccd1 _6355_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_12_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8019_ _8019_/CLK _8019_/D vssd1 vssd1 vccd1 vccd1 _8019_/Q sky130_fd_sc_hd__dfxtp_1
X_7237__115 _8473_/CLK vssd1 vssd1 vccd1 vccd1 _8247_/CLK sky130_fd_sc_hd__inv_2
Xhold1751 _8510_/Q vssd1 vssd1 vccd1 vccd1 _4040_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1740 _4021_/B vssd1 vssd1 vccd1 vccd1 _5988_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1762 _3799_/B vssd1 vssd1 vccd1 vccd1 _6204_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5292__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6445__B _6445_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1784 _3996_/B vssd1 vssd1 vccd1 vccd1 _5916_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1795 _8455_/Q vssd1 vssd1 vccd1 vccd1 _5731_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1773 _6240_/Y vssd1 vssd1 vccd1 vccd1 _7889_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5044__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6461__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4680__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8421_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4650__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5524__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4855__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5283__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4156__A _8516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6232__A1 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3981_ _3981_/A1 _4084_/A2 _6923_/A _4084_/B2 _3980_/X vssd1 vssd1 vccd1 vccd1 _3981_/X
+ sky130_fd_sc_hd__a221o_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3995__A _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5720_ _5704_/X _5719_/X _6251_/A vssd1 vssd1 vccd1 vccd1 _5721_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_9_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_42_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _8339_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5651_ _6967_/A _5652_/A2 _5652_/B1 hold605/X vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__a22o_1
X_5582_ _6740_/C _6704_/B vssd1 vssd1 vccd1 vccd1 _5582_/Y sky130_fd_sc_hd__nor2_2
X_8370_ _8370_/CLK _8370_/D _7264_/Y vssd1 vssd1 vccd1 vccd1 _8370_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5418__C _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4602_ _4601_/X _4600_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4602_/X sky130_fd_sc_hd__mux2_1
X_4533_ _4532_/X _4529_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7501_/D sky130_fd_sc_hd__mux2_1
X_7321_ _8365_/CLK _7321_/D vssd1 vssd1 vccd1 vccd1 _7321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold314 _7318_/Q vssd1 vssd1 vccd1 vccd1 _5415_/A sky130_fd_sc_hd__dlygate4sd3_1
X_7252_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7252_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold325 _5462_/X vssd1 vssd1 vccd1 vccd1 _7651_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold303 _5464_/X vssd1 vssd1 vccd1 vccd1 _7653_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _7437_/Q vssd1 vssd1 vccd1 vccd1 hold358/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold369 _5423_/X vssd1 vssd1 vccd1 vccd1 _7612_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _7343_/Q vssd1 vssd1 vccd1 vccd1 _5440_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6391_/A _6194_/X _6201_/Y _6202_/Y vssd1 vssd1 vccd1 vccd1 _6203_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4464_ _7018_/A _7923_/Q vssd1 vssd1 vccd1 vccd1 _8055_/D sky130_fd_sc_hd__and2_1
Xhold347 _5426_/X vssd1 vssd1 vccd1 vccd1 _7615_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6838__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5434__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4395_ _4398_/A _4395_/B vssd1 vssd1 vccd1 vccd1 _4395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6134_ _4077_/B _6417_/A2 _7267_/A vssd1 vssd1 vccd1 vccd1 _6134_/Y sky130_fd_sc_hd__a21oi_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6546__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6065_ _5981_/X _6064_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6066_/B sky130_fd_sc_hd__mux2_1
Xhold1003 _7809_/Q vssd1 vssd1 vccd1 vccd1 _5629_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1014 _7025_/X vssd1 vssd1 vccd1 vccd1 _8483_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout286_A _6775_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5274__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1025 _7576_/Q vssd1 vssd1 vccd1 vccd1 _5349_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _5631_/X vssd1 vssd1 vccd1 vccd1 _7811_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 _8461_/Q vssd1 vssd1 vccd1 vccd1 _7003_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5016_ _4434_/A _4448_/B _5140_/B1 _5015_/X vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3889__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1058 _5293_/X vssd1 vssd1 vccd1 vccd1 _7497_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1069 _8484_/Q vssd1 vssd1 vccd1 vccd1 _7026_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout453_A _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5026__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6967_ _6967_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6967_/X sky130_fd_sc_hd__and2_1
X_5918_ _5918_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _5921_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__6774__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6281__A _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_33_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8332_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7178__56 _8480_/CLK vssd1 vssd1 vccd1 vccd1 _8058_/CLK sky130_fd_sc_hd__inv_2
X_6898_ _7025_/A _6898_/A2 _6906_/A3 _6897_/X vssd1 vssd1 vccd1 vccd1 _6898_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5849_ _5850_/A _5850_/B vssd1 vssd1 vccd1 vccd1 _5849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1470_A _7300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4005__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7519_ _7519_/CLK _7519_/D vssd1 vssd1 vccd1 vccd1 _7519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4632__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8499_ _8501_/CLK _8499_/D vssd1 vssd1 vccd1 vccd1 _8499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold881 _8313_/Q vssd1 vssd1 vccd1 vccd1 hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold870 _6584_/X vssd1 vssd1 vccd1 vccd1 _8156_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 _6746_/X vssd1 vssd1 vccd1 vccd1 _8297_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4699__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1570 _7370_/Q vssd1 vssd1 vccd1 vccd1 _7076_/A sky130_fd_sc_hd__clkbuf_4
Xhold1581 _4231_/X vssd1 vssd1 vccd1 vccd1 _4232_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1592 _4332_/X vssd1 vssd1 vccd1 vccd1 _5576_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6191__A _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6903__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6765__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8425_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5519__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5725__B1 _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3754__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7192__70 _8071_/CLK vssd1 vssd1 vccd1 vccd1 _8105_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_1_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6150__B1 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4180_ _4180_/A _4181_/B vssd1 vssd1 vccd1 vccd1 _4180_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4585__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5256__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7870_ _8270_/CLK _7870_/D vssd1 vssd1 vccd1 vccd1 _7870_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5008__A2 _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6821_ _6953_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6821_/X sky130_fd_sc_hd__and2_1
XANTENNA__6756__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6813__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6752_ _6927_/A _6741_/B _6774_/B1 hold733/X vssd1 vssd1 vccd1 vccd1 _6752_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_15_clk _7871_/CLK vssd1 vssd1 vccd1 vccd1 _8451_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3964_ _7975_/Q _4068_/A2 _4068_/B1 _8007_/Q _3963_/X vssd1 vssd1 vccd1 vccd1 _3964_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_128_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6683_ _6933_/A _6669_/B _6702_/B1 hold342/X vssd1 vssd1 vccd1 vccd1 _6683_/X sky130_fd_sc_hd__a22o_1
X_5703_ _5699_/X _5702_/X _5879_/S vssd1 vssd1 vccd1 vccd1 _5703_/X sky130_fd_sc_hd__mux2_1
X_3895_ _3895_/A _3895_/B vssd1 vssd1 vccd1 vccd1 _3896_/D sky130_fd_sc_hd__and2_1
XANTENNA__5429__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8422_ _8468_/CLK _8422_/D vssd1 vssd1 vccd1 vccd1 _8422_/Q sky130_fd_sc_hd__dfxtp_1
X_5634_ _6933_/A _5620_/B _5653_/B1 hold431/X vssd1 vssd1 vccd1 vccd1 _5634_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3990__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6064__S0 _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5716__A0 _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5192__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4614__S1 _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8353_ _8353_/CLK _8353_/D vssd1 vssd1 vccd1 vccd1 _8353_/Q sky130_fd_sc_hd__dfxtp_1
Xhold100 _7844_/Q vssd1 vssd1 vccd1 vccd1 _6465_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5565_ _7022_/A _5565_/B vssd1 vssd1 vccd1 vccd1 _7754_/D sky130_fd_sc_hd__and2_1
X_7304_ _8378_/CLK _7304_/D _7114_/Y vssd1 vssd1 vccd1 vccd1 _7304_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_130_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5496_ _7517_/Q _5542_/B _7088_/B vssd1 vssd1 vccd1 vccd1 _7685_/D sky130_fd_sc_hd__and3_1
Xhold144 _7606_/Q vssd1 vssd1 vccd1 vccd1 _5664_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _5391_/A _5408_/B _6553_/A vssd1 vssd1 vccd1 vccd1 _5404_/C sky130_fd_sc_hd__and3b_1
Xhold133 _6496_/X vssd1 vssd1 vccd1 vccd1 _7978_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 _6507_/X vssd1 vssd1 vccd1 vccd1 _7989_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8284_ _8442_/CLK _8284_/D vssd1 vssd1 vccd1 vccd1 _8284_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold122 _7622_/Q vssd1 vssd1 vccd1 vccd1 _5680_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3742__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4447_ _4171_/Y _7030_/C _4446_/X _4445_/X vssd1 vssd1 vccd1 vccd1 _8360_/D sky130_fd_sc_hd__a31o_1
Xhold177 _5686_/X vssd1 vssd1 vccd1 vccd1 _7866_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _5681_/X vssd1 vssd1 vccd1 vccd1 _7861_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold166 _7855_/Q vssd1 vssd1 vccd1 vccd1 _6476_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6692__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold188 _7765_/Q vssd1 vssd1 vccd1 vccd1 _6516_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold199 _5431_/X vssd1 vssd1 vccd1 vccd1 _7620_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6117_ _6098_/A _6097_/A _6097_/B vssd1 vssd1 vccd1 vccd1 _6119_/B sky130_fd_sc_hd__a21bo_1
X_4378_ _5058_/A1 _4377_/Y _5468_/C vssd1 vssd1 vccd1 vccd1 _8385_/D sky130_fd_sc_hd__mux2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7097_/Y sky130_fd_sc_hd__inv_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5247__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6048_ _5840_/A _6309_/B _6047_/Y _6128_/A vssd1 vssd1 vccd1 vccd1 _6048_/X sky130_fd_sc_hd__o22a_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7999_ _8494_/CLK hold88/X vssd1 vssd1 vccd1 vccd1 _7999_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6747__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4853__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3981__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4605__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5238__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5521__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4541__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6738__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6199__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6633__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5410__A2 _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5961__A3 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3972__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3774__B1_N _3773_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3680_ _4067_/A_N _7964_/Q vssd1 vssd1 vccd1 vccd1 _3680_/X sky130_fd_sc_hd__and2b_1
X_5350_ _6935_/A _5335_/B _5368_/B1 hold977/X vssd1 vssd1 vccd1 vccd1 _5350_/X sky130_fd_sc_hd__a22o_1
X_5281_ _6877_/A _5262_/B _5295_/B1 _5281_/B2 vssd1 vssd1 vccd1 vccd1 _5281_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_64_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4301_ _4291_/Y _4295_/B _4293_/B vssd1 vssd1 vccd1 vccd1 _4302_/B sky130_fd_sc_hd__o21a_1
XANTENNA__6674__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4232_ _4232_/A _4232_/B vssd1 vssd1 vccd1 vccd1 _4232_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_57_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7020_ _7026_/A _7020_/B vssd1 vssd1 vccd1 vccd1 _7020_/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_4_clk clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _8431_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4780__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4163_ _4449_/B vssd1 vssd1 vccd1 vccd1 _4163_/Y sky130_fd_sc_hd__inv_2
X_4094_ _5789_/S _4094_/B _5838_/A vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__or3_2
X_7922_ _8472_/CLK _7922_/D vssd1 vssd1 vccd1 vccd1 _7922_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7853_ _8379_/CLK _7853_/D vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__6729__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6804_ _7029_/A _6804_/A2 _6776_/X _6803_/X vssd1 vssd1 vccd1 vccd1 _6804_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4996_ _8197_/Q _8229_/Q _8293_/Q _7801_/Q _4996_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4996_/X sky130_fd_sc_hd__mux4_1
X_7784_ _8402_/CLK _7784_/D vssd1 vssd1 vccd1 vccd1 _7784_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout249_A _6669_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3947_ _3947_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _3947_/X sky130_fd_sc_hd__or2_1
XANTENNA__4835__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6735_ _6965_/A _6737_/A2 _6737_/B1 hold771/X vssd1 vssd1 vccd1 vccd1 _6735_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_135_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7148__26 _8319_/CLK vssd1 vssd1 vccd1 vccd1 _7525_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6666_ _7029_/A _6666_/A2 _6666_/A3 _6665_/X vssd1 vssd1 vccd1 vccd1 _6666_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout416_A _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3878_ _4767_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__and2_1
X_8405_ _8473_/CLK _8405_/D vssd1 vssd1 vccd1 vccd1 _8405_/Q sky130_fd_sc_hd__dfxtp_1
X_6597_ _6977_/B _6597_/B vssd1 vssd1 vccd1 vccd1 _6597_/Y sky130_fd_sc_hd__nor2_1
X_5617_ _6971_/A _5584_/B _5617_/B1 hold689/X vssd1 vssd1 vccd1 vccd1 _5617_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8336_ _8466_/CLK _8336_/D vssd1 vssd1 vccd1 vccd1 _8336_/Q sky130_fd_sc_hd__dfxtp_1
X_5548_ _7090_/A _5548_/B vssd1 vssd1 vccd1 vccd1 _7737_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_112_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8267_ _8425_/CLK _8267_/D vssd1 vssd1 vccd1 vccd1 _8267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5479_ _7500_/Q _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7668_/D sky130_fd_sc_hd__and3_1
X_8198_ _8326_/CLK _8198_/D vssd1 vssd1 vccd1 vccd1 _8198_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout410 _4997_/S1 vssd1 vssd1 vccd1 vccd1 _4952_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout421 _7357_/Q vssd1 vssd1 vccd1 vccd1 _4997_/S0 sky130_fd_sc_hd__buf_4
Xfanout432 _7023_/A vssd1 vssd1 vccd1 vccd1 _7017_/A sky130_fd_sc_hd__buf_4
Xfanout454 _5667_/A vssd1 vssd1 vccd1 vccd1 _6999_/A sky130_fd_sc_hd__buf_4
Xfanout465 input63/X vssd1 vssd1 vccd1 vccd1 _7281_/A sky130_fd_sc_hd__clkbuf_8
Xfanout443 _6660_/A1 vssd1 vssd1 vccd1 vccd1 _7005_/A sky130_fd_sc_hd__clkbuf_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4523__S0 _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4428__B1 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4953__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4826__S1 _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5516__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7162__40 _8090_/CLK vssd1 vssd1 vccd1 vccd1 _8042_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6909__A _6909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6656__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5532__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7081__B2 _7044_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3890__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5092__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5631__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4850_ _8466_/Q _8398_/Q _8430_/Q _8304_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4850_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_0_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3801_ _4067_/A_N _7969_/Q vssd1 vssd1 vccd1 vccd1 _3801_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4781_ _4780_/X _4779_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__mux2_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5934__A3 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6520_ _6520_/A hold81/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__and2_1
XFILLER_0_7_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3732_ _3968_/A _6445_/B _3731_/Y vssd1 vssd1 vccd1 vccd1 _6279_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3663_ _7665_/Q _7664_/Q _7667_/Q _7666_/Q vssd1 vssd1 vccd1 vccd1 _3663_/X sky130_fd_sc_hd__or4_1
X_6451_ _6520_/A _6451_/B vssd1 vssd1 vccd1 vccd1 _7933_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5402_ _6553_/A _5402_/B vssd1 vssd1 vccd1 vccd1 _6554_/B sky130_fd_sc_hd__or2_1
X_6382_ _6391_/A _6373_/Y _6377_/X vssd1 vssd1 vccd1 vccd1 _6382_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5333_ _6558_/A _6740_/C vssd1 vssd1 vccd1 vccd1 _5333_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8121_ _8121_/CLK _8121_/D vssd1 vssd1 vccd1 vccd1 _8121_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6819__A _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8052_ _8052_/CLK _8052_/D vssd1 vssd1 vccd1 vccd1 _8052_/Q sky130_fd_sc_hd__dfxtp_1
X_5264_ _6777_/A _5262_/B _5295_/B1 hold352/X vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__a22o_1
X_4215_ _8508_/Q _4216_/B vssd1 vssd1 vccd1 vccd1 _4215_/Y sky130_fd_sc_hd__nor2_1
X_7003_ _7019_/A _7003_/B vssd1 vssd1 vccd1 vccd1 _7003_/X sky130_fd_sc_hd__and2_1
X_5195_ _6853_/A _5221_/A2 _5221_/B1 hold473/X vssd1 vssd1 vccd1 vccd1 _5195_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5442__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout199_A _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4146_ _5730_/A _5738_/A vssd1 vssd1 vccd1 vccd1 _5723_/B sky130_fd_sc_hd__nand2b_2
XANTENNA__4058__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6554__A _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7072__B2 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _4077_/A _4077_/B vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__and2_1
XFILLER_0_92_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7905_ _8480_/CLK _7905_/D vssd1 vssd1 vccd1 vccd1 _7905_/Q sky130_fd_sc_hd__dfxtp_1
X_7836_ _8456_/CLK _7836_/D vssd1 vssd1 vccd1 vccd1 _7836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6178__A3 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4808__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7767_ _8385_/CLK _7767_/D vssd1 vssd1 vccd1 vccd1 _7767_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6583__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4979_ _8355_/Q _7831_/Q _7497_/Q _7465_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4979_/X sky130_fd_sc_hd__mux4_1
X_7698_ _8354_/CLK _7698_/D vssd1 vssd1 vccd1 vccd1 _7698_/Q sky130_fd_sc_hd__dfxtp_1
X_6718_ _6931_/A _6737_/A2 _6737_/B1 hold863/X vssd1 vssd1 vccd1 vccd1 _6718_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_116_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6649_ _6955_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6649_/X sky130_fd_sc_hd__and2_1
XFILLER_0_131_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6886__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6638__A1 _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8319_ _8319_/CLK _8319_/D vssd1 vssd1 vccd1 vccd1 _8319_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6448__B _6448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5310__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout240 _5144_/A2 vssd1 vssd1 vccd1 vccd1 _4425_/B sky130_fd_sc_hd__buf_4
XANTENNA__4113__A2 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 _5262_/Y vssd1 vssd1 vccd1 vccd1 _5295_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout273 _3676_/A vssd1 vssd1 vccd1 vccd1 _4071_/A2 sky130_fd_sc_hd__buf_8
Xfanout251 _6559_/Y vssd1 vssd1 vccd1 vccd1 _6591_/B1 sky130_fd_sc_hd__buf_6
XANTENNA__5779__S _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout295 _6661_/B vssd1 vssd1 vccd1 vccd1 _6665_/B sky130_fd_sc_hd__clkbuf_8
Xfanout284 _6776_/X vssd1 vssd1 vccd1 vccd1 _6838_/A3 sky130_fd_sc_hd__buf_6
XANTENNA__5074__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6464__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4683__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6271__C1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6810__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5613__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6574__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5527__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6326__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6639__A _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4858__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4983__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5301__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5262__B _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4000_ _8077_/Q _3999_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4000_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3863__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5951_ _6411_/S _5951_/B vssd1 vssd1 vccd1 vccd1 _5957_/A sky130_fd_sc_hd__nand2_1
XANTENNA__5604__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4902_ _8344_/Q _7820_/Q _7486_/Q _7454_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4902_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5882_ _5873_/X _5875_/X _5879_/X _5880_/X _6028_/S _6198_/S vssd1 vssd1 vccd1 vccd1
+ _5882_/X sky130_fd_sc_hd__mux4_1
X_4833_ _8141_/Q _7540_/Q _7412_/Q _7572_/Q _7357_/Q _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4833_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5368__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7621_ _8090_/CLK _7621_/D vssd1 vssd1 vccd1 vccd1 _7621_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6821__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6565__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4040__A1 _4039_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4764_ _7024_/A _4764_/B vssd1 vssd1 vccd1 vccd1 _8121_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7552_ _8471_/CLK _7552_/D vssd1 vssd1 vccd1 vccd1 _7552_/Q sky130_fd_sc_hd__dfxtp_1
X_6503_ _6548_/A _6503_/B vssd1 vssd1 vccd1 vccd1 _6503_/X sky130_fd_sc_hd__and2_1
XANTENNA__5437__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3715_ _4067_/A_N _7965_/Q vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__and2b_1
X_7483_ _8471_/CLK _7483_/D vssd1 vssd1 vccd1 vccd1 _7483_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6868__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4695_ _8351_/Q _7827_/Q _7493_/Q _7461_/Q _4741_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4695_/X sky130_fd_sc_hd__mux4_1
X_6434_ _6434_/A _6434_/B vssd1 vssd1 vccd1 vccd1 _7916_/D sky130_fd_sc_hd__and2_1
XFILLER_0_102_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3646_ _7273_/A vssd1 vssd1 vccd1 vccd1 _3646_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6549__A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6365_ _3823_/B _5734_/X _7279_/A vssd1 vssd1 vccd1 vccd1 _6365_/Y sky130_fd_sc_hd__a21oi_1
X_8104_ _8104_/CLK hold6/A vssd1 vssd1 vccd1 vccd1 _8104_/Q sky130_fd_sc_hd__dfxtp_1
X_6296_ _6298_/A _6298_/B vssd1 vssd1 vccd1 vccd1 _6299_/A sky130_fd_sc_hd__and2_1
X_5316_ _6939_/A _5299_/B _5331_/B1 hold511/X vssd1 vssd1 vccd1 vccd1 _5316_/X sky130_fd_sc_hd__a22o_1
X_5247_ _6947_/A _5258_/A2 _5258_/B1 hold975/X vssd1 vssd1 vccd1 vccd1 _5247_/X sky130_fd_sc_hd__a22o_1
X_8035_ _8035_/CLK _8035_/D vssd1 vssd1 vccd1 vccd1 _8035_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4726__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _5178_/A1 _5069_/S _5182_/B1 _5177_/X vssd1 vssd1 vccd1 vccd1 _7401_/D sky130_fd_sc_hd__o211a_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5056__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4129_ _6244_/A _6242_/A vssd1 vssd1 vccd1 vccd1 _4129_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4516__B _5408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7819_ _8343_/CLK _7819_/D vssd1 vssd1 vccd1 vccd1 _7819_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5359__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1765_A _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6308__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3790__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4055__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7132__10 _8343_/CLK vssd1 vssd1 vccd1 vccd1 _7509_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6459__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4965__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5295__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4717__S0 _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6641__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4480_ _6999_/A _7907_/Q vssd1 vssd1 vccd1 vccd1 _8039_/D sky130_fd_sc_hd__and2_1
XFILLER_0_123_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold518 _5238_/X vssd1 vssd1 vccd1 vccd1 _7446_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3781__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold507 _7796_/Q vssd1 vssd1 vccd1 vccd1 hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _8201_/Q vssd1 vssd1 vccd1 vccd1 hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4588__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6369__A _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7903__D _7903_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6150_ _6309_/A _5719_/X _6130_/A vssd1 vssd1 vccd1 vccd1 _6150_/Y sky130_fd_sc_hd__o21ai_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5101_ _5472_/A _5523_/C vssd1 vssd1 vccd1 vccd1 _5101_/X sky130_fd_sc_hd__or2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 _8357_/Q vssd1 vssd1 vccd1 vccd1 _6840_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_6081_ _5963_/S _6079_/X _6080_/X vssd1 vssd1 vccd1 vccd1 _6081_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5825__A2 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1218 _6900_/X vssd1 vssd1 vccd1 vccd1 _8416_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _4412_/A _4416_/B _5166_/B1 _5031_/X vssd1 vssd1 vccd1 vccd1 _7328_/D sky130_fd_sc_hd__o211a_1
Xhold1229 _8435_/Q vssd1 vssd1 vccd1 vccd1 _6940_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5589__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5038__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6983_ _6982_/X _6983_/B vssd1 vssd1 vccd1 vccd1 _6983_/X sky130_fd_sc_hd__and2b_1
X_5934_ _5846_/A _5870_/A _5892_/A _5921_/A _5772_/S _5804_/A vssd1 vssd1 vccd1 vccd1
+ _5934_/X sky130_fd_sc_hd__mux4_1
X_5865_ _3910_/A _6063_/A _5864_/Y _6741_/A vssd1 vssd1 vccd1 vccd1 _7871_/D sky130_fd_sc_hd__a211oi_1
XANTENNA_fanout231_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4078__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4816_ _4815_/X _4814_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__mux2_1
X_7604_ _7977_/CLK _7604_/D vssd1 vssd1 vccd1 vccd1 _7604_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout329_A _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5796_ _5794_/X _5795_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5796_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5210__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7535_ _8136_/CLK _7535_/D vssd1 vssd1 vccd1 vccd1 _7535_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4747_ _7029_/A hold5/X vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__and2_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7466_ _8467_/CLK _7466_/D vssd1 vssd1 vccd1 vccd1 _7466_/Q sky130_fd_sc_hd__dfxtp_1
X_4678_ _8478_/Q _8410_/Q _8442_/Q _8316_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4678_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6710__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6417_ _6417_/A1 _6417_/A2 _6408_/X _6416_/Y _7279_/A vssd1 vssd1 vccd1 vccd1 _6417_/Y
+ sky130_fd_sc_hd__a221oi_1
XANTENNA__4947__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7397_ _8091_/CLK _7397_/D vssd1 vssd1 vccd1 vccd1 _7397_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5183__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6348_ _6339_/Y _6343_/X _6344_/Y _6346_/X _6347_/Y vssd1 vssd1 vccd1 vccd1 _7895_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5277__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6279_ _6279_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6281_/B sky130_fd_sc_hd__xnor2_1
X_8018_ _8019_/CLK _8018_/D vssd1 vssd1 vccd1 vccd1 _8018_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1741 _5989_/X vssd1 vssd1 vccd1 vccd1 _7876_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1752 _4044_/B vssd1 vssd1 vccd1 vccd1 _6011_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1730 _7727_/Q vssd1 vssd1 vccd1 vccd1 _3741_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1796 _7880_/Q vssd1 vssd1 vccd1 vccd1 hold1796/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1774 _7702_/Q vssd1 vssd1 vccd1 vccd1 _3914_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1763 _6204_/Y vssd1 vssd1 vccd1 vccd1 _7887_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1785 _7723_/Q vssd1 vssd1 vccd1 vccd1 _3876_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4246__B _4246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6742__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6792__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_40_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5201__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_55_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6189__A _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4938__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6701__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5093__A _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5524__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5268__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6917__A _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_113_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6768__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3980_ _4751_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3980_/X sky130_fd_sc_hd__and2_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5650_ _6965_/A _5652_/A2 _5652_/B1 hold613/X vssd1 vssd1 vccd1 vccd1 _5650_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _8467_/Q _8399_/Q _8431_/Q _8305_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4601_/X sky130_fd_sc_hd__mux4_1
X_5581_ _5581_/A _7940_/Q vssd1 vssd1 vccd1 vccd1 _6704_/B sky130_fd_sc_hd__or2_4
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4532_ _4531_/X _4530_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _4532_/X sky130_fd_sc_hd__mux2_1
X_7320_ _8365_/CLK _7320_/D vssd1 vssd1 vccd1 vccd1 _7320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold326 _7324_/Q vssd1 vssd1 vccd1 vccd1 _5421_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold304 _8135_/Q vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 _5415_/X vssd1 vssd1 vccd1 vccd1 _7604_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4463_ _7028_/A _7924_/Q vssd1 vssd1 vccd1 vccd1 _8056_/D sky130_fd_sc_hd__and2_1
Xhold359 _5229_/X vssd1 vssd1 vccd1 vccd1 _7437_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold348 _8519_/Q vssd1 vssd1 vccd1 vccd1 _5549_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 _5440_/X vssd1 vssd1 vccd1 vccd1 _7629_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _5740_/B _6198_/X _6200_/X vssd1 vssd1 vccd1 vccd1 _6202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4394_ _4394_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4394_/X sky130_fd_sc_hd__and2_1
XFILLER_0_110_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6827__A _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5259__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6133_ _6309_/A _6132_/X _6131_/X vssd1 vssd1 vccd1 vccd1 _6133_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6016_/A _5993_/A _6056_/A _6035_/A _5789_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6064_/X sky130_fd_sc_hd__mux4_1
Xhold1004 _5629_/X vssd1 vssd1 vccd1 vccd1 _7809_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1015 _8148_/Q vssd1 vssd1 vccd1 vccd1 _6576_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5450__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1026 _5349_/X vssd1 vssd1 vccd1 vccd1 _7576_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1037 _7485_/Q vssd1 vssd1 vccd1 vccd1 _5281_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 _7003_/X vssd1 vssd1 vccd1 vccd1 _8461_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5015_ _5417_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5015_/X sky130_fd_sc_hd__or2_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout181_A _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout279_A _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1059 _8323_/Q vssd1 vssd1 vccd1 vccd1 _6772_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6759__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4781__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout446_A _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6966_ _7017_/A _6966_/A2 _6970_/A3 _6965_/X vssd1 vssd1 vccd1 vccd1 _6966_/X sky130_fd_sc_hd__a31o_1
X_5917_ _5891_/Y _5895_/B _5893_/B vssd1 vssd1 vccd1 vccd1 _5923_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6897_ _6963_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6897_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5848_ _5823_/A _5820_/X _5822_/B vssd1 vssd1 vccd1 vccd1 _5850_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5779_ _6035_/A _6056_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5779_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7518_ _7518_/CLK _7518_/D vssd1 vssd1 vccd1 vccd1 _7518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8498_ _8501_/CLK _8498_/D vssd1 vssd1 vccd1 vccd1 _8498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7449_ _8339_/CLK _7449_/D vssd1 vssd1 vccd1 vccd1 _7449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold882 _6762_/X vssd1 vssd1 vccd1 vccd1 _8313_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold860 _5232_/X vssd1 vssd1 vccd1 vccd1 _7440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold871 _7826_/Q vssd1 vssd1 vccd1 vccd1 hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _8457_/Q vssd1 vssd1 vccd1 vccd1 _6999_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4956__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1560 _4238_/X vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1571 _7036_/Y vssd1 vssd1 vccd1 vccd1 _7037_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1582 _4232_/X vssd1 vssd1 vccd1 vccd1 _5562_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1593 hold1822/X vssd1 vssd1 vccd1 vccd1 _5081_/A sky130_fd_sc_hd__buf_1
XFILLER_0_98_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5519__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6411__S _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6150__A1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4866__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output75_A _8102_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6647__A _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5551__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6820_ _7019_/A _6820_/A2 _6779_/B _6819_/X vssd1 vssd1 vccd1 vccd1 _6820_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_49_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6751_ _6925_/A _6741_/B _6774_/B1 hold585/X vssd1 vssd1 vccd1 vccd1 _6751_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3963_ _4067_/A_N _7943_/Q vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__and2b_1
X_5702_ _5700_/X _5701_/X _5797_/S vssd1 vssd1 vccd1 vccd1 _5702_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3894_ _3894_/A _6223_/A vssd1 vssd1 vccd1 vccd1 _3895_/B sky130_fd_sc_hd__nand2_1
X_6682_ _6931_/A _6701_/A2 _6701_/B1 hold867/X vssd1 vssd1 vccd1 vccd1 _6682_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5429__C _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8421_ _8421_/CLK _8421_/D vssd1 vssd1 vccd1 vccd1 _8421_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6064__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5716__A1 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5633_ _6931_/A _5652_/A2 _5652_/B1 hold911/X vssd1 vssd1 vccd1 vccd1 _5633_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5564_ _6545_/A _5564_/B vssd1 vssd1 vccd1 vccd1 _7753_/D sky130_fd_sc_hd__and2_1
XANTENNA__3727__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8352_ _8353_/CLK _8352_/D vssd1 vssd1 vccd1 vccd1 _8352_/Q sky130_fd_sc_hd__dfxtp_1
Xhold101 _6465_/X vssd1 vssd1 vccd1 vccd1 _7947_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4515_ _5404_/A _5404_/B vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__nand2b_4
XANTENNA__5445__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7303_ _8071_/CLK _7303_/D _7113_/Y vssd1 vssd1 vccd1 vccd1 _7303_/Q sky130_fd_sc_hd__dfrtp_4
Xhold112 _7740_/Q vssd1 vssd1 vccd1 vccd1 _6491_/B sky130_fd_sc_hd__dlygate4sd3_1
X_8283_ _8283_/CLK _8283_/D vssd1 vssd1 vccd1 vccd1 _8283_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4116__A_N _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5495_ _7516_/Q _5538_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7684_/D sky130_fd_sc_hd__and3_1
XFILLER_0_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold134 _7854_/Q vssd1 vssd1 vccd1 vccd1 _6475_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold123 _5680_/X vssd1 vssd1 vccd1 vccd1 _7860_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _7739_/Q vssd1 vssd1 vccd1 vccd1 _6490_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _5664_/X vssd1 vssd1 vccd1 vccd1 _7844_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4449_/A _4449_/B _4171_/B vssd1 vssd1 vccd1 vccd1 _4446_/X sky130_fd_sc_hd__a21o_1
Xhold167 _6476_/X vssd1 vssd1 vccd1 vccd1 _7958_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6692__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold189 _6516_/X vssd1 vssd1 vccd1 vccd1 _7998_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ _4377_/A _4377_/B vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold178 _7333_/Q vssd1 vssd1 vccd1 vccd1 _5430_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6116_ _6116_/A _6116_/B vssd1 vssd1 vccd1 vccd1 _6119_/A sky130_fd_sc_hd__nor2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7096_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7096_/Y sky130_fd_sc_hd__inv_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6008_/A _5836_/Y _5955_/Y vssd1 vssd1 vccd1 vccd1 _6047_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5652__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7998_ _8030_/CLK _7998_/D vssd1 vssd1 vccd1 vccd1 _7998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6949_ _6949_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6949_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6683__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6467__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold690 _5617_/X vssd1 vssd1 vccd1 vccd1 _7801_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4686__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5371__A _7065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4541__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5643__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1390 _4431_/X vssd1 vssd1 vccd1 vccd1 _8366_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4434__B _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4139__A_N _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3709__B1 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6910__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5174__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5280_ _6941_/A _5294_/A2 _5294_/B1 hold523/X vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4300_ _4298_/Y _4300_/B vssd1 vssd1 vccd1 vccd1 _4300_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__6674__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4596__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4231_ _4221_/Y _4225_/B _4223_/B vssd1 vssd1 vccd1 vccd1 _4231_/X sky130_fd_sc_hd__o21a_1
XANTENNA__7911__D _7911_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4780__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4162_ _5551_/B _5003_/A0 _7073_/A vssd1 vssd1 vccd1 vccd1 _4449_/B sky130_fd_sc_hd__mux2_2
X_4093_ _5772_/S _3934_/B _5804_/A vssd1 vssd1 vccd1 vccd1 _4093_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5634__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7921_ _8457_/CLK _7921_/D vssd1 vssd1 vccd1 vccd1 _7921_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7001__A _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7852_ _8019_/CLK _7852_/D vssd1 vssd1 vccd1 vccd1 _7852_/Q sky130_fd_sc_hd__dfxtp_1
X_6803_ _6935_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6803_/X sky130_fd_sc_hd__and2_1
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7783_ _8473_/CLK _7783_/D vssd1 vssd1 vccd1 vccd1 _7783_/Q sky130_fd_sc_hd__dfxtp_1
X_4995_ _4993_/X _4994_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4995_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_105_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3948__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3946_ _5763_/A _5763_/B vssd1 vssd1 vccd1 vccd1 _3946_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6734_ _6963_/A _6737_/A2 _6737_/B1 hold973/X vssd1 vssd1 vccd1 vccd1 _6734_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6665_ _6971_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6665_/X sky130_fd_sc_hd__and2_1
X_8404_ _8472_/CLK _8404_/D vssd1 vssd1 vccd1 vccd1 _8404_/Q sky130_fd_sc_hd__dfxtp_1
X_3877_ _4767_/B _4071_/A2 _4071_/B1 _3875_/X _3876_/X vssd1 vssd1 vccd1 vccd1 _6262_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_104_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6596_ _8530_/Z _5388_/X _5399_/A vssd1 vssd1 vccd1 vccd1 _6596_/Y sky130_fd_sc_hd__a21oi_1
X_5616_ _6969_/A _5616_/A2 _5616_/B1 hold947/X vssd1 vssd1 vccd1 vccd1 _5616_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout311_A _5260_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout409_A hold1729/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8335_ _8343_/CLK _8335_/D vssd1 vssd1 vccd1 vccd1 _8335_/Q sky130_fd_sc_hd__dfxtp_1
X_5547_ _7090_/A _5547_/B vssd1 vssd1 vccd1 vccd1 _7736_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4373__B1 _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5478_ _7057_/A _7073_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _7667_/D sky130_fd_sc_hd__and3_1
X_8266_ _8460_/CLK _8266_/D vssd1 vssd1 vccd1 vccd1 _8266_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4429_ _5022_/A1 _5144_/A2 _4427_/X _4428_/Y vssd1 vssd1 vccd1 vccd1 _8367_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_112_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4125__B1 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _7357_/Q vssd1 vssd1 vccd1 vccd1 _4895_/S0 sky130_fd_sc_hd__buf_8
Xfanout411 _5476_/A vssd1 vssd1 vccd1 vccd1 _4997_/S1 sky130_fd_sc_hd__buf_4
X_8197_ _8451_/CLK _8197_/D vssd1 vssd1 vccd1 vccd1 _8197_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout400 _7059_/A vssd1 vssd1 vccd1 vccd1 _4991_/S sky130_fd_sc_hd__buf_8
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout455 _6552_/A vssd1 vssd1 vccd1 vccd1 _6534_/A sky130_fd_sc_hd__clkbuf_4
Xfanout466 _6911_/A vssd1 vssd1 vccd1 vccd1 _6741_/A sky130_fd_sc_hd__buf_6
Xfanout444 _7029_/A vssd1 vssd1 vccd1 vccd1 _7019_/A sky130_fd_sc_hd__buf_4
Xfanout433 _6660_/A1 vssd1 vssd1 vccd1 vccd1 _7023_/A sky130_fd_sc_hd__buf_4
X_7079_ _7079_/A _7079_/B _7079_/C vssd1 vssd1 vccd1 vccd1 _8514_/D sky130_fd_sc_hd__and3_1
XANTENNA__6417__A2 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6968__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4523__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6050__B1 _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5156__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4270__A _8500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5085__B _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6909__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6105__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5532__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6925__A _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3890__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5616__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4780_ _8456_/Q _8388_/Q _8420_/Q _8294_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4780_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4518__C_N _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _3800_/A _3800_/B _3800_/C _3800_/D vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__or4_1
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6592__A1 _3837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3731_ _3968_/A _4307_/A vssd1 vssd1 vccd1 vccd1 _3731_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_28_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7906__D _7906_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6344__A1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6450_ _7267_/A _6450_/B vssd1 vssd1 vccd1 vccd1 _7932_/D sky130_fd_sc_hd__nor2_1
X_5401_ _6600_/A _6600_/B _5401_/C vssd1 vssd1 vccd1 vccd1 _7596_/D sky130_fd_sc_hd__and3_1
X_6381_ _6412_/S _5899_/B _6362_/C _6379_/X _6380_/Y vssd1 vssd1 vccd1 vccd1 _6381_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_3_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5332_ _6971_/A _5332_/A2 _5332_/B1 hold487/X vssd1 vssd1 vccd1 vccd1 _5332_/X sky130_fd_sc_hd__a22o_1
X_8120_ _8120_/CLK _8120_/D vssd1 vssd1 vccd1 vccd1 _8120_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6819__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5263_ _7010_/A _5263_/B vssd1 vssd1 vccd1 vccd1 _5263_/Y sky130_fd_sc_hd__nand2_1
X_8051_ _8051_/CLK _8051_/D vssd1 vssd1 vccd1 vccd1 _8051_/Q sky130_fd_sc_hd__dfxtp_1
X_4214_ _4430_/A _4430_/B vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__and2b_1
X_7002_ _7024_/A _7002_/B vssd1 vssd1 vccd1 vccd1 _7002_/X sky130_fd_sc_hd__and2_1
X_5194_ _6917_/A _5188_/B _5220_/B1 _5194_/B2 vssd1 vssd1 vccd1 vccd1 _5194_/X sky130_fd_sc_hd__a22o_1
X_4145_ _5732_/C _4148_/B _8453_/Q vssd1 vssd1 vccd1 vccd1 _4153_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__6835__A _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5607__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4076_ _4076_/A _6112_/A vssd1 vssd1 vccd1 vccd1 _4077_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout261_A _5262_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7904_ _8431_/CLK _7904_/D vssd1 vssd1 vccd1 vccd1 _7904_/Q sky130_fd_sc_hd__dfxtp_1
X_7208__86 _8479_/CLK vssd1 vssd1 vccd1 vccd1 _8121_/CLK sky130_fd_sc_hd__inv_2
X_7835_ _8456_/CLK _7835_/D vssd1 vssd1 vccd1 vccd1 _7835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7766_ _8494_/CLK _7766_/D vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
X_4978_ _4977_/X _4974_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8258_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_46_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6583__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6717_ _6929_/A _6705_/B _6738_/B1 hold427/X vssd1 vssd1 vccd1 vccd1 _6717_/X sky130_fd_sc_hd__a22o_1
X_3929_ _4014_/A _6421_/B _3927_/Y vssd1 vssd1 vccd1 vccd1 _5716_/S sky130_fd_sc_hd__o21ai_4
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7697_ _8463_/CLK _7697_/D vssd1 vssd1 vccd1 vccd1 _7697_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5138__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6648_ _7025_/A _6648_/A2 _6666_/A3 _6647_/X vssd1 vssd1 vccd1 vccd1 _6648_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_116_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8318_ _8460_/CLK _8318_/D vssd1 vssd1 vccd1 vccd1 _8318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6579_ _6945_/A _6559_/B _6591_/B1 hold987/X vssd1 vssd1 vccd1 vccd1 _6579_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_131_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6099__A0 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8249_ _8249_/CLK _8249_/D vssd1 vssd1 vccd1 vccd1 _8249_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5310__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout230 _5451_/C vssd1 vssd1 vccd1 vccd1 _5453_/C sky130_fd_sc_hd__buf_4
Xfanout241 _5099_/B vssd1 vssd1 vccd1 vccd1 _5144_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout274 _3669_/Y vssd1 vssd1 vccd1 vccd1 _3676_/A sky130_fd_sc_hd__buf_12
Xfanout252 _6559_/Y vssd1 vssd1 vccd1 vccd1 _6592_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout263 _5226_/Y vssd1 vssd1 vccd1 vccd1 _5258_/B1 sky130_fd_sc_hd__buf_6
XANTENNA__4964__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout296 _6601_/Y vssd1 vssd1 vccd1 vccd1 _6661_/B sky130_fd_sc_hd__buf_8
Xfanout285 _6775_/Y vssd1 vssd1 vccd1 vccd1 _6837_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__5074__A1 input28/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6911__C _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5527__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6639__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4983__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5543__B _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6655__A _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3863__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5950_ _5831_/X _5834_/B _5950_/S vssd1 vssd1 vccd1 vccd1 _5951_/B sky130_fd_sc_hd__mux2_1
X_4901_ _4900_/X _4897_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8247_/D sky130_fd_sc_hd__mux2_1
X_5881_ _6008_/A _6307_/A _5881_/C _6362_/B vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__or4_1
X_7620_ _8090_/CLK _7620_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_118_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4832_ _8334_/Q _7810_/Q _7476_/Q _7444_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4832_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5368__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6565__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7551_ _8445_/CLK _7551_/D vssd1 vssd1 vccd1 vccd1 _7551_/Q sky130_fd_sc_hd__dfxtp_1
X_4763_ _7017_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _8120_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4671__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6502_ _6548_/A hold9/X vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__and2_1
X_7482_ _8413_/CLK _7482_/D vssd1 vssd1 vccd1 vccd1 _7482_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5437__C _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3714_ _3714_/A _3714_/B vssd1 vssd1 vccd1 vccd1 _3750_/A sky130_fd_sc_hd__and2_1
XFILLER_0_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4694_ _4693_/X _4690_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7524_/D sky130_fd_sc_hd__mux2_1
X_6433_ _6706_/A _6433_/B vssd1 vssd1 vccd1 vccd1 _7915_/D sky130_fd_sc_hd__and2_1
XFILLER_0_113_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5734__A _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6364_ _3848_/B _6414_/A2 _6130_/A _6361_/Y _6362_/X vssd1 vssd1 vccd1 vccd1 _6364_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5453__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8103_ _8103_/CLK _8103_/D vssd1 vssd1 vccd1 vccd1 _8103_/Q sky130_fd_sc_hd__dfxtp_2
X_5315_ _6937_/A _5332_/A2 _5332_/B1 hold907/X vssd1 vssd1 vccd1 vccd1 _5315_/X sky130_fd_sc_hd__a22o_1
X_6295_ _6295_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6298_/B sky130_fd_sc_hd__xnor2_1
X_7124__2 _8388_/CLK vssd1 vssd1 vccd1 vccd1 _7501_/CLK sky130_fd_sc_hd__inv_2
X_8034_ _8034_/CLK _8034_/D vssd1 vssd1 vccd1 vccd1 _8034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5246_ _6945_/A _5258_/A2 _5258_/B1 hold481/X vssd1 vssd1 vccd1 vccd1 _5246_/X sky130_fd_sc_hd__a22o_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4726__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _5468_/A _5468_/C vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__or2_1
X_4128_ _4122_/Y _4127_/X _3897_/D vssd1 vssd1 vccd1 vccd1 _4128_/X sky130_fd_sc_hd__a21o_1
X_4059_ _4059_/A1 _4084_/A2 _6933_/A _4084_/B2 _4058_/X vssd1 vssd1 vccd1 vccd1 _4059_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1493_A _7313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7818_ _8445_/CLK _7818_/D vssd1 vssd1 vccd1 vccd1 _7818_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5359__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7749_ _8079_/CLK _7749_/D vssd1 vssd1 vccd1 vccd1 _7749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4024__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3790__B2 _8022_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4965__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5295__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4717__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4694__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6475__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5598__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7199__77 _8086_/CLK vssd1 vssd1 vccd1 vccd1 _8112_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4442__B _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5538__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4653__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5770__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4869__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5554__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3781__B2 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 _5612_/X vssd1 vssd1 vccd1 vccd1 _7796_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold519 _7498_/Q vssd1 vssd1 vccd1 vccd1 hold519/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6080_ _6144_/S _6080_/B vssd1 vssd1 vccd1 vccd1 _6080_/X sky130_fd_sc_hd__or2_1
X_5100_ input11/X _5099_/B _5002_/X _5099_/Y vssd1 vssd1 vccd1 vccd1 _7362_/D sky130_fd_sc_hd__o211a_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5905__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5286__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5031_ _5425_/A _5454_/C vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__or2_1
Xhold1208 _6840_/X vssd1 vssd1 vccd1 vccd1 _8357_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1219 _8173_/Q vssd1 vssd1 vccd1 vccd1 _6618_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5589__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6982_ _5382_/X _6595_/A _6980_/X _6981_/Y vssd1 vssd1 vccd1 vccd1 _6982_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_76_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6786__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5933_ _3962_/X _6105_/A2 _5931_/X _5932_/X vssd1 vssd1 vccd1 vccd1 _5933_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_88_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4892__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5864_ _6163_/A _5842_/X _5851_/Y _5863_/X vssd1 vssd1 vccd1 vccd1 _5864_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6324__S _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5448__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4815_ _8461_/Q _8393_/Q _8425_/Q _8299_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4815_/X sky130_fd_sc_hd__mux4_1
X_7603_ _8360_/CLK _7603_/D vssd1 vssd1 vccd1 vccd1 _7603_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7534_ _8136_/CLK _7534_/D vssd1 vssd1 vccd1 vccd1 _7534_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4013__A2 _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5795_ _5921_/A _5946_/A _5974_/A _5993_/A _5744_/S _5797_/S vssd1 vssd1 vccd1 vccd1
+ _5795_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5210__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout224_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4746_ _7029_/A _4746_/B vssd1 vssd1 vccd1 vccd1 _8103_/D sky130_fd_sc_hd__and2_1
XFILLER_0_126_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3683__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4677_ _8188_/Q _8220_/Q _8284_/Q _7792_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4677_/X sky130_fd_sc_hd__mux4_1
X_7465_ _8355_/CLK _7465_/D vssd1 vssd1 vccd1 vccd1 _7465_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6710__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6416_ _6416_/A _6416_/B vssd1 vssd1 vccd1 vccd1 _6416_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6279__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4947__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7396_ _8382_/CLK _7396_/D vssd1 vssd1 vccd1 vccd1 _7396_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6347_ _3749_/B _6292_/A _6347_/B1 vssd1 vssd1 vccd1 vccd1 _6347_/Y sky130_fd_sc_hd__a21oi_1
X_6278_ _6261_/Y _6266_/B _6263_/B vssd1 vssd1 vccd1 vccd1 _6283_/A sky130_fd_sc_hd__a21o_1
X_5229_ _3939_/C _5227_/B _5227_/Y hold358/X vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__o22a_1
X_8017_ _8370_/CLK _8017_/D vssd1 vssd1 vccd1 vccd1 _8017_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3712__A _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1720 _8499_/Q vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__buf_1
XFILLER_0_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1731 _8165_/Q vssd1 vssd1 vccd1 vccd1 _5730_/A sky130_fd_sc_hd__clkbuf_2
Xhold1753 _8455_/Q vssd1 vssd1 vccd1 vccd1 _5738_/A sky130_fd_sc_hd__clkbuf_2
Xhold1742 _7729_/Q vssd1 vssd1 vccd1 vccd1 _3827_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1764 _7712_/Q vssd1 vssd1 vccd1 vccd1 _4062_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1775 _7707_/Q vssd1 vssd1 vccd1 vccd1 _3978_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1786 _6262_/A vssd1 vssd1 vccd1 vccd1 _3882_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1797 _7876_/Q vssd1 vssd1 vccd1 vccd1 hold1797/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4252__A2 _4246_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4022__A_N _7283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4004__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4635__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5201__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6701__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4938__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5268__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6917__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4437__B _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6768__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5549__A _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4874__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4515__A_N _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4600_ _8177_/Q _8209_/Q _8273_/Q _7781_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4600_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4626__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5580_ _6520_/A _5580_/B vssd1 vssd1 vccd1 vccd1 _7769_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6940__A1 _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4531_ _8457_/Q _8389_/Q _8421_/Q _8295_/Q _7362_/Q _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4531_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3754__A1 _3753_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4599__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4462_ _6999_/A _7925_/Q vssd1 vssd1 vccd1 vccd1 _8057_/D sky130_fd_sc_hd__and2_1
Xhold305 _6563_/X vssd1 vssd1 vccd1 vccd1 _8135_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold316 _7328_/Q vssd1 vssd1 vccd1 vccd1 _5425_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 _5421_/X vssd1 vssd1 vccd1 vccd1 _7610_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _7325_/Q vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 _5549_/X vssd1 vssd1 vccd1 vccd1 _7738_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _6309_/A _5837_/X _6130_/A vssd1 vssd1 vccd1 vccd1 _6201_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4393_ _5046_/A1 _4392_/Y _5454_/C vssd1 vssd1 vccd1 vccd1 _4393_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5259__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6132_ _5951_/B _5964_/X _6411_/S vssd1 vssd1 vccd1 vccd1 _6132_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6827__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ _6063_/A _6063_/B _6063_/C vssd1 vssd1 vccd1 vccd1 _6063_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_84_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1005 _8467_/Q vssd1 vssd1 vccd1 vccd1 _7009_/B sky130_fd_sc_hd__dlygate4sd3_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7004__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1038 _5281_/X vssd1 vssd1 vccd1 vccd1 _7485_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ _4437_/A _4448_/B _5140_/B1 _5013_/X vssd1 vssd1 vccd1 vccd1 _7319_/D sky130_fd_sc_hd__o211a_1
Xhold1016 _6576_/X vssd1 vssd1 vccd1 vccd1 _8148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 _7472_/Q vssd1 vssd1 vccd1 vccd1 _5268_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 _8153_/Q vssd1 vssd1 vccd1 vccd1 _6581_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6843__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout174_A hold1510/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6303__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6759__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ _6965_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6965_/X sky130_fd_sc_hd__and2_1
XANTENNA__4363__A _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5916_ _5916_/A1 _6011_/A2 _5914_/Y _5915_/X _6911_/A vssd1 vssd1 vccd1 vccd1 _7873_/D
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_88_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3993__A1 _6426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6896_ _7024_/A _6896_/A2 _6845_/B _6895_/X vssd1 vssd1 vccd1 vccd1 _6896_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout439_A _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5847_ _5847_/A _5847_/B vssd1 vssd1 vccd1 vccd1 _5850_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5195__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5778_ _5776_/X _5777_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7517_ _7517_/CLK _7517_/D vssd1 vssd1 vccd1 vccd1 _7517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8497_ _8501_/CLK _8497_/D vssd1 vssd1 vccd1 vccd1 _8497_/Q sky130_fd_sc_hd__dfxtp_1
X_4729_ _4728_/X _4725_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7529_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7448_ _8332_/CLK _7448_/D vssd1 vssd1 vccd1 vccd1 _7448_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_110_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8479_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6695__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7243__121 _8486_/CLK vssd1 vssd1 vccd1 vccd1 _8253_/CLK sky130_fd_sc_hd__inv_2
X_7379_ _8358_/CLK _7379_/D vssd1 vssd1 vccd1 vccd1 _7379_/Q sky130_fd_sc_hd__dfxtp_1
Xhold861 _7499_/Q vssd1 vssd1 vccd1 vccd1 hold861/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold850 _5212_/X vssd1 vssd1 vccd1 vccd1 _7426_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 _5646_/X vssd1 vssd1 vccd1 vccd1 _7826_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _6999_/X vssd1 vssd1 vccd1 vccd1 _8457_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _7881_/Q vssd1 vssd1 vccd1 vccd1 hold883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 _4239_/X vssd1 vssd1 vccd1 vccd1 _5563_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1550 _8437_/Q vssd1 vssd1 vccd1 vccd1 _6943_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 _7368_/Q vssd1 vssd1 vccd1 vccd1 _7078_/A sky130_fd_sc_hd__clkbuf_4
Xhold1594 _7684_/Q vssd1 vssd1 vccd1 vccd1 _3756_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1572 _7647_/Q vssd1 vssd1 vccd1 vccd1 _4271_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5369__A _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4856__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7169__47 _8010_/CLK vssd1 vssd1 vccd1 vccd1 _8049_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4608__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6922__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_101_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _8173_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_50_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6686__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6150__A2 _5719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6647__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6438__B1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5110__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6663__A _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4847__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6750_ _6923_/A _6773_/A2 _6773_/B1 hold817/X vssd1 vssd1 vccd1 vccd1 _6750_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_128_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3962_ _3962_/A _3962_/B vssd1 vssd1 vccd1 vccd1 _3962_/X sky130_fd_sc_hd__and2_1
X_5701_ _6096_/A _6115_/A _5744_/S vssd1 vssd1 vccd1 vccd1 _5701_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6681_ _6929_/A _6669_/B _6702_/B1 hold370/X vssd1 vssd1 vccd1 vccd1 _6681_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3893_ _6226_/A _6223_/A vssd1 vssd1 vccd1 vccd1 _3895_/A sky130_fd_sc_hd__or2_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8420_ _8421_/CLK _8420_/D vssd1 vssd1 vccd1 vccd1 _8420_/Q sky130_fd_sc_hd__dfxtp_1
X_5632_ _6929_/A _5620_/B _5653_/B1 hold533/X vssd1 vssd1 vccd1 vccd1 _5632_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5563_ _6534_/A _5563_/B vssd1 vssd1 vccd1 vccd1 _7752_/D sky130_fd_sc_hd__and2_1
X_8351_ _8451_/CLK _8351_/D vssd1 vssd1 vccd1 vccd1 _8351_/Q sky130_fd_sc_hd__dfxtp_1
X_7227__105 _8173_/CLK vssd1 vssd1 vccd1 vccd1 _8237_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4514_ _5124_/A1 _4449_/B _7082_/B vssd1 vssd1 vccd1 vccd1 _7284_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_53_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7183__61 _8476_/CLK vssd1 vssd1 vccd1 vccd1 _8063_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7302_ _8378_/CLK _7302_/D _7112_/Y vssd1 vssd1 vccd1 vccd1 _7302_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6677__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold124 _7752_/Q vssd1 vssd1 vccd1 vccd1 _6503_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _6491_/X vssd1 vssd1 vccd1 vccd1 _7973_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _7600_/Q vssd1 vssd1 vccd1 vccd1 _5658_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _6475_/X vssd1 vssd1 vccd1 vccd1 _7957_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5494_ _7515_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7683_/D sky130_fd_sc_hd__and3_1
XFILLER_0_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8282_ _8440_/CLK _8282_/D vssd1 vssd1 vccd1 vccd1 _8282_/Q sky130_fd_sc_hd__dfxtp_1
Xhold157 _6490_/X vssd1 vssd1 vccd1 vccd1 _7972_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _7748_/Q vssd1 vssd1 vccd1 vccd1 _6499_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4445_/A _5069_/S vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__and2_1
Xhold146 _7841_/Q vssd1 vssd1 vccd1 vccd1 _6462_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4376_ _5060_/A1 _5069_/S _4371_/Y _4375_/X vssd1 vssd1 vccd1 vccd1 _8386_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold179 _5430_/X vssd1 vssd1 vccd1 vccd1 _7619_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6115_ _6115_/A _6115_/B vssd1 vssd1 vccd1 vccd1 _6116_/B sky130_fd_sc_hd__nor2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7095_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7095_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout389_A _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout291_A _6667_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6046_ _6105_/A2 _6038_/A _6044_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6046_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6090__A1_N _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5652__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4792__S _7359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_54_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5189__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7997_ _8385_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 _7997_/Q sky130_fd_sc_hd__dfxtp_1
X_6948_ _7017_/A _6948_/A2 _6970_/A3 _6947_/X vssd1 vssd1 vccd1 vccd1 _6948_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6879_ _6945_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6879_/X sky130_fd_sc_hd__and2_1
XFILLER_0_134_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_69_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6904__A1 _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5168__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_112_clk_A clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4967__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold680 _5288_/X vssd1 vssd1 vccd1 vccd1 _7492_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 _8202_/Q vssd1 vssd1 vccd1 vccd1 hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5643__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5798__S _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6483__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1391 hold1804/X vssd1 vssd1 vccd1 vccd1 _4745_/B sky130_fd_sc_hd__buf_1
Xhold1380 _8179_/Q vssd1 vssd1 vccd1 vccd1 _6630_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6199__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4829__S0 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5099__A _7052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5546__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4230_ _4228_/Y _4230_/B vssd1 vssd1 vccd1 vccd1 _4232_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__5331__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4161_ _4161_/A _4161_/B vssd1 vssd1 vccd1 vccd1 _5551_/B sky130_fd_sc_hd__xor2_1
X_4092_ _4092_/A _4092_/B _4092_/C _4092_/D vssd1 vssd1 vccd1 vccd1 _4152_/A sky130_fd_sc_hd__or4_2
X_7920_ _8457_/CLK _7920_/D vssd1 vssd1 vccd1 vccd1 _7920_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6393__A _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3810__A _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7851_ _8019_/CLK hold78/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfxtp_1
X_6802_ _7010_/A _6802_/A2 _6779_/B _6801_/X vssd1 vssd1 vccd1 vccd1 _6802_/X sky130_fd_sc_hd__a31o_1
X_7782_ _8466_/CLK _7782_/D vssd1 vssd1 vccd1 vccd1 _7782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4994_ _8164_/Q _7563_/Q _7435_/Q _7595_/Q _5475_/A _4997_/S1 vssd1 vssd1 vccd1 vccd1
+ _4994_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3948__B2 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3945_ _5763_/A _5763_/B vssd1 vssd1 vccd1 vccd1 _3945_/Y sky130_fd_sc_hd__nor2_1
X_6733_ _6961_/A _6737_/A2 _6737_/B1 hold555/X vssd1 vssd1 vccd1 vccd1 _6733_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6664_ _7026_/A _6664_/A2 _6666_/A3 _6663_/X vssd1 vssd1 vccd1 vccd1 _6664_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5615_ _6967_/A _5616_/A2 _5616_/B1 _5615_/B2 vssd1 vssd1 vccd1 vccd1 _5615_/X sky130_fd_sc_hd__a22o_1
X_8403_ _8471_/CLK _8403_/D vssd1 vssd1 vccd1 vccd1 _8403_/Q sky130_fd_sc_hd__dfxtp_1
X_3876_ _3876_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3876_/X sky130_fd_sc_hd__or2_1
XFILLER_0_104_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6595_ _6595_/A vssd1 vssd1 vccd1 vccd1 _6595_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout304_A _5618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5546_ _5546_/A _7088_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _7735_/D sky130_fd_sc_hd__and3_1
X_8334_ _8428_/CLK _8334_/D vssd1 vssd1 vccd1 vccd1 _8334_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5477_ _5477_/A _7088_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _7666_/D sky130_fd_sc_hd__and3_1
X_8265_ _8338_/CLK _8265_/D vssd1 vssd1 vccd1 vccd1 _8265_/Q sky130_fd_sc_hd__dfxtp_1
X_4428_ _4427_/A _4427_/B _4425_/B vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5472__A _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5322__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout412 _5476_/A vssd1 vssd1 vccd1 vccd1 _4896_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout423 _7357_/Q vssd1 vssd1 vccd1 vccd1 _4896_/S0 sky130_fd_sc_hd__buf_4
Xfanout401 _7059_/A vssd1 vssd1 vccd1 vccd1 _4988_/S sky130_fd_sc_hd__buf_4
X_8196_ _8442_/CLK _8196_/D vssd1 vssd1 vccd1 vccd1 _8196_/Q sky130_fd_sc_hd__dfxtp_1
X_4359_ _5472_/A _7733_/Q vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__xnor2_1
Xfanout456 _6552_/A vssd1 vssd1 vccd1 vccd1 _6548_/A sky130_fd_sc_hd__clkbuf_2
Xfanout445 _7029_/A vssd1 vssd1 vccd1 vccd1 _7015_/A sky130_fd_sc_hd__clkbuf_4
Xfanout434 _6660_/A1 vssd1 vssd1 vccd1 vccd1 _7026_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7078_ _7078_/A _7079_/B _7079_/C vssd1 vssd1 vccd1 vccd1 _8513_/D sky130_fd_sc_hd__and3_1
Xfanout467 input63/X vssd1 vssd1 vccd1 vccd1 _6911_/A sky130_fd_sc_hd__buf_6
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5625__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6029_ _5694_/Y _6028_/X _6027_/Y _6083_/A vssd1 vssd1 vccd1 vccd1 _6029_/X sky130_fd_sc_hd__o2bb2a_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3720__A _4770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7139__17 _8445_/CLK vssd1 vssd1 vccd1 vccd1 _7516_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6105__A2 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4697__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6478__A _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5313__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5864__A1 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6656__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7066__B1 _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6925__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5616__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7102__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4106__A_N _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4445__B _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6941__A _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__B1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5557__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6592__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3730_ _4768_/B _4072_/B _3730_/B1 vssd1 vssd1 vccd1 vccd1 _6445_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _7666_/Q vssd1 vssd1 vccd1 vccd1 _3661_/Y sky130_fd_sc_hd__inv_2
X_5400_ _8531_/Z _6976_/A _5399_/Y _5382_/X _6597_/B vssd1 vssd1 vccd1 vccd1 _5401_/C
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6380_ _6380_/A _6380_/B vssd1 vssd1 vccd1 vccd1 _6380_/Y sky130_fd_sc_hd__nor2_1
X_7153__31 _8484_/CLK vssd1 vssd1 vccd1 vccd1 _7530_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6388__A _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5331_ _6969_/A _5299_/B _5331_/B1 hold531/X vssd1 vssd1 vccd1 vccd1 _5331_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4107__B2 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8050_ _8050_/CLK _8050_/D vssd1 vssd1 vccd1 vccd1 _8050_/Q sky130_fd_sc_hd__dfxtp_1
X_7001_ _7010_/A _7001_/B vssd1 vssd1 vccd1 vccd1 _7001_/X sky130_fd_sc_hd__and2_1
XANTENNA__5855__A1 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5262_ _7267_/A _5262_/B vssd1 vssd1 vccd1 vccd1 _5262_/Y sky130_fd_sc_hd__nor2_2
X_5193_ _6849_/A _5189_/B _5189_/Y hold284/X vssd1 vssd1 vccd1 vccd1 _5193_/X sky130_fd_sc_hd__o22a_1
X_4213_ _4212_/X _5020_/A1 _5453_/B vssd1 vssd1 vccd1 vccd1 _4430_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5855__B2 _5739_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4144_ _8454_/Q _4144_/B vssd1 vssd1 vccd1 vccd1 _4144_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5607__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6835__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7012__A _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4075_ _6115_/A _6112_/A vssd1 vssd1 vccd1 vccd1 _4077_/A sky130_fd_sc_hd__or2_1
X_7903_ _7903_/CLK _7903_/D vssd1 vssd1 vccd1 vccd1 _7903_/Q sky130_fd_sc_hd__dfxtp_1
X_7834_ _8079_/CLK _7834_/D vssd1 vssd1 vccd1 vccd1 _7834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout254_A _5620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6851__A _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_90_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _8378_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7765_ _8030_/CLK _7765_/D vssd1 vssd1 vccd1 vccd1 _7765_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6716_ _6927_/A _6705_/B _6738_/B1 hold551/X vssd1 vssd1 vccd1 vccd1 _6716_/X sky130_fd_sc_hd__a22o_1
X_4977_ _4976_/X _4975_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6583__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3928_ _4014_/A _6421_/B _3927_/Y vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__o21a_2
XANTENNA_fanout421_A _7357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7696_ _8419_/CLK _7696_/D vssd1 vssd1 vccd1 vccd1 _7696_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3859_ _3859_/A _3859_/B vssd1 vssd1 vccd1 vccd1 _3896_/A sky130_fd_sc_hd__and2_1
X_6647_ _6953_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6647_/X sky130_fd_sc_hd__and2_1
XFILLER_0_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6886__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6578_ _6877_/A _6592_/A2 _6592_/B1 hold981/X vssd1 vssd1 vccd1 vccd1 _6578_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8317_ _8476_/CLK _8317_/D vssd1 vssd1 vccd1 vccd1 _8317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5529_ _8248_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7718_/D sky130_fd_sc_hd__and3_1
XFILLER_0_131_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6099__A1 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6298__A _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6638__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8248_ _8248_/CLK _8248_/D vssd1 vssd1 vccd1 vccd1 _8248_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout231 _7073_/B vssd1 vssd1 vccd1 vccd1 _5451_/C sky130_fd_sc_hd__clkbuf_4
X_8179_ _8328_/CLK _8179_/D vssd1 vssd1 vccd1 vccd1 _8179_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout220 _5470_/C vssd1 vssd1 vccd1 vccd1 _5468_/C sky130_fd_sc_hd__buf_4
Xfanout242 _4369_/Y vssd1 vssd1 vccd1 vccd1 _5099_/B sky130_fd_sc_hd__buf_12
XANTENNA_hold1703_A _6422_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout264 _5226_/Y vssd1 vssd1 vccd1 vccd1 _5259_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout253 _5620_/Y vssd1 vssd1 vccd1 vccd1 _5652_/B1 sky130_fd_sc_hd__buf_6
Xfanout286 _6775_/Y vssd1 vssd1 vccd1 vccd1 _6839_/B sky130_fd_sc_hd__buf_4
Xfanout297 _6557_/Y vssd1 vssd1 vccd1 vccd1 _6559_/B sky130_fd_sc_hd__buf_6
XANTENNA__4129__A_N _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout275 _6943_/B vssd1 vssd1 vccd1 vccd1 _6970_/A3 sky130_fd_sc_hd__buf_8
XANTENNA__5074__A2 _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6271__A1 _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6810__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _8385_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6574__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4034__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6326__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4220__S _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7039__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6655__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4456__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5696__S0 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4900_ _4899_/X _4898_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4900_/X sky130_fd_sc_hd__mux2_1
X_5880_ _5702_/X _5707_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5880_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4890__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_72_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _8513_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4831_ _4830_/X _4827_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8237_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6565__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4762_ _7005_/A _4762_/B vssd1 vssd1 vccd1 vccd1 _8119_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7550_ _8218_/CLK _7550_/D vssd1 vssd1 vccd1 vccd1 _7550_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4671__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6501_ _6534_/A hold96/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__and2_1
X_7481_ _8339_/CLK _7481_/D vssd1 vssd1 vccd1 vccd1 _7481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3713_ _6298_/A _6295_/A vssd1 vssd1 vccd1 vccd1 _3714_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4693_ _4692_/X _4691_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6868__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6432_ _7015_/A _6432_/B vssd1 vssd1 vccd1 vccd1 _7914_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5734__B _6380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7007__A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8102_ _8102_/CLK _8102_/D vssd1 vssd1 vccd1 vccd1 _8102_/Q sky130_fd_sc_hd__dfxtp_1
X_6363_ _3823_/A _6414_/B1 _6398_/B1 _6350_/A _5734_/X vssd1 vssd1 vccd1 vccd1 _6363_/X
+ sky130_fd_sc_hd__a221o_1
X_5314_ _6935_/A _5332_/A2 _5332_/B1 hold915/X vssd1 vssd1 vccd1 vccd1 _5314_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_87_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6294_ _6294_/A1 _6292_/A _6293_/X _6347_/B1 vssd1 vssd1 vccd1 vccd1 _7892_/D sky130_fd_sc_hd__a211oi_1
X_5245_ _6877_/A _5226_/B _5259_/B1 hold927/X vssd1 vssd1 vccd1 vccd1 _5245_/X sky130_fd_sc_hd__a22o_1
X_8033_ _8033_/CLK _8033_/D vssd1 vssd1 vccd1 vccd1 _8033_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3839__B1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _5176_/A1 _5069_/S _5182_/B1 _5175_/X vssd1 vssd1 vccd1 vccd1 _7400_/D sky130_fd_sc_hd__o211a_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4366__A _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout469_A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6253__A1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5056__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4127_ _4123_/Y _4126_/Y _3800_/D vssd1 vssd1 vccd1 vccd1 _4127_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout371_A _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4058_ _4756_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _4058_/X sky130_fd_sc_hd__and2_1
XFILLER_0_97_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_63_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _8510_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7817_ _8218_/CLK _7817_/D vssd1 vssd1 vccd1 vccd1 _7817_/Q sky130_fd_sc_hd__dfxtp_1
X_7748_ _8510_/CLK _7748_/D vssd1 vssd1 vccd1 vccd1 _7748_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5764__B1 _5971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7679_ _8319_/CLK _7679_/D vssd1 vssd1 vccd1 vccd1 _7679_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6308__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5925__A _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1653_A _7346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3790__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4040__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5295__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5660__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6491__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_54_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _7907_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5819__B _5971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5538__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4653__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5835__A _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold509 _8310_/Q vssd1 vssd1 vccd1 vccd1 hold509/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3781__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output98_A _7293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5905__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5030_/A1 _4416_/B _5166_/B1 _5029_/X vssd1 vssd1 vccd1 vccd1 _7327_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5570__A _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5286__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1209 _8410_/Q vssd1 vssd1 vccd1 vccd1 _6888_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_6981_ _6981_/A _6981_/B vssd1 vssd1 vccd1 vccd1 _6981_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5932_ _3962_/A _6398_/A2 _6413_/B1 _5918_/A _6011_/A2 vssd1 vssd1 vccd1 vccd1 _5932_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5863_ _6198_/S _5694_/Y _5862_/X _5855_/X _5854_/X vssd1 vssd1 vccd1 vccd1 _5863_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_75_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4892__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _8171_/Q _8203_/Q _8267_/Q _7775_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4814_/X sky130_fd_sc_hd__mux4_1
X_5794_ _5846_/A _5820_/A _5892_/A _5870_/A _5772_/S _5797_/S vssd1 vssd1 vccd1 vccd1
+ _5794_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5746__A0 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7602_ _8387_/CLK _7602_/D vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__dfxtp_1
X_7533_ _8428_/CLK _7533_/D vssd1 vssd1 vccd1 vccd1 _7533_/Q sky130_fd_sc_hd__dfxtp_1
X_4745_ _7006_/A _4745_/B vssd1 vssd1 vccd1 vccd1 _8102_/D sky130_fd_sc_hd__and2_1
XFILLER_0_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5210__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7464_ _8354_/CLK _7464_/D vssd1 vssd1 vccd1 vccd1 _7464_/Q sky130_fd_sc_hd__dfxtp_1
X_4676_ _4674_/X _4675_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4676_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout217_A _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6710__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6415_ _5953_/B _6309_/Y _6412_/X _5740_/B vssd1 vssd1 vccd1 vccd1 _6416_/B sky130_fd_sc_hd__a22o_1
X_7395_ _8379_/CLK _7395_/D vssd1 vssd1 vccd1 vccd1 _7395_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5464__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6346_ _5840_/Y _6309_/Y _6338_/A _6414_/A2 _6345_/X vssd1 vssd1 vccd1 vccd1 _6346_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4795__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8016_ _8034_/CLK _8016_/D vssd1 vssd1 vccd1 vccd1 _8016_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5277__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6277_ _6267_/Y _6274_/X _6275_/X _6276_/Y vssd1 vssd1 vccd1 vccd1 _6277_/X sky130_fd_sc_hd__o31a_1
X_5228_ _6777_/A _5227_/B _5227_/Y hold334/X vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__o22a_1
Xhold1710 _8454_/Q vssd1 vssd1 vccd1 vccd1 _4148_/B sky130_fd_sc_hd__buf_1
XANTENNA__6295__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4580__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1732 _5725_/X vssd1 vssd1 vccd1 vccd1 _6030_/A1 sky130_fd_sc_hd__clkbuf_2
Xhold1743 _7716_/Q vssd1 vssd1 vccd1 vccd1 _3760_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1721 _4281_/X vssd1 vssd1 vccd1 vccd1 _5569_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5159_ _5459_/A _5454_/C vssd1 vssd1 vccd1 vccd1 _5159_/X sky130_fd_sc_hd__or2_1
Xhold1754 _5942_/Y vssd1 vssd1 vccd1 vccd1 _7874_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1765 _6056_/A vssd1 vssd1 vccd1 vccd1 _4065_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1776 _7713_/Q vssd1 vssd1 vccd1 vccd1 _4081_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1787 _6277_/X vssd1 vssd1 vccd1 vccd1 _7891_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1798 _7895_/Q vssd1 vssd1 vccd1 vccd1 hold1798/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_36_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _8468_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4035__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4635__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5201__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5655__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6701__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6486__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5268__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6933__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6768__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_27_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8175_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__7110__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4874__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4626__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3784__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4530_ _8167_/Q _8199_/Q _8263_/Q _7771_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4530_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4461_ _7022_/A _7926_/Q vssd1 vssd1 vccd1 vccd1 _8058_/D sky130_fd_sc_hd__and2_1
Xhold317 _5425_/X vssd1 vssd1 vccd1 vccd1 _7614_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold306 _7396_/Q vssd1 vssd1 vccd1 vccd1 _5463_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold339 _5422_/X vssd1 vssd1 vccd1 vccd1 _7611_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _7402_/Q vssd1 vssd1 vccd1 vccd1 _5469_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6200_ _5841_/X _6130_/B _6194_/A _6414_/A2 _6199_/X vssd1 vssd1 vccd1 vccd1 _6200_/X
+ sky130_fd_sc_hd__a221o_1
X_6131_ _5953_/B _6362_/C _6130_/X vssd1 vssd1 vccd1 vccd1 _6131_/X sky130_fd_sc_hd__a21o_1
X_4392_ _4392_/A _4392_/B vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__xnor2_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5259__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7930__D _7930_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _4090_/B _6105_/A2 _6060_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _6063_/C sky130_fd_sc_hd__a22o_1
Xhold1006 _7009_/X vssd1 vssd1 vccd1 vccd1 _8467_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1039 _7572_/Q vssd1 vssd1 vccd1 vccd1 _5345_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5013_ _5416_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__or2_1
Xhold1017 _7433_/Q vssd1 vssd1 vccd1 vccd1 _5219_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1028 _6581_/X vssd1 vssd1 vccd1 vccd1 _8153_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3959__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6759__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6303__S1 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8154_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout167_A hold1510/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6964_ _7024_/A _6964_/A2 _6943_/B _6963_/X vssd1 vssd1 vccd1 vccd1 _6964_/X sky130_fd_sc_hd__a31o_1
XANTENNA__7020__A _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5915_ _5734_/A _5895_/X _5912_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _5915_/X sky130_fd_sc_hd__o22a_1
X_6895_ _6961_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6895_/X sky130_fd_sc_hd__and2_1
XANTENNA__5459__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5846_ _5846_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5847_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_64_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5475__A _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5195__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5777_ _5921_/A _5892_/A _5974_/A _5946_/A _5782_/S _5797_/S vssd1 vssd1 vccd1 vccd1
+ _5777_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6392__A0 _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7516_ _7516_/CLK _7516_/D vssd1 vssd1 vccd1 vccd1 _7516_/Q sky130_fd_sc_hd__dfxtp_1
X_8496_ _8501_/CLK _8496_/D vssd1 vssd1 vccd1 vccd1 _8496_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4728_ _4727_/X _4726_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3707__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4659_ _4658_/X _4655_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7519_/D sky130_fd_sc_hd__mux2_1
X_7447_ _8467_/CLK _7447_/D vssd1 vssd1 vccd1 vccd1 _7447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6695__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold873 _7444_/Q vssd1 vssd1 vccd1 vccd1 hold873/X sky130_fd_sc_hd__dlygate4sd3_1
X_7378_ _8362_/CLK _7378_/D vssd1 vssd1 vccd1 vccd1 _7378_/Q sky130_fd_sc_hd__dfxtp_1
Xhold862 _5295_/X vssd1 vssd1 vccd1 vccd1 _7499_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _8144_/Q vssd1 vssd1 vccd1 vccd1 hold851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold840 _6689_/X vssd1 vssd1 vccd1 vccd1 _8216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 _6454_/X vssd1 vssd1 vccd1 vccd1 _7936_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ _6391_/A _6320_/Y _6321_/X _6412_/S _6328_/Y vssd1 vssd1 vccd1 vccd1 _6329_/X
+ sky130_fd_sc_hd__o221a_1
Xhold895 _8485_/Q vssd1 vssd1 vccd1 vccd1 _7027_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1540 _7356_/Q vssd1 vssd1 vccd1 vccd1 _7065_/A sky130_fd_sc_hd__buf_2
Xhold1551 _6943_/X vssd1 vssd1 vccd1 vccd1 _6944_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1562 hold1562/A vssd1 vssd1 vccd1 vccd1 _4775_/B sky130_fd_sc_hd__clkbuf_2
Xhold1595 _3757_/B vssd1 vssd1 vccd1 vccd1 _6437_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1584 _7040_/Y vssd1 vssd1 vccd1 vccd1 _7041_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1573 _4271_/Y vssd1 vssd1 vccd1 vccd1 _4272_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4856__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4608__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6383__B1 _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6686__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7105__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4544__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4448__B _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6663__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3779__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4464__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6610__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4847__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3961_ _5921_/A _5918_/A vssd1 vssd1 vccd1 vccd1 _3962_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6071__C1 _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5700_ _6056_/A _6075_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5700_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6680_ _6927_/A _6669_/B _6702_/B1 hold573/X vssd1 vssd1 vccd1 vccd1 _6680_/X sky130_fd_sc_hd__a22o_1
X_3892_ _6223_/A vssd1 vssd1 vccd1 vccd1 _3892_/Y sky130_fd_sc_hd__inv_2
X_5631_ _6927_/A _5620_/B _5653_/B1 _5631_/B2 vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6374__A0 _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5562_ _6548_/A _5562_/B vssd1 vssd1 vccd1 vccd1 _7751_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3727__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8350_ _8350_/CLK _8350_/D vssd1 vssd1 vccd1 vccd1 _8350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4513_ _5126_/A1 _4449_/A _5442_/C vssd1 vssd1 vccd1 vccd1 _7285_/D sky130_fd_sc_hd__mux2_1
X_8281_ _8475_/CLK _8281_/D vssd1 vssd1 vccd1 vccd1 _8281_/Q sky130_fd_sc_hd__dfxtp_1
X_7301_ _8501_/CLK _7301_/D _7111_/Y vssd1 vssd1 vccd1 vccd1 _7301_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__6677__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold125 _6503_/X vssd1 vssd1 vccd1 vccd1 _7985_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 _5658_/X vssd1 vssd1 vccd1 vccd1 _7838_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ _7514_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7682_/D sky130_fd_sc_hd__and3_1
Xhold114 _7601_/Q vssd1 vssd1 vccd1 vccd1 _5659_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4444_ _4440_/A _5442_/C _4443_/X _4442_/X vssd1 vssd1 vccd1 vccd1 _8361_/D sky130_fd_sc_hd__a31o_1
Xhold147 _6462_/X vssd1 vssd1 vccd1 vccd1 _7944_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _8445_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold158 _7863_/Q vssd1 vssd1 vccd1 vccd1 _6484_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold136 _7858_/Q vssd1 vssd1 vccd1 vccd1 _6479_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4783__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold169 _6499_/X vssd1 vssd1 vccd1 vccd1 _7981_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4375_ _4383_/A _4383_/B _4341_/C _4377_/B _4354_/C vssd1 vssd1 vccd1 vccd1 _4375_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7015__A _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7094_ _5389_/A _5374_/A _5409_/A vssd1 vssd1 vccd1 vccd1 _7094_/X sky130_fd_sc_hd__o21a_1
X_6114_ _6115_/A _6115_/B vssd1 vssd1 vccd1 vccd1 _6114_/Y sky130_fd_sc_hd__nand2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _4032_/A _6398_/A2 _6413_/B1 _6032_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _6045_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4535__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5652__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_A _6776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout451_A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7996_ _8385_/CLK hold48/X vssd1 vssd1 vccd1 vccd1 _7996_/Q sky130_fd_sc_hd__dfxtp_1
X_6947_ _6947_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6947_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6878_ _4775_/A _6878_/A2 _6845_/B _6877_/X vssd1 vssd1 vccd1 vccd1 _6878_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5829_ _5816_/Y _5827_/X _5828_/X _4775_/A vssd1 vssd1 vccd1 vccd1 _7870_/D sky130_fd_sc_hd__o211a_1
XANTENNA__6365__B1 _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8479_ _8479_/CLK _8479_/D vssd1 vssd1 vccd1 vccd1 _8479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4391__A2 _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5340__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold670 _5202_/X vssd1 vssd1 vccd1 vccd1 _7416_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold681 _8147_/Q vssd1 vssd1 vccd1 vccd1 hold681/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5371__C _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold692 _6675_/X vssd1 vssd1 vccd1 vccd1 _8202_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5643__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6840__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1370 _6948_/X vssd1 vssd1 vccd1 vccd1 _8439_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1381 _6630_/X vssd1 vssd1 vccd1 vccd1 _8179_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1392 _8372_/Q vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_115_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4829__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5099__B _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3709__A2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6939__A _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5331__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4459__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4160_ _5552_/B _4448_/A _7082_/A vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4091_ _3950_/X _3951_/Y _4045_/X _3935_/X _3922_/Y vssd1 vssd1 vccd1 vccd1 _4092_/D
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4893__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5634__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7850_ _8370_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_6801_ _6933_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6801_/X sky130_fd_sc_hd__and2_1
XANTENNA__5398__A1 _7065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4993_ _8357_/Q _7833_/Q _7499_/Q _7467_/Q _4997_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4993_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7781_ _8431_/CLK _7781_/D vssd1 vssd1 vccd1 vccd1 _7781_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3948__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3944_ _3944_/A vssd1 vssd1 vccd1 vccd1 _5763_/B sky130_fd_sc_hd__inv_2
XFILLER_0_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6732_ _6959_/A _6737_/A2 _6737_/B1 _6732_/B2 vssd1 vssd1 vccd1 vccd1 _6732_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6347__B1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6663_ _6969_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6663_/X sky130_fd_sc_hd__and2_1
X_3875_ _8090_/Q _3874_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3875_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8402_ _8402_/CLK _8402_/D vssd1 vssd1 vccd1 vccd1 _8402_/Q sky130_fd_sc_hd__dfxtp_1
X_5614_ _6965_/A _5616_/A2 _5616_/B1 hold831/X vssd1 vssd1 vccd1 vccd1 _5614_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6898__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5456__C _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6594_ _7074_/A _7069_/A _6597_/B _7067_/A vssd1 vssd1 vccd1 vccd1 _6595_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_61_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6849__A _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5545_ _5545_/A _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7734_/D sky130_fd_sc_hd__and3_1
X_8333_ _8478_/CLK _8333_/D vssd1 vssd1 vccd1 vccd1 _8333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8264_ _8458_/CLK _8264_/D vssd1 vssd1 vccd1 vccd1 _8264_/Q sky130_fd_sc_hd__dfxtp_1
X_5476_ _5476_/A _7088_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _7665_/D sky130_fd_sc_hd__and3_1
X_4427_ _4427_/A _4427_/B vssd1 vssd1 vccd1 vccd1 _4427_/X sky130_fd_sc_hd__or2_1
XANTENNA__5472__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5322__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8195_ _8195_/CLK _8195_/D vssd1 vssd1 vccd1 vccd1 _8195_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout413 _5476_/A vssd1 vssd1 vccd1 vccd1 _4867_/S1 sky130_fd_sc_hd__buf_4
Xfanout402 hold1746/X vssd1 vssd1 vccd1 vccd1 _7059_/A sky130_fd_sc_hd__buf_6
Xfanout457 _5667_/A vssd1 vssd1 vccd1 vccd1 _6552_/A sky130_fd_sc_hd__buf_2
Xfanout424 hold1747/X vssd1 vssd1 vccd1 vccd1 _5475_/A sky130_fd_sc_hd__buf_8
Xfanout446 _4775_/A vssd1 vssd1 vccd1 vccd1 _7029_/A sky130_fd_sc_hd__buf_4
X_4358_ _5580_/B _5062_/A1 _7030_/B vssd1 vssd1 vccd1 vccd1 _4358_/X sky130_fd_sc_hd__mux2_1
Xfanout435 _6545_/A vssd1 vssd1 vccd1 vccd1 _7022_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__5086__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout468 input63/X vssd1 vssd1 vccd1 vccd1 _7258_/A sky130_fd_sc_hd__buf_8
X_7077_ _7077_/A _7079_/B _7079_/C vssd1 vssd1 vccd1 vccd1 _8512_/D sky130_fd_sc_hd__and3_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _5570_/B _5042_/A1 _5540_/B vssd1 vssd1 vccd1 vccd1 _4397_/B sky130_fd_sc_hd__mux2_1
X_6028_ _5799_/X _5810_/B _6028_/S vssd1 vssd1 vccd1 vccd1 _6028_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6822__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3720__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7979_ _8365_/CLK _7979_/D vssd1 vssd1 vccd1 vccd1 _7979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6586__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6050__A2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5010__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5663__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4978__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7066__A1 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6494__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5616__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6941__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6577__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5838__A _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4052__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3660_ _7667_/Q vssd1 vssd1 vccd1 vccd1 _3660_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_70_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6669__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4986__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5330_ _6967_/A _5299_/B _5331_/B1 hold410/X vssd1 vssd1 vccd1 vccd1 _5330_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5573__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_53_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5261_ _6908_/C _6776_/A vssd1 vssd1 vccd1 vccd1 _5263_/B sky130_fd_sc_hd__or2_1
XANTENNA__5304__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4107__A2 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7000_ _7010_/A _7000_/B vssd1 vssd1 vccd1 vccd1 _7000_/X sky130_fd_sc_hd__and2_1
X_4212_ _4212_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__xor2_1
XANTENNA__4738__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5192_ _6847_/A _5189_/B _5189_/Y hold286/X vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3866__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4143_ _7596_/Q _8165_/Q _8455_/Q vssd1 vssd1 vccd1 vccd1 _4143_/X sky130_fd_sc_hd__and3b_1
XANTENNA__5607__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6804__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_68_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4074_ _4074_/A0 _4073_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6112_/A sky130_fd_sc_hd__mux2_2
X_7902_ _8507_/CLK _7902_/D vssd1 vssd1 vccd1 vccd1 _7902_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_111_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4910__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7833_ _8469_/CLK _7833_/D vssd1 vssd1 vccd1 vccd1 _7833_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6568__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6851__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5748__A _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7764_ _8382_/CLK _7764_/D vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5240__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6715_ _6925_/A _6705_/B _6738_/B1 hold581/X vssd1 vssd1 vccd1 vccd1 _6715_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5467__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4976_ _8484_/Q _8416_/Q _8448_/Q _8322_/Q _7063_/A _4976_/S1 vssd1 vssd1 vccd1 vccd1
+ _4976_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout247_A _6705_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3927_ _4014_/A _5549_/B vssd1 vssd1 vccd1 vccd1 _3927_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4371__B _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7695_ _8195_/CLK _7695_/D vssd1 vssd1 vccd1 vccd1 _7695_/Q sky130_fd_sc_hd__dfxtp_1
X_6646_ _7019_/A _6646_/A2 _6605_/B _6645_/X vssd1 vssd1 vccd1 vccd1 _6646_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_74_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout414_A hold1729/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3858_ _6244_/A _6242_/A vssd1 vssd1 vccd1 vccd1 _3859_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6577_ _6941_/A _6592_/A2 _6591_/B1 hold843/X vssd1 vssd1 vccd1 vccd1 _6577_/X sky130_fd_sc_hd__a22o_1
X_3789_ _4067_/A_N _7958_/Q vssd1 vssd1 vccd1 vccd1 _3789_/X sky130_fd_sc_hd__and2b_1
X_5528_ _8247_/Q _5528_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7717_/D sky130_fd_sc_hd__and3_1
X_8316_ _8478_/CLK _8316_/D vssd1 vssd1 vccd1 vccd1 _8316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8247_ _8247_/CLK _8247_/D vssd1 vssd1 vccd1 vccd1 _8247_/Q sky130_fd_sc_hd__dfxtp_1
X_5459_ _5459_/A _5503_/B _5462_/C vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__and3_1
X_8178_ _8338_/CLK _8178_/D vssd1 vssd1 vccd1 vccd1 _8178_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout232 _4370_/X vssd1 vssd1 vccd1 vccd1 _7073_/B sky130_fd_sc_hd__buf_6
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout210 _5734_/X vssd1 vssd1 vccd1 vccd1 _6063_/A sky130_fd_sc_hd__buf_4
Xfanout221 _5470_/C vssd1 vssd1 vccd1 vccd1 _7030_/C sky130_fd_sc_hd__buf_4
Xfanout254 _5620_/Y vssd1 vssd1 vccd1 vccd1 _5653_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout243 _4082_/B1 vssd1 vssd1 vccd1 vccd1 _4071_/B1 sky130_fd_sc_hd__buf_8
Xfanout265 _5188_/Y vssd1 vssd1 vccd1 vccd1 _5220_/B1 sky130_fd_sc_hd__buf_6
Xfanout276 _6908_/X vssd1 vssd1 vccd1 vccd1 _6943_/B sky130_fd_sc_hd__clkbuf_16
Xfanout298 _6557_/Y vssd1 vssd1 vccd1 vccd1 _6592_/A2 sky130_fd_sc_hd__buf_6
XANTENNA__3731__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout287 _6741_/B vssd1 vssd1 vccd1 vccd1 _6773_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5658__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4034__B2 _8012_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3793__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6489__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4968__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6731__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7113__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5696__S1 _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4472__A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _4829_/X _4828_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4830_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5568__A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7213__91 _8419_/CLK vssd1 vssd1 vccd1 vccd1 _8126_/CLK sky130_fd_sc_hd__inv_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4761_ _6534_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _8118_/D sky130_fd_sc_hd__and2_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6500_ _7006_/A _6500_/B vssd1 vssd1 vccd1 vccd1 _6500_/X sky130_fd_sc_hd__and2_1
X_7480_ _8332_/CLK _7480_/D vssd1 vssd1 vccd1 vccd1 _7480_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3712_ _6298_/A _6295_/A vssd1 vssd1 vccd1 vccd1 _3714_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4692_ _8480_/Q _8412_/Q _8444_/Q _8318_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4692_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6431_ _6552_/A _6431_/B vssd1 vssd1 vccd1 vccd1 _7913_/D sky130_fd_sc_hd__and2_1
XFILLER_0_43_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4959__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6722__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6362_ _6412_/S _6362_/B _6362_/C vssd1 vssd1 vccd1 vccd1 _6362_/X sky130_fd_sc_hd__and3_1
XFILLER_0_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5313_ _6933_/A _5332_/A2 _5332_/B1 _5313_/B2 vssd1 vssd1 vccd1 vccd1 _5313_/X sky130_fd_sc_hd__a22o_1
X_8101_ _8101_/CLK _8101_/D vssd1 vssd1 vccd1 vccd1 _8101_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_577 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5289__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6293_ _6391_/A _6283_/X _6292_/X vssd1 vssd1 vccd1 vccd1 _6293_/X sky130_fd_sc_hd__o21ba_1
X_5244_ _6941_/A _5258_/A2 _5258_/B1 hold419/X vssd1 vssd1 vccd1 vccd1 _5244_/X sky130_fd_sc_hd__a22o_1
X_8032_ _8032_/CLK _8032_/D vssd1 vssd1 vccd1 vccd1 _8032_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3839__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5175_ hold67/X _5468_/C vssd1 vssd1 vccd1 vccd1 _5175_/X sky130_fd_sc_hd__or2_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7023__A _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4126_ _4124_/X _4125_/Y _3788_/A vssd1 vssd1 vccd1 vccd1 _4126_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4057_ _8079_/Q _4056_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__mux2_2
XANTENNA_fanout364_A _3657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5478__A _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7816_ _8154_/CLK _7816_/D vssd1 vssd1 vccd1 vccd1 _7816_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5213__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7747_ _8510_/CLK _7747_/D vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4959_ _8159_/Q _7558_/Q _7430_/Q _7590_/Q _4990_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4959_/X sky130_fd_sc_hd__mux4_1
X_7678_ _8428_/CLK _7678_/D vssd1 vssd1 vccd1 vccd1 _7678_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6629_ _6935_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6629_/X sky130_fd_sc_hd__and2_1
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6713__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4991__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5755__A1 _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3766__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7108__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6947__A _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4467__A _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6980_ _6597_/B _5385_/Y _6978_/X _6979_/X vssd1 vssd1 vccd1 vccd1 _6980_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5931_ _5927_/X _5930_/Y _6251_/A vssd1 vssd1 vccd1 vccd1 _5931_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6786__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5862_ _5858_/X _5861_/X _6302_/A vssd1 vssd1 vccd1 vccd1 _5862_/X sky130_fd_sc_hd__mux2_1
X_4813_ _4811_/X _4812_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__mux2_1
X_5793_ _6028_/S _6083_/A vssd1 vssd1 vccd1 vccd1 _5793_/Y sky130_fd_sc_hd__nor2_2
X_7601_ _8361_/CLK _7601_/D vssd1 vssd1 vccd1 vccd1 _7601_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5746__A1 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4744_ _7006_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _8101_/D sky130_fd_sc_hd__and2_1
X_7532_ _8136_/CLK _7532_/D vssd1 vssd1 vccd1 vccd1 _7532_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4119__A_N _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4675_ _8155_/Q _7554_/Q _7426_/Q _7586_/Q _4720_/S0 _4741_/S1 vssd1 vssd1 vccd1
+ vccd1 _4675_/X sky130_fd_sc_hd__mux4_1
XANTENNA__7018__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7463_ _8353_/CLK _7463_/D vssd1 vssd1 vccd1 vccd1 _7463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6414_ _6405_/A _6414_/A2 _6414_/B1 _3846_/B _6413_/X vssd1 vssd1 vccd1 vccd1 _6416_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5464__C _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7394_ _8373_/CLK _7394_/D vssd1 vssd1 vccd1 vccd1 _7394_/Q sky130_fd_sc_hd__dfxtp_1
X_6345_ _3749_/A _6414_/B1 _6398_/B1 _6331_/A _6292_/A vssd1 vssd1 vccd1 vccd1 _6345_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__6857__A _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6276_ _3883_/B _6292_/A _6347_/B1 vssd1 vssd1 vccd1 vccd1 _6276_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5227_ _7010_/A _5227_/B vssd1 vssd1 vccd1 vccd1 _5227_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5480__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8015_ _8034_/CLK _8015_/D vssd1 vssd1 vccd1 vccd1 _8015_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1711 _7639_/Q vssd1 vssd1 vccd1 vccd1 _4216_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1700 _7688_/Q vssd1 vssd1 vccd1 vccd1 _3863_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1722 _7668_/Q vssd1 vssd1 vccd1 vccd1 _3926_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4580__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1733 _6030_/X vssd1 vssd1 vccd1 vccd1 _6031_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1744 _6140_/A vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _5158_/A1 _5069_/S _5002_/X _5157_/X vssd1 vssd1 vccd1 vccd1 _7391_/D sky130_fd_sc_hd__o211a_1
Xhold1766 _6071_/Y vssd1 vssd1 vccd1 vccd1 _7880_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _4109_/A _4109_/B vssd1 vssd1 vccd1 vccd1 _4109_/X sky130_fd_sc_hd__or2_1
Xhold1777 _6092_/X vssd1 vssd1 vccd1 vccd1 _7881_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5089_ _5089_/A _5538_/C vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__or2_1
Xhold1755 _7718_/Q vssd1 vssd1 vccd1 vccd1 _3780_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1799 _7877_/Q vssd1 vssd1 vccd1 vccd1 hold1799/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5700__S _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1788 _7722_/Q vssd1 vssd1 vccd1 vccd1 _3852_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5001__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3903__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4226__S _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3987__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6007__A _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4750__A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3739__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6940__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4460_ _6552_/A _7927_/Q vssd1 vssd1 vccd1 vccd1 _8059_/D sky130_fd_sc_hd__and2_1
XFILLER_0_53_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold307 _5463_/X vssd1 vssd1 vccd1 vccd1 _7652_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _7870_/Q vssd1 vssd1 vccd1 vccd1 _4746_/B sky130_fd_sc_hd__buf_1
Xhold329 _5469_/X vssd1 vssd1 vccd1 vccd1 _7658_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4391_ _4387_/A _5465_/C _4390_/X _4389_/X vssd1 vssd1 vccd1 vccd1 _8380_/D sky130_fd_sc_hd__a31o_1
X_6130_ _6130_/A _6130_/B vssd1 vssd1 vccd1 vccd1 _6130_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ _4066_/A _6398_/A2 _6413_/B1 _6053_/A vssd1 vssd1 vccd1 vccd1 _6063_/B sky130_fd_sc_hd__a22o_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4562__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1029 _7541_/Q vssd1 vssd1 vccd1 vccd1 _5310_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_5012_ hold212/X _5085_/B _5140_/B1 _5011_/X vssd1 vssd1 vccd1 vccd1 _5012_/X sky130_fd_sc_hd__o211a_1
Xhold1007 _8475_/Q vssd1 vssd1 vccd1 vccd1 _7017_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1018 _5219_/X vssd1 vssd1 vccd1 vccd1 _7433_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6843__C _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5967__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6963_ _6963_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6963_/X sky130_fd_sc_hd__and2_1
X_5914_ _5914_/A _5914_/B vssd1 vssd1 vccd1 vccd1 _5914_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6894_ _7019_/A _6894_/A2 _6906_/A3 _6893_/X vssd1 vssd1 vccd1 vccd1 _6894_/X sky130_fd_sc_hd__a31o_1
X_5845_ _5846_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5845_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5756__A _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5475__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5195__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5776_ _5846_/A _5765_/A _5870_/A _5820_/A _5804_/A _5789_/S vssd1 vssd1 vccd1 vccd1
+ _5776_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6392__A1 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8495_ _8501_/CLK _8495_/D vssd1 vssd1 vccd1 vccd1 _8495_/Q sky130_fd_sc_hd__dfxtp_1
X_7515_ _7515_/CLK _7515_/D vssd1 vssd1 vccd1 vccd1 _7515_/Q sky130_fd_sc_hd__dfxtp_1
X_4727_ _8485_/Q _8417_/Q _8449_/Q _8323_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4727_/X sky130_fd_sc_hd__mux4_1
X_7446_ _8332_/CLK _7446_/D vssd1 vssd1 vccd1 vccd1 _7446_/Q sky130_fd_sc_hd__dfxtp_1
X_4658_ _4657_/X _4656_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4658_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold830 _5638_/X vssd1 vssd1 vccd1 vccd1 _7818_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6695__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4589_ _4588_/X _4585_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7509_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_101_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3902__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold841 _8229_/Q vssd1 vssd1 vccd1 vccd1 hold841/X sky130_fd_sc_hd__dlygate4sd3_1
X_7377_ _8515_/CLK _7377_/D vssd1 vssd1 vccd1 vccd1 _7377_/Q sky130_fd_sc_hd__dfxtp_1
Xhold852 _6572_/X vssd1 vssd1 vccd1 vccd1 _8144_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 _8273_/Q vssd1 vssd1 vccd1 vccd1 hold863/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold874 _5236_/X vssd1 vssd1 vccd1 vccd1 _7444_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 _7787_/Q vssd1 vssd1 vccd1 vccd1 hold885/X sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ _6412_/S _6325_/X _6327_/X vssd1 vssd1 vccd1 vccd1 _6328_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold896 _7027_/X vssd1 vssd1 vccd1 vccd1 _8485_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6259_ _6259_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6262_/B sky130_fd_sc_hd__xnor2_1
Xhold1530 _6844_/X vssd1 vssd1 vccd1 vccd1 _8388_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1541 _7065_/Y vssd1 vssd1 vccd1 vccd1 _7066_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 _6944_/X vssd1 vssd1 vccd1 vccd1 _8437_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1563 _8425_/Q vssd1 vssd1 vccd1 vccd1 _6919_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1585 hold1811/X vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__clkbuf_2
Xhold1574 _4272_/Y vssd1 vssd1 vccd1 vccd1 _4274_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1596 _8491_/Q vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5666__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6922__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5385__B _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6686__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6497__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5110__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5646__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4544__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4745__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7121__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3960_ _5921_/A _5918_/A vssd1 vssd1 vccd1 vccd1 _3962_/A sky130_fd_sc_hd__or2_1
XFILLER_0_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5576__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3891_ _3891_/A0 _3890_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6223_/A sky130_fd_sc_hd__mux2_2
XANTENNA__4480__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5630_ _6925_/A _5620_/B _5653_/B1 hold491/X vssd1 vssd1 vccd1 vccd1 _5630_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6374__A1 _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5561_ _6534_/A _5561_/B vssd1 vssd1 vccd1 vccd1 _7750_/D sky130_fd_sc_hd__and2_1
XFILLER_0_41_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5492_ _7513_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7681_/D sky130_fd_sc_hd__and3_1
XFILLER_0_81_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4512_ _5128_/A1 _4171_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _7286_/D sky130_fd_sc_hd__mux2_1
XANTENNA__3801__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7300_ _8501_/CLK _7300_/D _7110_/Y vssd1 vssd1 vccd1 vccd1 _7300_/Q sky130_fd_sc_hd__dfrtp_4
X_8280_ _8476_/CLK _8280_/D vssd1 vssd1 vccd1 vccd1 _8280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6677__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold126 _7610_/Q vssd1 vssd1 vccd1 vccd1 _5668_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _5659_/X vssd1 vssd1 vccd1 vccd1 _7839_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 _7615_/Q vssd1 vssd1 vccd1 vccd1 _5673_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _7607_/Q vssd1 vssd1 vccd1 vccd1 _5665_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _4449_/A _4449_/B _4171_/B _4178_/B vssd1 vssd1 vccd1 vccd1 _4443_/X sky130_fd_sc_hd__a31o_1
Xhold159 _6484_/X vssd1 vssd1 vccd1 vccd1 _7966_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold137 _6479_/X vssd1 vssd1 vccd1 vccd1 _7961_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4783__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4374_ _5062_/A1 _5182_/A2 _4372_/Y _4373_/X vssd1 vssd1 vccd1 vccd1 _8387_/D sky130_fd_sc_hd__a22o_1
X_7093_ _5389_/A _5374_/A _5409_/A vssd1 vssd1 vccd1 vccd1 _7093_/X sky130_fd_sc_hd__o21a_1
X_6113_ _6115_/A _6115_/B vssd1 vssd1 vccd1 vccd1 _6116_/A sky130_fd_sc_hd__and2_1
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ _5694_/Y _6043_/X _6042_/Y vssd1 vssd1 vccd1 vccd1 _6044_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5637__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4535__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7031__A _7031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout277_A _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7995_ _8020_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 _7995_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6062__B1 _6060_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout444_A _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6946_ _7028_/A _6946_/A2 _6970_/A3 _6945_/X vssd1 vssd1 vccd1 vccd1 _6946_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_119_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6877_ _6877_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6877_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5828_ _5820_/A _5963_/S _6063_/A vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5168__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5759_ _5759_/A vssd1 vssd1 vccd1 vccd1 _5759_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6904__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3718__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7174__52 _8472_/CLK vssd1 vssd1 vccd1 vccd1 _8054_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_44_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8478_ _8478_/CLK _8478_/D vssd1 vssd1 vccd1 vccd1 _8478_/Q sky130_fd_sc_hd__dfxtp_1
X_7429_ _8413_/CLK _7429_/D vssd1 vssd1 vccd1 vccd1 _7429_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold660 _5628_/X vssd1 vssd1 vccd1 vccd1 _7808_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold671 _7833_/Q vssd1 vssd1 vccd1 vccd1 hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold682 _6575_/X vssd1 vssd1 vccd1 vccd1 _8147_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold693 _7554_/Q vssd1 vssd1 vccd1 vccd1 hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5628__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1360 _8343_/Q vssd1 vssd1 vccd1 vccd1 _6812_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1393 _8365_/Q vssd1 vssd1 vccd1 vccd1 _5018_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1371 _8405_/Q vssd1 vssd1 vccd1 vccd1 _6878_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1382 _8374_/Q vssd1 vssd1 vccd1 vccd1 _5036_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3824__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4504__S _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5843__B _5971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6939__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5828__B1_N _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7116__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5331__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6955__A _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4090_ _4090_/A _4090_/B _4115_/A _4090_/D vssd1 vssd1 vccd1 vccd1 _4092_/C sky130_fd_sc_hd__or4_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4475__A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7233__111 _8328_/CLK vssd1 vssd1 vccd1 vccd1 _8243_/CLK sky130_fd_sc_hd__inv_2
X_6800_ _7023_/A _6800_/A2 _6838_/A3 _6799_/X vssd1 vssd1 vccd1 vccd1 _6800_/X sky130_fd_sc_hd__a31o_1
X_7780_ _8332_/CLK _7780_/D vssd1 vssd1 vccd1 vccd1 _7780_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4992_ _4991_/X _4988_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8260_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_105_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _4014_/A _8518_/Q vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6731_ _6891_/A _6737_/A2 _6737_/B1 hold797/X vssd1 vssd1 vccd1 vccd1 _6731_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3874_ _7994_/Q _4068_/A2 _4068_/B1 _8026_/Q _3873_/X vssd1 vssd1 vccd1 vccd1 _3874_/X
+ sky130_fd_sc_hd__a221o_1
X_6662_ _7027_/A _6662_/A2 _6605_/B _6661_/X vssd1 vssd1 vccd1 vccd1 _6662_/X sky130_fd_sc_hd__a31o_1
X_8401_ _8469_/CLK _8401_/D vssd1 vssd1 vccd1 vccd1 _8401_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5613_ _6963_/A _5616_/A2 _5616_/B1 hold761/X vssd1 vssd1 vccd1 vccd1 _5613_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8332_ _8332_/CLK _8332_/D vssd1 vssd1 vccd1 vccd1 _8332_/Q sky130_fd_sc_hd__dfxtp_1
X_6593_ _6597_/B _7067_/A _7069_/A vssd1 vssd1 vccd1 vccd1 _6593_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_54_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6849__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5544_ _5544_/A _7088_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5544_/X sky130_fd_sc_hd__and3_1
XFILLER_0_112_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8263_ _8458_/CLK _8263_/D vssd1 vssd1 vccd1 vccd1 _8263_/Q sky130_fd_sc_hd__dfxtp_1
X_5475_ _5475_/A _7088_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _7664_/D sky130_fd_sc_hd__and3_1
X_4426_ _5024_/A1 _4425_/B _4424_/X _4425_/Y vssd1 vssd1 vccd1 vccd1 _8368_/D sky130_fd_sc_hd__a22o_1
XANTENNA__5472__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5322__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8194_ _8354_/CLK _8194_/D vssd1 vssd1 vccd1 vccd1 _8194_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7026__A _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout403 _5477_/A vssd1 vssd1 vccd1 vccd1 _4998_/S sky130_fd_sc_hd__buf_8
Xfanout414 hold1729/X vssd1 vssd1 vccd1 vccd1 _5476_/A sky130_fd_sc_hd__buf_6
XANTENNA_fanout394_A _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout447 _7007_/A vssd1 vssd1 vccd1 vccd1 _7008_/A sky130_fd_sc_hd__buf_4
X_4357_ _4357_/A _4357_/B vssd1 vssd1 vccd1 vccd1 _4357_/Y sky130_fd_sc_hd__xnor2_1
Xfanout425 _7283_/Q vssd1 vssd1 vccd1 vccd1 _4067_/A_N sky130_fd_sc_hd__buf_4
XANTENNA__6865__A _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _7027_/A vssd1 vssd1 vccd1 vccd1 _6545_/A sky130_fd_sc_hd__clkbuf_4
Xfanout458 _4775_/A vssd1 vssd1 vccd1 vccd1 _5667_/A sky130_fd_sc_hd__clkbuf_4
Xfanout469 input63/X vssd1 vssd1 vccd1 vccd1 _7264_/A sky130_fd_sc_hd__clkbuf_8
X_7076_ _7076_/A _7079_/B _7079_/C vssd1 vssd1 vccd1 vccd1 _8511_/D sky130_fd_sc_hd__and3_1
XANTENNA__5086__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4288_/A _4288_/B vssd1 vssd1 vccd1 vccd1 _4288_/X sky130_fd_sc_hd__xor2_1
X_6027_ _6250_/S _5792_/Y _6026_/X vssd1 vssd1 vccd1 vccd1 _6027_/Y sky130_fd_sc_hd__o21ai_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6586__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7978_ _8387_/CLK _7978_/D vssd1 vssd1 vccd1 vccd1 _7978_/Q sky130_fd_sc_hd__dfxtp_1
X_6929_ _6929_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6929_/X sky130_fd_sc_hd__and2_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1676_A _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4692__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5944__A _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5313__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold490 _5242_/X vssd1 vssd1 vccd1 vccd1 _7450_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1190 _6652_/X vssd1 vssd1 vccd1 vccd1 _8190_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6121__S0 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6577__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4052__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6015__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6329__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_467 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6329__B2 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6669__B _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4986__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5260_ _6908_/C _6776_/A vssd1 vssd1 vccd1 vccd1 _5260_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4211_ _4201_/Y _4205_/B _4203_/B vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__o21a_1
XANTENNA__4738__S1 _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5191_ _3939_/C _5189_/B _5189_/Y hold344/X vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3866__A2 _6441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4142_ _4117_/Y _4141_/Y _4152_/A vssd1 vssd1 vccd1 vccd1 _4144_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__3821__B _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4073_ _4073_/A1 _4073_/A2 _6939_/A _4073_/B2 _4072_/X vssd1 vssd1 vccd1 vccd1 _4073_/X
+ sky130_fd_sc_hd__a221o_2
X_7901_ _8507_/CLK _7901_/D vssd1 vssd1 vccd1 vccd1 _7901_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4910__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6568__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7832_ _8484_/CLK _7832_/D vssd1 vssd1 vccd1 vccd1 _7832_/Q sky130_fd_sc_hd__dfxtp_1
X_4975_ _8194_/Q _8226_/Q _8290_/Q _7798_/Q _7063_/A _4976_/S1 vssd1 vssd1 vccd1 vccd1
+ _4975_/X sky130_fd_sc_hd__mux4_1
X_7763_ _8071_/CLK _7763_/D vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3926_ _3926_/A1 _4084_/A2 _6777_/A _4084_/B2 _3925_/X vssd1 vssd1 vccd1 vccd1 _6421_/B
+ sky130_fd_sc_hd__a221oi_4
X_6714_ _6923_/A _6737_/A2 _6737_/B1 hold591/X vssd1 vssd1 vccd1 vccd1 _6714_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4674__S0 _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7694_ _8355_/CLK _7694_/D vssd1 vssd1 vccd1 vccd1 _7694_/Q sky130_fd_sc_hd__dfxtp_1
X_6645_ _6951_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6645_/X sky130_fd_sc_hd__and2_1
XFILLER_0_61_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3857_ _6244_/A _6242_/A vssd1 vssd1 vccd1 vccd1 _3859_/A sky130_fd_sc_hd__or2_1
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7144__22 _8413_/CLK vssd1 vssd1 vccd1 vccd1 _7521_/CLK sky130_fd_sc_hd__inv_2
X_3788_ _3788_/A vssd1 vssd1 vccd1 vccd1 _3800_/C sky130_fd_sc_hd__inv_2
X_6576_ _6939_/A _6559_/B _6591_/B1 _6576_/B2 vssd1 vssd1 vccd1 vccd1 _6576_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout407_A _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8315_ _8477_/CLK _8315_/D vssd1 vssd1 vccd1 vccd1 _8315_/Q sky130_fd_sc_hd__dfxtp_1
X_5527_ _8246_/Q _5542_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7716_/D sky130_fd_sc_hd__and3_1
XFILLER_0_112_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8246_ _8246_/CLK _8246_/D vssd1 vssd1 vccd1 vccd1 _8246_/Q sky130_fd_sc_hd__dfxtp_1
X_5458_ _5458_/A _5465_/B _5463_/C vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5389_ _5389_/A _6553_/A _5391_/A vssd1 vssd1 vccd1 vccd1 _5389_/X sky130_fd_sc_hd__or3b_1
Xfanout200 _3919_/X vssd1 vssd1 vccd1 vccd1 _6393_/A sky130_fd_sc_hd__clkbuf_4
Xfanout211 _5734_/X vssd1 vssd1 vccd1 vccd1 _6011_/A2 sky130_fd_sc_hd__buf_4
Xfanout222 _7073_/B vssd1 vssd1 vccd1 vccd1 _5470_/C sky130_fd_sc_hd__clkbuf_4
X_8177_ _8467_/CLK _8177_/D vssd1 vssd1 vccd1 vccd1 _8177_/Q sky130_fd_sc_hd__dfxtp_1
X_4409_ _4419_/A _4415_/B _4413_/B _4262_/C vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__a31o_1
Xfanout244 _3676_/Y vssd1 vssd1 vccd1 vccd1 _4082_/B1 sky130_fd_sc_hd__clkbuf_16
Xfanout255 _5584_/Y vssd1 vssd1 vccd1 vccd1 _5616_/B1 sky130_fd_sc_hd__buf_8
Xfanout233 _5182_/A2 vssd1 vssd1 vccd1 vccd1 _4416_/B sky130_fd_sc_hd__buf_4
Xfanout288 _6739_/Y vssd1 vssd1 vccd1 vccd1 _6741_/B sky130_fd_sc_hd__buf_8
Xfanout266 _5188_/Y vssd1 vssd1 vccd1 vccd1 _5221_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout299 _6398_/A2 vssd1 vssd1 vccd1 vccd1 _6414_/B1 sky130_fd_sc_hd__clkbuf_8
X_7059_ _7059_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7059_/Y sky130_fd_sc_hd__nand2_1
Xfanout277 _6963_/B vssd1 vssd1 vccd1 vccd1 _6969_/B sky130_fd_sc_hd__buf_6
XFILLER_0_5_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4319__S _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5004__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4034__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3793__B2 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5674__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4968__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6731__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6798__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4753__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4656__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _7026_/A _4760_/B vssd1 vssd1 vccd1 vccd1 _8117_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6970__A1 _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5584__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3711_ _6295_/A vssd1 vssd1 vccd1 vccd1 _3711_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3784__A1 _3783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4691_ _8190_/Q _8222_/Q _8286_/Q _7794_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4691_/X sky130_fd_sc_hd__mux4_1
X_6430_ _7007_/A _6430_/B vssd1 vssd1 vccd1 vccd1 _7912_/D sky130_fd_sc_hd__and2_1
XANTENNA__6183__C1 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6722__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6361_ _6412_/S _6361_/B vssd1 vssd1 vccd1 vccd1 _6361_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4959__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8100_ _8513_/CLK _8100_/D vssd1 vssd1 vccd1 vccd1 _8100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5312_ _6931_/A _5299_/B _5331_/B1 hold398/X vssd1 vssd1 vccd1 vccd1 _5312_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5289__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6292_ _6292_/A _6292_/B _6292_/C _6292_/D vssd1 vssd1 vccd1 vccd1 _6292_/X sky130_fd_sc_hd__or4_1
XFILLER_0_3_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8031_ _8465_/CLK _8031_/D vssd1 vssd1 vccd1 vccd1 _8031_/Q sky130_fd_sc_hd__dfxtp_2
X_5243_ _6939_/A _5258_/A2 _5258_/B1 hold607/X vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3839__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5174_ _5174_/A1 _5069_/S _5182_/B1 _5173_/X vssd1 vssd1 vccd1 vccd1 _7399_/D sky130_fd_sc_hd__o211a_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_4125_ _3759_/A _3759_/B _6140_/A _3800_/B vssd1 vssd1 vccd1 vccd1 _4125_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_127_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4056_ _7983_/Q _4079_/A2 _4079_/B1 _8015_/Q _4055_/X vssd1 vssd1 vccd1 vccd1 _4056_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4895__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5478__B _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7815_ _8339_/CLK _7815_/D vssd1 vssd1 vccd1 vccd1 _7815_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout357_A _3837_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4382__B _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5213__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4647__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7746_ _8365_/CLK _7746_/D vssd1 vssd1 vccd1 vccd1 _7746_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4958_ _8352_/Q _7828_/Q _7494_/Q _7462_/Q _5089_/A _4969_/S1 vssd1 vssd1 vccd1 vccd1
+ _4958_/X sky130_fd_sc_hd__mux4_1
X_7677_ _8339_/CLK _7677_/D vssd1 vssd1 vccd1 vccd1 _7677_/Q sky130_fd_sc_hd__dfxtp_1
X_3909_ _5846_/A _6302_/A vssd1 vssd1 vccd1 vccd1 _3910_/B sky130_fd_sc_hd__or2_1
XFILLER_0_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4889_ _8149_/Q _7548_/Q _7420_/Q _7580_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4889_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6713__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6628_ _7010_/A _6628_/A2 _6605_/B _6627_/X vssd1 vssd1 vccd1 vccd1 _6628_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4602__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6559_ _6741_/A _6559_/B vssd1 vssd1 vccd1 vccd1 _6559_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8229_ _8487_/CLK _8229_/D vssd1 vssd1 vccd1 vccd1 _8229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5204__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6952__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_67_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4512__S _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6165__C1 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_110_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6947__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4748__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5140__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6963__A _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4877__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5930_ _6128_/A _5930_/B vssd1 vssd1 vccd1 vccd1 _5930_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5579__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4483__A _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7600_ _8364_/CLK _7600_/D vssd1 vssd1 vccd1 vccd1 _7600_/Q sky130_fd_sc_hd__dfxtp_1
X_5861_ _5859_/X _5860_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4629__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4812_ _8138_/Q _7537_/Q _7409_/Q _7569_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4812_/X sky130_fd_sc_hd__mux4_1
X_5792_ _5879_/S _5792_/B vssd1 vssd1 vccd1 vccd1 _5792_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5746__A2 _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4743_ _4742_/X _4739_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7531_/D sky130_fd_sc_hd__mux2_1
X_7531_ _7531_/CLK _7531_/D vssd1 vssd1 vccd1 vccd1 _7531_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7462_ _8353_/CLK _7462_/D vssd1 vssd1 vccd1 vccd1 _7462_/Q sky130_fd_sc_hd__dfxtp_1
X_6413_ _6126_/A _5881_/C _6413_/B1 _4118_/A _6292_/A vssd1 vssd1 vccd1 vccd1 _6413_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4674_ _8348_/Q _7824_/Q _7490_/Q _7458_/Q _4720_/S0 _4741_/S1 vssd1 vssd1 vccd1
+ vccd1 _4674_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4801__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7393_ _8071_/CLK _7393_/D vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6344_ _6412_/S _6047_/Y _6128_/X vssd1 vssd1 vccd1 vccd1 _6344_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6857__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6275_ _5957_/Y _6130_/A _6266_/A _6414_/A2 _6272_/X vssd1 vssd1 vccd1 vccd1 _6275_/X
+ sky130_fd_sc_hd__a221o_1
X_8014_ _8462_/CLK _8014_/D vssd1 vssd1 vccd1 vccd1 _8014_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5480__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5226_ _7267_/A _5226_/B vssd1 vssd1 vccd1 vccd1 _5226_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__7034__A _7075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1701 _7669_/Q vssd1 vssd1 vccd1 vccd1 _3941_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold1712 _4217_/B vssd1 vssd1 vccd1 vccd1 _4224_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1734 _6031_/Y vssd1 vssd1 vccd1 vccd1 _7878_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1723 _8494_/Q vssd1 vssd1 vccd1 vccd1 _3710_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5157_ _5458_/A _5463_/C vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__or2_1
XANTENNA__6873__A _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5088_ input5/X _4425_/B _5146_/B1 _5087_/X vssd1 vssd1 vccd1 vccd1 _7356_/D sky130_fd_sc_hd__o211a_1
Xhold1778 _7717_/Q vssd1 vssd1 vccd1 vccd1 _3768_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4108_ _4045_/A _4107_/X _4106_/Y vssd1 vssd1 vccd1 vccd1 _4109_/B sky130_fd_sc_hd__o21a_1
Xhold1767 _7714_/Q vssd1 vssd1 vccd1 vccd1 _4049_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1745 _6153_/X vssd1 vssd1 vccd1 vccd1 _7884_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1756 _7720_/Q vssd1 vssd1 vccd1 vccd1 _3868_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1789 _7701_/Q vssd1 vssd1 vccd1 vccd1 _3947_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4039_ _4039_/A1 _4084_/A2 _4035_/X _4084_/B2 _4038_/X vssd1 vssd1 vccd1 vccd1 _4039_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__4868__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1491_A _7310_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6934__A1 _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5198__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6395__C1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7729_ _8463_/CLK _7729_/D vssd1 vssd1 vccd1 vccd1 _7729_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_113_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8346_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6147__C1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6113__A _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6698__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5122__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6783__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3987__B2 _8008_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3647__A _7365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7119__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_104_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8442_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6023__A _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6689__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold308 _7340_/Q vssd1 vssd1 vccd1 vccd1 _5437_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold319 _8103_/D vssd1 vssd1 vccd1 vccd1 _8069_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5361__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4390_ _4390_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4478__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6060_ _6128_/A _6361_/B _6362_/C _6362_/B vssd1 vssd1 vccd1 vccd1 _6060_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _7318_/Q _5449_/C vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__or2_1
Xhold1008 _7017_/X vssd1 vssd1 vccd1 vccd1 _8475_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1019 _8227_/Q vssd1 vssd1 vccd1 vccd1 _6700_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6962_ _7024_/A _6962_/A2 _6970_/A3 _6961_/X vssd1 vssd1 vccd1 vccd1 _6962_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_16_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5913_ _6105_/A2 _5895_/A _5903_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _5914_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_88_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6893_ _6959_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6893_/X sky130_fd_sc_hd__and2_1
XANTENNA__6916__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5844_ _5846_/A _5846_/B vssd1 vssd1 vccd1 vccd1 _5847_/A sky130_fd_sc_hd__and2_1
XFILLER_0_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5756__B _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5775_ _5734_/A _5769_/Y _6163_/B _5740_/Y _5771_/Y vssd1 vssd1 vccd1 vccd1 _5775_/X
+ sky130_fd_sc_hd__o221a_1
X_7514_ _7514_/CLK _7514_/D vssd1 vssd1 vccd1 vccd1 _7514_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7029__A _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6392__A2 _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout222_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8494_ _8494_/CLK _8494_/D vssd1 vssd1 vccd1 vccd1 _8494_/Q sky130_fd_sc_hd__dfxtp_1
X_4726_ _8195_/Q _8227_/Q _8291_/Q _7799_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4726_/X sky130_fd_sc_hd__mux4_1
X_7445_ _8175_/CLK _7445_/D vssd1 vssd1 vccd1 vccd1 _7445_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4657_ _8475_/Q _8407_/Q _8439_/Q _8313_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4657_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7376_ _8360_/CLK _7376_/D vssd1 vssd1 vccd1 vccd1 _7376_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5352__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold820 _5637_/X vssd1 vssd1 vccd1 vccd1 _7817_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4588_ _4587_/X _4586_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4588_/X sky130_fd_sc_hd__mux2_1
Xhold842 _6702_/X vssd1 vssd1 vccd1 vccd1 _8229_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold831 _7798_/Q vssd1 vssd1 vccd1 vccd1 hold831/X sky130_fd_sc_hd__dlygate4sd3_1
X_6327_ _3750_/B _6414_/A2 _6019_/X _6130_/A _6326_/X vssd1 vssd1 vccd1 vccd1 _6327_/X
+ sky130_fd_sc_hd__a221o_1
Xhold864 _6718_/X vssd1 vssd1 vccd1 vccd1 _8273_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold853 _8312_/Q vssd1 vssd1 vccd1 vccd1 hold853/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold886 _5603_/X vssd1 vssd1 vccd1 vccd1 _7787_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3902__B2 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold875 _7578_/Q vssd1 vssd1 vccd1 vccd1 hold875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold897 _7559_/Q vssd1 vssd1 vccd1 vccd1 hold897/X sky130_fd_sc_hd__dlygate4sd3_1
X_6258_ _6253_/Y _6255_/X _6256_/Y _6257_/Y vssd1 vssd1 vccd1 vccd1 _7890_/D sky130_fd_sc_hd__o31a_1
XANTENNA__5104__B1 _5002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5209_ _6947_/A _5188_/B _5220_/B1 hold997/X vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__a22o_1
X_6189_ _6191_/A _6191_/B vssd1 vssd1 vccd1 vccd1 _6192_/A sky130_fd_sc_hd__and2_1
Xhold1531 _7734_/Q vssd1 vssd1 vccd1 vccd1 _5656_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1520 _7685_/Q vssd1 vssd1 vccd1 vccd1 hold1520/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 _7066_/Y vssd1 vssd1 vccd1 vccd1 _8505_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1553 _7682_/Q vssd1 vssd1 vccd1 vccd1 _4052_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1586 hold1799/X vssd1 vssd1 vccd1 vccd1 _4753_/B sky130_fd_sc_hd__clkbuf_2
Xhold1564 _6920_/X vssd1 vssd1 vccd1 vccd1 _8425_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1575 _4274_/X vssd1 vssd1 vccd1 vccd1 _5568_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 _4339_/X vssd1 vssd1 vccd1 vccd1 _5577_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3969__A1 _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7250__128 _8484_/CLK vssd1 vssd1 vccd1 vccd1 _8260_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5591__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5343__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5682__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3914__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5646__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4082__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4761__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3890_ _3890_/A1 _4084_/A2 _6951_/A _4084_/B2 _3889_/X vssd1 vssd1 vccd1 vccd1 _3890_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6374__A2 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5560_ _7006_/A _5560_/B vssd1 vssd1 vccd1 vccd1 _7749_/D sky130_fd_sc_hd__and2_1
X_5491_ _7512_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7680_/D sky130_fd_sc_hd__and3_1
X_4511_ _5130_/A1 _4178_/B _5442_/C vssd1 vssd1 vccd1 vccd1 _7287_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_111_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold116 _7604_/Q vssd1 vssd1 vccd1 vccd1 _5662_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _4442_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4442_/X sky130_fd_sc_hd__and2_1
XANTENNA__4700__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold105 _5673_/X vssd1 vssd1 vccd1 vccd1 _7853_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 _5668_/X vssd1 vssd1 vccd1 vccd1 _7848_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold138 _7901_/Q vssd1 vssd1 vccd1 vccd1 _5001_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _5665_/X vssd1 vssd1 vccd1 vccd1 _7845_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4373_ _4372_/A _4358_/X _5470_/C vssd1 vssd1 vccd1 vccd1 _4373_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7092_ _5389_/A _5374_/A _5409_/A vssd1 vssd1 vccd1 vccd1 _7092_/X sky130_fd_sc_hd__o21a_1
X_6112_ _6112_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6115_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ _5832_/X _5861_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6043_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5637__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7031__B _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout172_A _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7994_ _8090_/CLK hold54/X vssd1 vssd1 vccd1 vccd1 _7994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6062__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6945_ _6945_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6945_/X sky130_fd_sc_hd__and2_1
XANTENNA__4073__B1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6876_ _7017_/A _6876_/A2 _6906_/A3 _6875_/X vssd1 vssd1 vccd1 vccd1 _6876_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3820__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5486__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout437_A _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5827_ _6198_/S _5801_/X _5825_/X _5826_/Y vssd1 vssd1 vccd1 vccd1 _5827_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_9_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5758_ _5950_/S _5898_/B _5750_/Y vssd1 vssd1 vccd1 vccd1 _5759_/A sky130_fd_sc_hd__a21o_1
X_8477_ _8477_/CLK _8477_/D vssd1 vssd1 vccd1 vccd1 _8477_/Q sky130_fd_sc_hd__dfxtp_1
X_4709_ _8353_/Q _7829_/Q _7495_/Q _7463_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4709_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4610__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5689_ _5690_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _5881_/C sky130_fd_sc_hd__nor2_4
XANTENNA__5706__S _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1454_A _7302_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5325__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7428_ _8160_/CLK _7428_/D vssd1 vssd1 vccd1 vccd1 _7428_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3734__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7359_ _8456_/CLK _7359_/D vssd1 vssd1 vccd1 vccd1 _7359_/Q sky130_fd_sc_hd__dfxtp_2
Xhold672 _5653_/X vssd1 vssd1 vccd1 vccd1 _7833_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold650 _5239_/X vssd1 vssd1 vccd1 vccd1 _7447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _7825_/Q vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 _7791_/Q vssd1 vssd1 vccd1 vccd1 hold683/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _5323_/X vssd1 vssd1 vccd1 vccd1 _7554_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5628__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1361 _6812_/X vssd1 vssd1 vccd1 vccd1 _8343_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6840__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1350 _8337_/Q vssd1 vssd1 vccd1 vccd1 _6800_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4057__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1372 _6878_/X vssd1 vssd1 vccd1 vccd1 _8405_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1383 _7348_/Q vssd1 vssd1 vccd1 vccd1 _6553_/A sky130_fd_sc_hd__clkbuf_4
Xhold1394 hold1506/X vssd1 vssd1 vccd1 vccd1 _6453_/B sky130_fd_sc_hd__buf_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5677__A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5316__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6955__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output66_A _8112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4756__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6971__A _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5070__C_N _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4991_ _4990_/X _4989_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__mux2_1
X_6730_ _6955_/A _6737_/A2 _6737_/B1 hold537/X vssd1 vssd1 vccd1 vccd1 _6730_/X sky130_fd_sc_hd__a22o_1
X_3942_ _3939_/X _3940_/X _3941_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _5763_/A sky130_fd_sc_hd__o31a_1
XFILLER_0_86_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3802__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3819__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3873_ _4067_/A_N _7962_/Q vssd1 vssd1 vccd1 vccd1 _3873_/X sky130_fd_sc_hd__and2b_1
X_6661_ _6967_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6661_/X sky130_fd_sc_hd__and2_1
XFILLER_0_128_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8400_ _8468_/CLK _8400_/D vssd1 vssd1 vccd1 vccd1 _8400_/Q sky130_fd_sc_hd__dfxtp_1
X_6592_ _3837_/X _6592_/A2 _6592_/B1 hold633/X vssd1 vssd1 vccd1 vccd1 _6592_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6898__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5612_ _6961_/A _5616_/A2 _5616_/B1 hold507/X vssd1 vssd1 vccd1 vccd1 _5612_/X sky130_fd_sc_hd__a22o_1
X_5543_ _5543_/A _7090_/A vssd1 vssd1 vccd1 vccd1 _7732_/D sky130_fd_sc_hd__nor2_1
X_8331_ _8461_/CLK _8331_/D vssd1 vssd1 vccd1 vccd1 _8331_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3835__A _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7127__5 _8485_/CLK vssd1 vssd1 vccd1 vccd1 _7504_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__5307__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8262_ _8326_/CLK _8262_/D vssd1 vssd1 vccd1 vccd1 _8262_/Q sky130_fd_sc_hd__dfxtp_1
X_5474_ _5474_/A _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7663_/D sky130_fd_sc_hd__and3_1
XFILLER_0_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4425_ _4425_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3869__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8193_ _8350_/CLK _8193_/D vssd1 vssd1 vccd1 vccd1 _8193_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout404 hold1746/X vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__buf_8
X_4356_ _8488_/Q _4356_/B vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout426 _7283_/Q vssd1 vssd1 vccd1 vccd1 _3923_/B sky130_fd_sc_hd__clkbuf_8
Xfanout448 _4775_/A vssd1 vssd1 vccd1 vccd1 _7007_/A sky130_fd_sc_hd__buf_4
Xfanout415 _7063_/A vssd1 vssd1 vccd1 vccd1 _5089_/A sky130_fd_sc_hd__buf_8
XANTENNA__6865__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 _6660_/A1 vssd1 vssd1 vccd1 vccd1 _7027_/A sky130_fd_sc_hd__clkbuf_4
X_7075_ _7075_/A _7079_/B _7079_/C vssd1 vssd1 vccd1 vccd1 _8510_/D sky130_fd_sc_hd__and3_1
XANTENNA__5086__A2 _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout459 _6660_/A1 vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__clkbuf_8
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout387_A _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4287_ _4277_/Y _4281_/B _4278_/Y vssd1 vssd1 vccd1 vccd1 _4288_/B sky130_fd_sc_hd__o21a_1
X_6026_ _6028_/S _6026_/B vssd1 vssd1 vccd1 vccd1 _6026_/X sky130_fd_sc_hd__or2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6822__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6881__A _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _8019_/CLK sky130_fd_sc_hd__clkbuf_16
X_7977_ _7977_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 _7977_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6586__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6928_ _7007_/A _6928_/A2 _6943_/B _6927_/X vssd1 vssd1 vccd1 vccd1 _6928_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6859_ _6925_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6859_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4692__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5010__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8529_ _8529_/A _7092_/X vssd1 vssd1 vccd1 vccd1 _8529_/Z sky130_fd_sc_hd__ebufn_1
XANTENNA__3745__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4340__S _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold480 _5258_/X vssd1 vssd1 vccd1 vccd1 _7466_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 _7810_/Q vssd1 vssd1 vccd1 vccd1 hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6274__A1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6791__A _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1191 _8353_/Q vssd1 vssd1 vccd1 vccd1 _6832_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_84_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _8033_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1180 _5038_/X vssd1 vssd1 vccd1 vccd1 _7331_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4037__B1 _3676_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6121__S1 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6577__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output104_A _7299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3941__A_N _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4210_ _4208_/Y _4210_/B vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__5870__A _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5190_ _6777_/A _5221_/A2 _5221_/B1 hold543/X vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__a22o_1
X_4141_ _6405_/A _4121_/X _4140_/X _4118_/Y vssd1 vssd1 vccd1 vccd1 _4141_/Y sky130_fd_sc_hd__o211ai_2
XANTENNA__6804__A3 _6776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5699__S0 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4072_ _4759_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _4072_/X sky130_fd_sc_hd__and2_1
X_7900_ _8507_/CLK _7900_/D vssd1 vssd1 vccd1 vccd1 _7900_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_75_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _8494_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4028__B1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6568__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7831_ _8355_/CLK _7831_/D vssd1 vssd1 vccd1 vccd1 _7831_/Q sky130_fd_sc_hd__dfxtp_1
X_4974_ _4972_/X _4973_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__mux2_1
X_7762_ _8091_/CLK _7762_/D vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5240__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6713_ _6921_/A _6705_/B _6738_/B1 hold773/X vssd1 vssd1 vccd1 vccd1 _6713_/X sky130_fd_sc_hd__a22o_1
X_3925_ _4744_/B _3966_/B vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__and2_1
XFILLER_0_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7693_ _8086_/CLK _7693_/D vssd1 vssd1 vccd1 vccd1 _7693_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4674__S1 _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6644_ _7028_/A _6644_/A2 _6666_/A3 _6643_/X vssd1 vssd1 vccd1 vccd1 _6644_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_132_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3856_ _3856_/A0 _3855_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6242_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_6_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6575_ _6937_/A _6592_/A2 _6592_/B1 hold681/X vssd1 vssd1 vccd1 vccd1 _6575_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3787_ _3787_/A _3787_/B vssd1 vssd1 vccd1 vccd1 _3788_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4160__S _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5526_ _8245_/Q _5538_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7715_/D sky130_fd_sc_hd__and3_1
X_8314_ _8440_/CLK _8314_/D vssd1 vssd1 vccd1 vccd1 _8314_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8245_ _8245_/CLK _8245_/D vssd1 vssd1 vccd1 vccd1 _8245_/Q sky130_fd_sc_hd__dfxtp_1
X_5457_ _5457_/A _5503_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__and3_1
XFILLER_0_112_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5700__A0 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4408_ _5036_/A1 _5067_/S _4406_/X _4407_/Y vssd1 vssd1 vccd1 vccd1 _8374_/D sky130_fd_sc_hd__a22o_1
X_8176_ _8332_/CLK _8176_/D vssd1 vssd1 vccd1 vccd1 _8176_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout223 _7073_/B vssd1 vssd1 vccd1 vccd1 _5542_/C sky130_fd_sc_hd__buf_4
X_5388_ _6553_/A _5389_/A _5388_/C vssd1 vssd1 vccd1 vccd1 _5388_/X sky130_fd_sc_hd__or3_2
Xfanout201 _6028_/S vssd1 vssd1 vccd1 vccd1 _6302_/A sky130_fd_sc_hd__buf_4
Xfanout212 _5538_/C vssd1 vssd1 vccd1 vccd1 _5541_/C sky130_fd_sc_hd__buf_4
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout256 _5584_/Y vssd1 vssd1 vccd1 vccd1 _5617_/B1 sky130_fd_sc_hd__clkbuf_8
X_4339_ _4339_/A _4339_/B vssd1 vssd1 vccd1 vccd1 _4339_/X sky130_fd_sc_hd__xor2_1
Xfanout245 _6774_/B1 vssd1 vssd1 vccd1 vccd1 _6773_/B1 sky130_fd_sc_hd__buf_8
Xfanout234 _5182_/A2 vssd1 vssd1 vccd1 vccd1 _4407_/B sky130_fd_sc_hd__buf_2
Xfanout278 _6971_/B vssd1 vssd1 vccd1 vccd1 _6963_/B sky130_fd_sc_hd__buf_8
Xfanout267 _4084_/A2 vssd1 vssd1 vccd1 vccd1 _4073_/A2 sky130_fd_sc_hd__buf_6
XANTENNA__6256__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 _6703_/Y vssd1 vssd1 vccd1 vccd1 _6737_/A2 sky130_fd_sc_hd__buf_8
X_7058_ _7071_/B _7057_/Y _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8501_/D sky130_fd_sc_hd__a21oi_1
X_6009_ _6128_/A _6307_/B _6309_/B _5759_/A vssd1 vssd1 vccd1 vccd1 _6009_/X sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_66_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _7977_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_69_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1786_A _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3793__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6731__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_57_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _8368_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4753__B _4753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4656__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3710_/A0 _3709_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6295_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_125_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4690_ _4688_/X _4689_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4690_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5584__B _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6183__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6722__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6360_ _5739_/Y _6067_/X _6359_/X _6251_/A vssd1 vssd1 vccd1 vccd1 _6360_/X sky130_fd_sc_hd__o22a_1
X_5311_ _6929_/A _5332_/A2 _5332_/B1 hold413/X vssd1 vssd1 vccd1 vccd1 _5311_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5289__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6291_ _6008_/A _5718_/X _6130_/X _6287_/X vssd1 vssd1 vccd1 vccd1 _6292_/D sky130_fd_sc_hd__a31o_1
X_8030_ _8030_/CLK _8030_/D vssd1 vssd1 vccd1 vccd1 _8030_/Q sky130_fd_sc_hd__dfxtp_1
X_5242_ _6937_/A _5226_/B _5259_/B1 hold489/X vssd1 vssd1 vccd1 vccd1 _5242_/X sky130_fd_sc_hd__a22o_1
X_5173_ hold63/X _5468_/C vssd1 vssd1 vccd1 vccd1 _5173_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5105__A _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6238__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4124_ _6157_/A _6154_/A vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__and2b_1
Xinput1 i_instr_ID[10] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_1
XFILLER_0_127_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4055_ _3923_/B _7951_/Q vssd1 vssd1 vccd1 vccd1 _4055_/X sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_48_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8080_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5997__A0 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4895__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7814_ _8332_/CLK _7814_/D vssd1 vssd1 vccd1 vccd1 _7814_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5749__A0 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4647__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5213__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7204__82 _8451_/CLK vssd1 vssd1 vccd1 vccd1 _8117_/CLK sky130_fd_sc_hd__inv_2
X_4957_ _4956_/X _4953_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8255_/D sky130_fd_sc_hd__mux2_1
X_7745_ _8387_/CLK _7745_/D vssd1 vssd1 vccd1 vccd1 _7745_/Q sky130_fd_sc_hd__dfxtp_1
X_7676_ _8517_/CLK _7676_/D vssd1 vssd1 vccd1 vccd1 _7676_/Q sky130_fd_sc_hd__dfxtp_1
X_3908_ _5846_/A _6302_/A vssd1 vssd1 vccd1 vccd1 _3910_/A sky130_fd_sc_hd__nand2_1
X_4888_ _8342_/Q _7818_/Q _7484_/Q _7452_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4888_/X sky130_fd_sc_hd__mux4_1
X_6627_ _6933_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6627_/X sky130_fd_sc_hd__and2_1
X_3839_ _3839_/A1 _4073_/A2 _6971_/A _4073_/B2 _3838_/X vssd1 vssd1 vccd1 vccd1 _6452_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_62_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5494__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6713__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6558_ _6558_/A _6776_/B vssd1 vssd1 vccd1 vccd1 _6560_/B sky130_fd_sc_hd__or2_1
XFILLER_0_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6489_ _7006_/A _6489_/B vssd1 vssd1 vccd1 vccd1 _6489_/X sky130_fd_sc_hd__and2_1
XANTENNA__5714__S _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5509_ _7530_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7698_/D sky130_fd_sc_hd__and3_1
X_8228_ _8442_/CLK _8228_/D vssd1 vssd1 vccd1 vccd1 _8228_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4583__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8159_ _8442_/CLK _8159_/D vssd1 vssd1 vccd1 vccd1 _8159_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_39_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _7805_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5988__B1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5204__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5685__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3766__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6165__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3933__A _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6963__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6455__S _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5979__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4764__A _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4877__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6640__A1 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6079__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5860_ _5744_/X _5781_/X _5860_/S vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__mux2_1
X_4811_ _8331_/Q _7807_/Q _7473_/Q _7441_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4811_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4629__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5791_ _5792_/B vssd1 vssd1 vccd1 vccd1 _5791_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5746__A3 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4742_ _4741_/X _4740_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__mux2_1
X_7530_ _7530_/CLK _7530_/D vssd1 vssd1 vccd1 vccd1 _7530_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4673_ _4672_/X _4669_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7521_/D sky130_fd_sc_hd__mux2_1
X_7461_ _8481_/CLK _7461_/D vssd1 vssd1 vccd1 vccd1 _7461_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3827__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6412_ _6123_/X _6411_/X _6412_/S vssd1 vssd1 vccd1 vccd1 _6412_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7392_ _8378_/CLK _7392_/D vssd1 vssd1 vccd1 vccd1 _7392_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4801__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6343_ _5740_/Y _6042_/Y _6342_/X _6309_/A vssd1 vssd1 vccd1 vccd1 _6343_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3843__A _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6274_ _6309_/A _5954_/Y _6271_/X _6273_/X vssd1 vssd1 vccd1 vccd1 _6274_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4565__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5225_ _6740_/C _6776_/A vssd1 vssd1 vccd1 vccd1 _5227_/B sky130_fd_sc_hd__or2_1
X_8013_ _8465_/CLK _8013_/D vssd1 vssd1 vccd1 vccd1 _8013_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__7034__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1702 _3941_/X vssd1 vssd1 vccd1 vccd1 _6422_/A3 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1735 _7596_/Q vssd1 vssd1 vccd1 vccd1 _5732_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1713 _8493_/Q vssd1 vssd1 vccd1 vccd1 _3722_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_5156_ _5156_/A1 _4416_/B _5166_/B1 _5155_/X vssd1 vssd1 vccd1 vccd1 _7390_/D sky130_fd_sc_hd__o211a_1
XANTENNA__6873__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1724 _8496_/Q vssd1 vssd1 vccd1 vccd1 _3880_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1746 _7359_/Q vssd1 vssd1 vccd1 vccd1 hold1746/X sky130_fd_sc_hd__buf_2
X_5087_ _7065_/A _5451_/C vssd1 vssd1 vccd1 vccd1 _5087_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4107_ _5971_/A _5974_/A _4045_/D _4041_/Y _5993_/A vssd1 vssd1 vccd1 vccd1 _4107_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA_fanout467_A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1768 _6096_/A vssd1 vssd1 vccd1 vccd1 _6110_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1757 _7728_/Q vssd1 vssd1 vccd1 vccd1 _3819_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4038_ _4753_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _4038_/X sky130_fd_sc_hd__and2_1
XANTENNA__4868__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1779 _7715_/Q vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7050__A _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5198__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5989_ _5979_/X _5980_/X _5987_/X _5988_/Y vssd1 vssd1 vccd1 vccd1 _5989_/X sky130_fd_sc_hd__o31a_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5709__S _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4613__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7728_ _8419_/CLK _7728_/D vssd1 vssd1 vccd1 vccd1 _7728_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1484_A _7298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3737__B _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7659_ _8360_/CLK _7659_/D vssd1 vssd1 vccd1 vccd1 _7659_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6698__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7055__C_N _7031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3920__A2 _3917_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5122__A1 input23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4556__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6870__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6622__A1 _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3987__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3739__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7195__73 _8515_/CLK vssd1 vssd1 vccd1 vccd1 _8108_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_65_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6233__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6689__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold309 _5437_/X vssd1 vssd1 vccd1 vccd1 _7626_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5361__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4759__A _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _4442_/A _5069_/S _5182_/B1 _5009_/X vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__o211a_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1009 _8456_/Q vssd1 vssd1 vccd1 vccd1 _6998_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6961_ _6961_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6961_/X sky130_fd_sc_hd__and2_1
XFILLER_0_88_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5912_ _6302_/A _6083_/A _5907_/X _5911_/Y _5786_/B vssd1 vssd1 vccd1 vccd1 _5912_/X
+ sky130_fd_sc_hd__o32a_1
X_6892_ _7022_/A _6892_/A2 _6906_/A3 _6891_/X vssd1 vssd1 vccd1 vccd1 _6892_/X sky130_fd_sc_hd__a31o_1
X_5843_ _6342_/S _5971_/B vssd1 vssd1 vccd1 vccd1 _5846_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3838__A _4775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7513_ _7513_/CLK _7513_/D vssd1 vssd1 vccd1 vccd1 _7513_/Q sky130_fd_sc_hd__dfxtp_1
X_5774_ _6302_/A _5774_/B vssd1 vssd1 vccd1 vccd1 _6163_/B sky130_fd_sc_hd__or2_1
XANTENNA__6392__A3 _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8493_ _8501_/CLK _8493_/D vssd1 vssd1 vccd1 vccd1 _8493_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4725_ _4723_/X _4724_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7444_ _8136_/CLK _7444_/D vssd1 vssd1 vccd1 vccd1 _7444_/Q sky130_fd_sc_hd__dfxtp_1
X_4656_ _8185_/Q _8217_/Q _8281_/Q _7789_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4656_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout215_A _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4786__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold821 _7413_/Q vssd1 vssd1 vccd1 vccd1 hold821/X sky130_fd_sc_hd__dlygate4sd3_1
X_4587_ _8465_/Q _8397_/Q _8429_/Q _8303_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4587_/X sky130_fd_sc_hd__mux4_1
Xhold810 _5207_/X vssd1 vssd1 vccd1 vccd1 _7421_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7375_ _8362_/CLK _7375_/D vssd1 vssd1 vccd1 vccd1 _7375_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5888__C1 _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5352__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5491__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3902__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold843 _8149_/Q vssd1 vssd1 vccd1 vccd1 hold843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 _5614_/X vssd1 vssd1 vccd1 vccd1 _7798_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6326_ _3725_/B _6414_/B1 _6398_/B1 _6315_/A _6292_/A vssd1 vssd1 vccd1 vccd1 _6326_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold854 _6761_/X vssd1 vssd1 vccd1 vccd1 _8312_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold865 _7538_/Q vssd1 vssd1 vccd1 vccd1 hold865/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 _5351_/X vssd1 vssd1 vccd1 vccd1 _7578_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 _7829_/Q vssd1 vssd1 vccd1 vccd1 hold887/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 _5328_/X vssd1 vssd1 vccd1 vccd1 _7559_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4538__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6257_ _3859_/B _6292_/A _6347_/B1 vssd1 vssd1 vccd1 vccd1 _6257_/Y sky130_fd_sc_hd__a21oi_1
Xhold1510 _4155_/Y vssd1 vssd1 vccd1 vccd1 hold1510/X sky130_fd_sc_hd__buf_4
X_6188_ _6188_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6191_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__6852__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5208_ _6945_/A _5188_/B _5220_/B1 hold833/X vssd1 vssd1 vccd1 vccd1 _5208_/X sky130_fd_sc_hd__a22o_1
Xhold1521 _6438_/Y vssd1 vssd1 vccd1 vccd1 _7920_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1532 hold1796/X vssd1 vssd1 vccd1 vccd1 _4756_/B sky130_fd_sc_hd__clkbuf_2
X_5139_ _5449_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__or2_1
Xhold1543 _7697_/Q vssd1 vssd1 vccd1 vccd1 _3829_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6604__A1 _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1576 _7365_/Q vssd1 vssd1 vccd1 vccd1 _7083_/B2 sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_66_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1565 _7347_/Q vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__buf_2
Xhold1554 _4052_/X vssd1 vssd1 vccd1 vccd1 _6435_/B sky130_fd_sc_hd__buf_1
Xhold1587 _7671_/Q vssd1 vssd1 vccd1 vccd1 _3904_/A1 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold1598 _7631_/Q vssd1 vssd1 vccd1 vccd1 _4156_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3969__A2 _3967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4710__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__8026__D _8026_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3748__A _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5040__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5591__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6215__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5343__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4777__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5646__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3930__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6071__A2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4082__A1 _4757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4761__B _4761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6034__A _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6374__A3 _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6969__A _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4510_ _5132_/A1 _4440_/B _5442_/C vssd1 vssd1 vccd1 vccd1 _7288_/D sky130_fd_sc_hd__mux2_1
X_5490_ _7511_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7679_/D sky130_fd_sc_hd__and3_1
XFILLER_0_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold117 _5662_/X vssd1 vssd1 vccd1 vccd1 _7842_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ hold212/X _4440_/Y _5442_/C vssd1 vssd1 vccd1 vccd1 _8362_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold106 _7618_/Q vssd1 vssd1 vccd1 vccd1 _5676_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _5001_/X vssd1 vssd1 vccd1 vccd1 _7283_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5885__A2 _5739_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold128 _7867_/Q vssd1 vssd1 vccd1 vccd1 _6488_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7087__A1 _5544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6111_ _6106_/X _6109_/Y _6111_/B1 _7029_/A vssd1 vssd1 vccd1 vccd1 _6111_/X sky130_fd_sc_hd__o211a_1
X_4372_ _4372_/A _4372_/B vssd1 vssd1 vccd1 vccd1 _4372_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4001__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7087__B2 _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7091_ _5389_/A _5374_/A _5409_/A vssd1 vssd1 vccd1 vccd1 _7091_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5098__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6042_ _6302_/A _6040_/X _6041_/X _5740_/B vssd1 vssd1 vccd1 vccd1 _6042_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__6834__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5637__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A _7077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6209__A _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4940__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7993_ _8379_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _7993_/Q sky130_fd_sc_hd__dfxtp_1
X_6944_ _6877_/A _6963_/B _6944_/B1 _7015_/A vssd1 vssd1 vccd1 vccd1 _6944_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6062__A2 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout165_A _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5270__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4073__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6875_ _6941_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6875_/X sky130_fd_sc_hd__and2_1
XANTENNA__3820__B2 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3820__A1 _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5022__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5826_ _3922_/B _6380_/A _5823_/Y _5734_/A vssd1 vssd1 vccd1 vccd1 _5826_/Y sky130_fd_sc_hd__o22ai_1
XANTENNA__5486__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout332_A _3875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5757_ _5804_/A _5838_/B _5752_/X vssd1 vssd1 vccd1 vccd1 _5898_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__4376__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6770__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6879__A _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8476_ _8476_/CLK _8476_/D vssd1 vssd1 vccd1 vccd1 _8476_/Q sky130_fd_sc_hd__dfxtp_1
X_4708_ _4707_/X _4704_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7526_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5688_ _5688_/A _7596_/Q _8453_/Q vssd1 vssd1 vccd1 vccd1 _5730_/B sky130_fd_sc_hd__or3b_2
X_7427_ _8486_/CLK _7427_/D vssd1 vssd1 vccd1 vccd1 _7427_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5325__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4639_ _8343_/Q _7819_/Q _7485_/Q _7453_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4639_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_8_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold651 _7778_/Q vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 _5211_/X vssd1 vssd1 vccd1 vccd1 _7425_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7358_ _8032_/CLK _7358_/D vssd1 vssd1 vccd1 vccd1 _7358_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_13_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold662 _5645_/X vssd1 vssd1 vccd1 vccd1 _7825_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 _7804_/Q vssd1 vssd1 vccd1 vccd1 hold695/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 _5607_/X vssd1 vssd1 vccd1 vccd1 _7791_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7289_ _8358_/CLK _7289_/D _7099_/Y vssd1 vssd1 vccd1 vccd1 _7289_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5007__B _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6309_ _6309_/A _6309_/B vssd1 vssd1 vccd1 vccd1 _6309_/Y sky130_fd_sc_hd__nor2_2
Xhold673 _7424_/Q vssd1 vssd1 vccd1 vccd1 hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5628__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1351 _6800_/X vssd1 vssd1 vccd1 vccd1 _8337_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4931__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1340 _8333_/Q vssd1 vssd1 vccd1 vccd1 _6792_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 _8335_/Q vssd1 vssd1 vccd1 vccd1 _6796_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1373 _8328_/Q vssd1 vssd1 vccd1 vccd1 _6782_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 _5389_/X vssd1 vssd1 vccd1 vccd1 _7079_/C sky130_fd_sc_hd__buf_4
XANTENNA__6589__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1395 _8380_/Q vssd1 vssd1 vccd1 vccd1 _4389_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6789__A _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6761__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7165__43 _8011_/CLK vssd1 vssd1 vccd1 vccd1 _8045_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_51_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3925__B _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5316__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6816__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4756__B _4756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6971__B _6971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5868__A _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4772__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4990_ _8486_/Q _8418_/Q _8450_/Q _8324_/Q _4990_/S0 _4990_/S1 vssd1 vssd1 vccd1
+ vccd1 _4990_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5252__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3941_ _4083_/B _3941_/B _3941_/C vssd1 vssd1 vccd1 vccd1 _3941_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6660_ _6660_/A1 _6660_/A2 _6666_/A3 _6659_/X vssd1 vssd1 vccd1 vccd1 _6660_/X sky130_fd_sc_hd__a31o_1
X_3872_ _3872_/A _3872_/B vssd1 vssd1 vccd1 vccd1 _3896_/B sky130_fd_sc_hd__and2_1
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6752__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5611_ _6959_/A _5616_/A2 _5616_/B1 hold879/X vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6591_ _6969_/A _6559_/B _6591_/B1 hold963/X vssd1 vssd1 vccd1 vccd1 _6591_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4989__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5542_ _8261_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7731_/D sky130_fd_sc_hd__and3_1
XANTENNA__5807__S _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4711__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8330_ _8350_/CLK _8330_/D vssd1 vssd1 vccd1 vccd1 _8330_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5307__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5473_ _5473_/A _7088_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _7662_/D sky130_fd_sc_hd__and3_1
X_8261_ _8261_/CLK _8261_/D vssd1 vssd1 vccd1 vccd1 _8261_/Q sky130_fd_sc_hd__dfxtp_1
X_4424_ _4427_/A _4427_/B _4504_/A1 vssd1 vssd1 vccd1 vccd1 _4424_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3869__A1 _4764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8192_ _8483_/CLK _8192_/D vssd1 vssd1 vccd1 vccd1 _8192_/Q sky130_fd_sc_hd__dfxtp_1
X_4355_ _4352_/A _4351_/X _4350_/B vssd1 vssd1 vccd1 vccd1 _4357_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout405 _4976_/S1 vssd1 vssd1 vccd1 vccd1 _4990_/S1 sky130_fd_sc_hd__clkbuf_8
X_7074_ _7074_/A _7079_/B _7079_/C vssd1 vssd1 vccd1 vccd1 _8509_/D sky130_fd_sc_hd__and3_1
Xfanout427 _7028_/A vssd1 vssd1 vccd1 vccd1 _7018_/A sky130_fd_sc_hd__buf_4
Xfanout416 _7063_/A vssd1 vssd1 vccd1 vccd1 _4990_/S0 sky130_fd_sc_hd__buf_4
Xfanout438 _6551_/A vssd1 vssd1 vccd1 vccd1 _6550_/A sky130_fd_sc_hd__clkbuf_4
Xfanout449 _6706_/A vssd1 vssd1 vccd1 vccd1 _7010_/A sky130_fd_sc_hd__buf_4
XANTENNA__7042__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4284_/Y _4286_/B vssd1 vssd1 vccd1 vccd1 _4286_/Y sky130_fd_sc_hd__nand2b_1
X_6025_ _5934_/X _6024_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6026_/B sky130_fd_sc_hd__mux2_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4913__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6881__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7976_ _8361_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 _7976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5497__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5243__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6927_ _6927_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6927_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6858_ _7005_/A _6858_/A2 _6906_/A3 _6857_/X vssd1 vssd1 vccd1 vccd1 _6858_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_134_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5809_ _5807_/X _5808_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5810_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6789_ _6921_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6789_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8528_ _8528_/A _7091_/X vssd1 vssd1 vccd1 vccd1 _8528_/Z sky130_fd_sc_hd__ebufn_1
XANTENNA__5717__S _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8459_ _8468_/CLK _8459_/D vssd1 vssd1 vccd1 vccd1 _8459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold470 _6672_/X vssd1 vssd1 vccd1 vccd1 _8199_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _7454_/Q vssd1 vssd1 vccd1 vccd1 hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _5630_/X vssd1 vssd1 vccd1 vccd1 _7810_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6791__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1170 _6824_/X vssd1 vssd1 vccd1 vccd1 _8349_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1181 _8167_/Q vssd1 vssd1 vccd1 vccd1 _6606_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 _6832_/X vssd1 vssd1 vccd1 vccd1 _8353_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5234__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4037__A1 _4753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4037__B2 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6409__S0 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3936__A _7282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6734__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6458__S _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4140_ _4134_/X _4138_/X _4139_/Y _3897_/C vssd1 vssd1 vccd1 vccd1 _4140_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5699__S1 _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4071_ _4759_/B _4071_/A2 _4071_/B1 _4069_/X _4070_/X vssd1 vssd1 vccd1 vccd1 _6115_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_116_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7830_ _8354_/CLK _7830_/D vssd1 vssd1 vccd1 vccd1 _7830_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4028__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4973_ _8161_/Q _7560_/Q _7432_/Q _7592_/Q _7063_/A _4976_/S1 vssd1 vssd1 vccd1 vccd1
+ _4973_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6206__B _6406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7761_ _8379_/CLK _7761_/D vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
X_3924_ _8067_/Q _3677_/Y _4079_/B1 _8003_/Q _3923_/X vssd1 vssd1 vccd1 vccd1 _6909_/A
+ sky130_fd_sc_hd__a221o_2
XANTENNA__4007__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6712_ _6853_/A _6705_/B _6738_/B1 hold435/X vssd1 vssd1 vccd1 vccd1 _6712_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7692_ _8195_/CLK _7692_/D vssd1 vssd1 vccd1 vccd1 _7692_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6643_ _6949_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6643_/X sky130_fd_sc_hd__and2_1
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3855_ _3855_/A1 _4084_/A2 _3851_/X _4084_/B2 _3854_/X vssd1 vssd1 vccd1 vccd1 _3855_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6725__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6574_ _6935_/A _6592_/A2 _6592_/B1 _6574_/B2 vssd1 vssd1 vccd1 vccd1 _6574_/X sky130_fd_sc_hd__a22o_1
X_3786_ _6175_/A _6172_/A vssd1 vssd1 vccd1 vccd1 _3787_/B sky130_fd_sc_hd__or2_1
XFILLER_0_131_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5525_ _8244_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7714_/D sky130_fd_sc_hd__and3_1
X_8313_ _8475_/CLK _8313_/D vssd1 vssd1 vccd1 vccd1 _8313_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8244_ _8244_/CLK _8244_/D vssd1 vssd1 vccd1 vccd1 _8244_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5456_ _5456_/A _5540_/B _5456_/C vssd1 vssd1 vccd1 vccd1 _5456_/X sky130_fd_sc_hd__and3_1
X_4407_ _4407_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _4407_/Y sky130_fd_sc_hd__nor2_1
X_8175_ _8175_/CLK _8175_/D vssd1 vssd1 vccd1 vccd1 _8175_/Q sky130_fd_sc_hd__dfxtp_1
X_5387_ _6553_/A _5389_/A _5388_/C vssd1 vssd1 vccd1 vccd1 _6976_/A sky130_fd_sc_hd__nor3_1
Xfanout202 _3907_/Y vssd1 vssd1 vccd1 vccd1 _6028_/S sky130_fd_sc_hd__buf_4
Xfanout213 _7073_/B vssd1 vssd1 vccd1 vccd1 _5538_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout224 _7073_/B vssd1 vssd1 vccd1 vccd1 _5523_/C sky130_fd_sc_hd__buf_4
Xfanout246 _6741_/Y vssd1 vssd1 vccd1 vccd1 _6774_/B1 sky130_fd_sc_hd__buf_8
X_4338_ _4328_/Y _4332_/B _4330_/B vssd1 vssd1 vccd1 vccd1 _4339_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout235 _5182_/A2 vssd1 vssd1 vccd1 vccd1 _5067_/S sky130_fd_sc_hd__clkbuf_8
Xfanout268 _3708_/Y vssd1 vssd1 vccd1 vccd1 _4084_/A2 sky130_fd_sc_hd__buf_8
Xfanout279 _6845_/B vssd1 vssd1 vccd1 vccd1 _6906_/A3 sky130_fd_sc_hd__buf_8
Xfanout257 _5335_/Y vssd1 vssd1 vccd1 vccd1 _5367_/B1 sky130_fd_sc_hd__buf_6
X_7057_ _7057_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7057_/Y sky130_fd_sc_hd__nand2_1
X_4269_ _4410_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4407_/A sky130_fd_sc_hd__and2_1
X_6008_ _6008_/A _6008_/B vssd1 vssd1 vccd1 vccd1 _6309_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4616__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5216__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7959_ _8020_/CLK hold93/X vssd1 vssd1 vccd1 vccd1 _7959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3778__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6716__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7873__D _7873_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7135__13 _8338_/CLK vssd1 vssd1 vccd1 vccd1 _7512_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7223__101 _8339_/CLK vssd1 vssd1 vccd1 vccd1 _8233_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_20_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6798__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3789__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5207__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4526__S _7365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6970__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6707__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4261__S _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5310_ _6927_/A _5332_/A2 _5332_/B1 _5310_/B2 vssd1 vssd1 vccd1 vccd1 _5310_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6290_ _6270_/A _6309_/A _5881_/C _6126_/A vssd1 vssd1 vccd1 vccd1 _6292_/C sky130_fd_sc_hd__o211a_1
X_5241_ _6935_/A _5226_/B _5259_/B1 _5241_/B2 vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_53_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5172_ _5172_/A1 _5067_/S _5172_/B1 _5171_/X vssd1 vssd1 vccd1 vccd1 _7398_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5105__B _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4123_ _6175_/A _6172_/A vssd1 vssd1 vccd1 vccd1 _4123_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput2 i_instr_ID[11] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_1
X_4054_ _6096_/A _6094_/A vssd1 vssd1 vccd1 vccd1 _4090_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_127_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5997__A1 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5121__A _7031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5749__A1 _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7813_ _8467_/CLK _7813_/D vssd1 vssd1 vccd1 vccd1 _7813_/Q sky130_fd_sc_hd__dfxtp_1
X_7744_ _8362_/CLK _7744_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4956_ _4955_/X _4954_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout245_A _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3907_ _3968_/A _3904_/Y _3905_/Y vssd1 vssd1 vccd1 vccd1 _3907_/Y sky130_fd_sc_hd__o21ai_2
X_7675_ _8173_/CLK _7675_/D vssd1 vssd1 vccd1 vccd1 _7675_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7048__A _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4887_ _4886_/X _4883_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8245_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout412_A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3838_ _4775_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3838_/X sky130_fd_sc_hd__and2_1
X_6626_ _7023_/A _6626_/A2 _6666_/A3 _6625_/X vssd1 vssd1 vccd1 vccd1 _6626_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5494__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6557_ _6558_/A _6776_/B vssd1 vssd1 vccd1 vccd1 _6557_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6887__A _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3769_ _4761_/B _3676_/A _4082_/B1 _3767_/X _3768_/X vssd1 vssd1 vccd1 vccd1 _6157_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_70_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5508_ _7529_/Q _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _7697_/D sky130_fd_sc_hd__and3_1
X_6488_ _6520_/A _6488_/B vssd1 vssd1 vccd1 vccd1 _6488_/X sky130_fd_sc_hd__and2_1
XFILLER_0_42_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5439_ _5439_/A _5470_/B _5470_/C vssd1 vssd1 vccd1 vccd1 _5439_/X sky130_fd_sc_hd__and3_1
X_8227_ _8350_/CLK _8227_/D vssd1 vssd1 vccd1 vccd1 _8227_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4583__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5780__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8158_ _8481_/CLK _8158_/D vssd1 vssd1 vccd1 vccd1 _8158_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5015__B _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7109_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7109_/Y sky130_fd_sc_hd__inv_2
X_8089_ _8501_/CLK _8123_/D vssd1 vssd1 vccd1 vccd1 _8089_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3999__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6952__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6797__A _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5140__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4764__B _4764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6079__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _4809_/X _4806_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8234_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5600__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5790_ _5838_/A _5789_/X _4093_/Y vssd1 vssd1 vccd1 vccd1 _5792_/B sky130_fd_sc_hd__o21bai_1
XANTENNA__3837__S0 _7282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4741_ _8487_/Q _8419_/Q _8451_/Q _8325_/Q _4741_/S0 _4741_/S1 vssd1 vssd1 vccd1
+ vccd1 _4741_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4672_ _4671_/X _4670_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7460_ _8160_/CLK _7460_/D vssd1 vssd1 vccd1 vccd1 _7460_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6411_ _6270_/B _6410_/X _6411_/S vssd1 vssd1 vccd1 vccd1 _6411_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7391_ _8071_/CLK _7391_/D vssd1 vssd1 vccd1 vccd1 _7391_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6500__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6342_ _6196_/X _6341_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6342_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6273_ _6126_/A _5881_/C _5793_/Y _5962_/X _6412_/S vssd1 vssd1 vccd1 vccd1 _6273_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5224_ _6740_/C _6776_/A vssd1 vssd1 vccd1 vccd1 _5224_/Y sky130_fd_sc_hd__nor2_1
X_8012_ _8479_/CLK _8012_/D vssd1 vssd1 vccd1 vccd1 _8012_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4565__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1725 _8100_/Q vssd1 vssd1 vccd1 vccd1 hold1725/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1714 _8454_/Q vssd1 vssd1 vccd1 vccd1 _5688_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1703 _6422_/X vssd1 vssd1 vccd1 vccd1 _7904_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5155_ _5457_/A _5540_/C vssd1 vssd1 vccd1 vccd1 _5155_/X sky130_fd_sc_hd__or2_1
X_4106_ _6016_/A _6013_/A vssd1 vssd1 vccd1 vccd1 _4106_/Y sky130_fd_sc_hd__nand2b_1
X_5086_ input4/X _5085_/B _5140_/B1 _5085_/Y vssd1 vssd1 vccd1 vccd1 _7355_/D sky130_fd_sc_hd__o211a_1
Xhold1769 _6110_/X vssd1 vssd1 vccd1 vccd1 _6111_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1736 _4149_/X vssd1 vssd1 vccd1 vccd1 _5742_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1758 _7726_/Q vssd1 vssd1 vccd1 vccd1 _3718_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1747 _7357_/Q vssd1 vssd1 vccd1 vccd1 hold1747/X sky130_fd_sc_hd__clkbuf_4
XANTENNA__5489__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4037_ _4753_/B _3669_/Y _3676_/Y _6927_/A _4036_/X vssd1 vssd1 vccd1 vccd1 _5993_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__7050__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5786__A _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5198__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5988_ _5988_/A1 _6011_/A2 _6911_/A vssd1 vssd1 vccd1 vccd1 _5988_/Y sky130_fd_sc_hd__a21oi_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6395__A1 _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6934__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4939_ _4937_/X _4938_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__mux2_1
X_7727_ _8195_/CLK _7727_/D vssd1 vssd1 vccd1 vccd1 _7727_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6147__A1 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7658_ _8030_/CLK _7658_/D vssd1 vssd1 vccd1 vccd1 _7658_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6609_ _6849_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6609_/X sky130_fd_sc_hd__and2_1
XANTENNA__6698__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7589_ _8413_/CLK _7589_/D vssd1 vssd1 vccd1 vccd1 _7589_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5122__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4556__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6783__C _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5830__A0 _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6689__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6233__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5361__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output89_A _8104_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5649__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6310__A1 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4775__A _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6960_ _7023_/A _6960_/A2 _6970_/A3 _6959_/X vssd1 vssd1 vccd1 vccd1 _6960_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5911_ _5911_/A vssd1 vssd1 vccd1 vccd1 _5911_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_124_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6891_ _6891_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6891_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5842_ _5881_/C _5837_/X _5841_/X _6008_/B vssd1 vssd1 vccd1 vccd1 _5842_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4714__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6916__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5773_ _5963_/S _5797_/S _5773_/C vssd1 vssd1 vccd1 vccd1 _5774_/B sky130_fd_sc_hd__or3_1
XANTENNA__3838__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7512_ _7512_/CLK _7512_/D vssd1 vssd1 vccd1 vccd1 _7512_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_4_8_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4724_ _8162_/Q _7561_/Q _7433_/Q _7593_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4724_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_133_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8492_ _8494_/CLK _8492_/D vssd1 vssd1 vccd1 vccd1 _8492_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4655_ _4653_/X _4654_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4655_/X sky130_fd_sc_hd__mux2_1
X_7443_ _8478_/CLK _7443_/D vssd1 vssd1 vccd1 vccd1 _7443_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4786__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4586_ _8175_/Q _8207_/Q _8271_/Q _7779_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4586_/X sky130_fd_sc_hd__mux4_1
Xhold811 _7489_/Q vssd1 vssd1 vccd1 vccd1 hold811/X sky130_fd_sc_hd__dlygate4sd3_1
X_7374_ _8363_/CLK _7374_/D vssd1 vssd1 vccd1 vccd1 _7374_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout208_A _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold800 _6771_/X vssd1 vssd1 vccd1 vccd1 _8322_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput60 i_read_data_M[7] vssd1 vssd1 vccd1 vccd1 _6528_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5352__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold822 _5199_/X vssd1 vssd1 vccd1 vccd1 _7413_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold855 _8215_/Q vssd1 vssd1 vccd1 vccd1 hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 _6577_/X vssd1 vssd1 vccd1 vccd1 _8149_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6325_ _5806_/B _6362_/C _6324_/X _5740_/B vssd1 vssd1 vccd1 vccd1 _6325_/X sky130_fd_sc_hd__a22o_1
Xhold833 _7422_/Q vssd1 vssd1 vccd1 vccd1 hold833/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 _5307_/X vssd1 vssd1 vccd1 vccd1 _7538_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 _8469_/Q vssd1 vssd1 vccd1 vccd1 _7011_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 _5649_/X vssd1 vssd1 vccd1 vccd1 _7829_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4538__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold899 _7574_/Q vssd1 vssd1 vccd1 vccd1 hold899/X sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ _6391_/A _6247_/Y _6252_/X vssd1 vssd1 vccd1 vccd1 _6256_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5104__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5207_ _6877_/A _5221_/A2 _5221_/B1 hold809/X vssd1 vssd1 vccd1 vccd1 _5207_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6376__S _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1500 hold1810/X vssd1 vssd1 vccd1 vccd1 _4769_/B sky130_fd_sc_hd__buf_1
X_6187_ _3787_/A _6417_/A2 _6186_/X _6347_/B1 vssd1 vssd1 vccd1 vccd1 _7886_/D sky130_fd_sc_hd__a211oi_1
XANTENNA__7061__A _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1522 _7354_/Q vssd1 vssd1 vccd1 vccd1 _7069_/A sky130_fd_sc_hd__clkbuf_4
X_5138_ _5138_/A1 _4425_/B _5146_/B1 _5137_/X vssd1 vssd1 vccd1 vccd1 _7381_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1544 _7899_/Q vssd1 vssd1 vccd1 vccd1 hold1562/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1511 _7371_/Q vssd1 vssd1 vccd1 vccd1 hold1511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1533 _7692_/Q vssd1 vssd1 vccd1 vccd1 _3729_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 _7083_/X vssd1 vssd1 vccd1 vccd1 _7084_/C sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 _7670_/Q vssd1 vssd1 vccd1 vccd1 _3917_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1566 _5392_/X vssd1 vssd1 vccd1 vccd1 _5402_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1588 _3904_/Y vssd1 vssd1 vccd1 vccd1 _6424_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1599 _4165_/Y vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6160__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5069_ input26/X _5408_/B _5069_/S vssd1 vssd1 vccd1 vccd1 _5070_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4710__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4624__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1761_A _8500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5591__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6215__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5343__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6140__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4777__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7871__CLK _7871_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4082__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcore_473 vssd1 vssd1 vccd1 vccd1 core_473/HI o_pc_IF[0] sky130_fd_sc_hd__conb_1
XFILLER_0_116_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6969__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4440_ _4440_/A _4440_/B vssd1 vssd1 vccd1 vccd1 _4440_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold107 _5676_/X vssd1 vssd1 vccd1 vccd1 _7856_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _6488_/X vssd1 vssd1 vccd1 vccd1 _7970_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _7603_/Q vssd1 vssd1 vccd1 vccd1 _5661_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6110_ _6110_/A1 _6094_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _6110_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__6985__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4371_ _4372_/A _5069_/S vssd1 vssd1 vccd1 vccd1 _4371_/Y sky130_fd_sc_hd__nor2_1
X_7090_ _7090_/A _7090_/B vssd1 vssd1 vccd1 vccd1 _8519_/D sky130_fd_sc_hd__nor2_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6041_ _6144_/S _5853_/C _6342_/S vssd1 vssd1 vccd1 vccd1 _6041_/X sky130_fd_sc_hd__a21o_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4940__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7992_ _8504_/CLK _7992_/D vssd1 vssd1 vccd1 vccd1 _7992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5270__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6943_ _6943_/A _6943_/B vssd1 vssd1 vccd1 vccd1 _6943_/X sky130_fd_sc_hd__and2_1
XANTENNA__4073__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6225__A _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6874_ _7028_/A _6874_/A2 _6906_/A3 _6873_/X vssd1 vssd1 vccd1 vccd1 _6874_/X sky130_fd_sc_hd__a31o_1
X_5825_ _5963_/S _6413_/B1 _6063_/A _5824_/X vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3820__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5756_ _6126_/A _5772_/S vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6879__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6770__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5687_ _6520_/A _5687_/B vssd1 vssd1 vccd1 vccd1 _5687_/X sky130_fd_sc_hd__and2_1
X_8475_ _8475_/CLK _8475_/D vssd1 vssd1 vccd1 vccd1 _8475_/Q sky130_fd_sc_hd__dfxtp_1
X_4707_ _4706_/X _4705_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4638_ _4637_/X _4634_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7516_/D sky130_fd_sc_hd__mux2_1
X_7426_ _8484_/CLK _7426_/D vssd1 vssd1 vccd1 vccd1 _7426_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5325__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 _5279_/X vssd1 vssd1 vccd1 vccd1 _7483_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold652 _5594_/X vssd1 vssd1 vccd1 vccd1 _7778_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 _8299_/Q vssd1 vssd1 vccd1 vccd1 hold663/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 _7487_/Q vssd1 vssd1 vccd1 vccd1 hold641/X sky130_fd_sc_hd__dlygate4sd3_1
X_4569_ _8333_/Q _7809_/Q _7475_/Q _7443_/Q _7362_/Q _7050_/A vssd1 vssd1 vccd1 vccd1
+ _4569_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6895__A _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7357_ _8476_/CLK _7357_/D vssd1 vssd1 vccd1 vccd1 _7357_/Q sky130_fd_sc_hd__dfxtp_4
Xhold696 _5624_/X vssd1 vssd1 vccd1 vccd1 _7804_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 _8219_/Q vssd1 vssd1 vccd1 vccd1 hold685/X sky130_fd_sc_hd__dlygate4sd3_1
X_7288_ _8362_/CLK _7288_/D _7098_/Y vssd1 vssd1 vccd1 vccd1 _7288_/Q sky130_fd_sc_hd__dfrtp_2
X_6308_ _3714_/A _6414_/B1 _6398_/B1 _6295_/A _6292_/A vssd1 vssd1 vccd1 vccd1 _6308_/X
+ sky130_fd_sc_hd__a221o_1
Xhold674 _5210_/X vssd1 vssd1 vccd1 vccd1 _7424_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6239_ _6309_/A _5900_/X _6232_/Y _6238_/X vssd1 vssd1 vccd1 vccd1 _6239_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5023__B _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1330 _8336_/Q vssd1 vssd1 vccd1 vccd1 _6798_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 _7349_/Q vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1341 _6792_/X vssd1 vssd1 vccd1 vccd1 _8333_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4931__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1374 _6782_/X vssd1 vssd1 vccd1 vccd1 _8328_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1363 _6796_/X vssd1 vssd1 vccd1 vccd1 _8335_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1385 _8387_/Q vssd1 vssd1 vccd1 vccd1 _5062_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6589__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1396 _7875_/Q vssd1 vssd1 vccd1 vccd1 hold412/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4695__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5974__A _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6789__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6761__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5316__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7180__58 _8008_/CLK vssd1 vssd1 vccd1 vccd1 _8060_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_31_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4529__S _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4772__B _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3940_ _4745_/B _3966_/B vssd1 vssd1 vccd1 vccd1 _3940_/X sky130_fd_sc_hd__and2_1
XFILLER_0_86_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5252__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3802__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_50_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6201__B1 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3871_ _3871_/A _6209_/A vssd1 vssd1 vccd1 vccd1 _3872_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6752__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6590_ _6967_/A _6559_/B _6591_/B1 hold645/X vssd1 vssd1 vccd1 vccd1 _6590_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_38_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5610_ _6891_/A _5616_/A2 _5616_/B1 _5610_/B2 vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4989__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5541_ _8260_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7730_/D sky130_fd_sc_hd__and3_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_65_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8260_ _8260_/CLK _8260_/D vssd1 vssd1 vccd1 vccd1 _8260_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5307__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5472_ _5472_/A _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7661_/D sky130_fd_sc_hd__and3_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4423_ _4234_/Y _5453_/C _4422_/X _4421_/X vssd1 vssd1 vccd1 vccd1 _8369_/D sky130_fd_sc_hd__a31o_1
X_8191_ _8319_/CLK _8191_/D vssd1 vssd1 vccd1 vccd1 _8191_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3869__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6268__A0 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4354_ _4377_/A _4377_/B _4354_/C vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__and3b_1
X_7240__118 _8218_/CLK vssd1 vssd1 vccd1 vccd1 _8250_/CLK sky130_fd_sc_hd__inv_2
X_7073_ _7073_/A _7073_/B _7073_/C vssd1 vssd1 vccd1 vccd1 _8508_/D sky130_fd_sc_hd__and3_1
Xfanout417 _7063_/A vssd1 vssd1 vccd1 vccd1 _4987_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout406 _4976_/S1 vssd1 vssd1 vccd1 vccd1 _4969_/S1 sky130_fd_sc_hd__buf_4
Xfanout428 _6434_/A vssd1 vssd1 vccd1 vccd1 _7028_/A sky130_fd_sc_hd__buf_4
Xfanout439 _6660_/A1 vssd1 vssd1 vccd1 vccd1 _6551_/A sky130_fd_sc_hd__buf_4
X_6024_ _5946_/A _5974_/A _5993_/A _6016_/A _5772_/S _5804_/A vssd1 vssd1 vccd1 vccd1
+ _6024_/X sky130_fd_sc_hd__mux4_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ _8498_/Q _4285_/B vssd1 vssd1 vccd1 vccd1 _4285_/Y sky130_fd_sc_hd__nand2_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4913__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout275_A _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7975_ _8387_/CLK _7975_/D vssd1 vssd1 vccd1 vccd1 _7975_/Q sky130_fd_sc_hd__dfxtp_1
X_6926_ _7006_/A _6926_/A2 _6943_/B _6925_/X vssd1 vssd1 vccd1 vccd1 _6926_/X sky130_fd_sc_hd__a31o_1
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5497__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5243__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4677__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5794__A2 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout442_A _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6857_ _6923_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6857_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6743__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6788_ _7015_/A _6788_/A2 _6779_/B _6787_/X vssd1 vssd1 vccd1 vccd1 _6788_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5808_ _5709_/X _5712_/X _5838_/A vssd1 vssd1 vccd1 vccd1 _5808_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8527_ _8527_/A _4519_/X vssd1 vssd1 vccd1 vccd1 _8527_/Z sky130_fd_sc_hd__ebufn_1
X_5739_ _6251_/A _6083_/A vssd1 vssd1 vccd1 vccd1 _5739_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_134_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1557_A _8517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8458_ _8458_/CLK _8458_/D vssd1 vssd1 vccd1 vccd1 _8458_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8389_ _8421_/CLK _8389_/D vssd1 vssd1 vccd1 vccd1 _8389_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7409_ _8283_/CLK _7409_/D vssd1 vssd1 vccd1 vccd1 _7409_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold471 _7553_/Q vssd1 vssd1 vccd1 vccd1 hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 _6685_/X vssd1 vssd1 vccd1 vccd1 _8212_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4601__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold493 _7401_/Q vssd1 vssd1 vccd1 vccd1 _5468_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 _5246_/X vssd1 vssd1 vccd1 vccd1 _7454_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1160 _6589_/X vssd1 vssd1 vccd1 vccd1 _8161_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 _6606_/X vssd1 vssd1 vccd1 vccd1 _8167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1193 _8408_/Q vssd1 vssd1 vccd1 vccd1 _6884_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 _8449_/Q vssd1 vssd1 vccd1 vccd1 _6968_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5234__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4037__A2 _3669_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4668__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6409__S1 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__A1 _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6734__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3936__B _7283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4840__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5942__C1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5170__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output71_A _8117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4767__B _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _4070_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _4070_/X sky130_fd_sc_hd__or2_1
XFILLER_0_92_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6422__B1 _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4028__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5776__A2 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4972_ _8354_/Q _7830_/Q _7496_/Q _7464_/Q _7063_/A _4987_/S1 vssd1 vssd1 vccd1 vccd1
+ _4972_/X sky130_fd_sc_hd__mux4_1
X_7760_ _8378_/CLK _7760_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _7282_/Q _3923_/B _7971_/Q vssd1 vssd1 vccd1 vccd1 _3923_/X sky130_fd_sc_hd__and3_1
XFILLER_0_86_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6711_ _6917_/A _6737_/A2 _6737_/B1 _6711_/B2 vssd1 vssd1 vccd1 vccd1 _6711_/X sky130_fd_sc_hd__a22o_1
X_7691_ _8195_/CLK _7691_/D vssd1 vssd1 vccd1 vccd1 _7691_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6642_ _7017_/A _6642_/A2 _6666_/A3 _6641_/X vssd1 vssd1 vccd1 vccd1 _6642_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4722__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3854_ _4766_/B _3966_/B vssd1 vssd1 vccd1 vccd1 _3854_/X sky130_fd_sc_hd__and2_1
XANTENNA__6725__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6573_ _6933_/A _6592_/A2 _6592_/B1 hold937/X vssd1 vssd1 vccd1 vccd1 _6573_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5119__A _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3785_ _6175_/A _6172_/A vssd1 vssd1 vccd1 vccd1 _3787_/A sky130_fd_sc_hd__nand2_1
X_8312_ _8476_/CLK _8312_/D vssd1 vssd1 vccd1 vccd1 _8312_/Q sky130_fd_sc_hd__dfxtp_1
X_5524_ _8243_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7713_/D sky130_fd_sc_hd__and3_1
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8243_ _8243_/CLK _8243_/D vssd1 vssd1 vccd1 vccd1 _8243_/Q sky130_fd_sc_hd__dfxtp_1
X_5455_ _5455_/A _5503_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _5455_/X sky130_fd_sc_hd__and3_1
X_8174_ _8517_/CLK _8174_/D vssd1 vssd1 vccd1 vccd1 _8174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4406_ _4410_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__or2_1
X_5386_ _5385_/Y _5386_/B vssd1 vssd1 vccd1 vccd1 _6983_/B sky130_fd_sc_hd__nand2b_1
Xfanout203 _3907_/Y vssd1 vssd1 vccd1 vccd1 _6270_/A sky130_fd_sc_hd__buf_4
Xfanout214 _5456_/C vssd1 vssd1 vccd1 vccd1 _5454_/C sky130_fd_sc_hd__buf_4
Xfanout225 _5449_/C vssd1 vssd1 vccd1 vccd1 _7082_/B sky130_fd_sc_hd__buf_4
XANTENNA_fanout392_A _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 _5182_/A2 vssd1 vssd1 vccd1 vccd1 _5069_/S sky130_fd_sc_hd__buf_4
X_4337_ _4335_/Y _4337_/B vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__nand2b_1
Xfanout247 _6705_/Y vssd1 vssd1 vccd1 vccd1 _6737_/B1 sky130_fd_sc_hd__buf_8
XFILLER_0_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout258 _5335_/Y vssd1 vssd1 vccd1 vccd1 _5368_/B1 sky130_fd_sc_hd__clkbuf_8
X_7056_ hold90/X _7071_/B _7064_/B1 vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__a21oi_1
Xfanout269 _4084_/B2 vssd1 vssd1 vccd1 vccd1 _4073_/B2 sky130_fd_sc_hd__buf_6
XFILLER_0_66_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4268_ _5567_/B _5036_/A1 _5465_/B vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4898__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6007_ _6270_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6362_/C sky130_fd_sc_hd__nor2_2
XFILLER_0_97_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4199_ _5557_/B _4434_/A _7073_/A vssd1 vssd1 vccd1 vccd1 _4200_/B sky130_fd_sc_hd__mux2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6413__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5216__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6964__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7958_ _8504_/CLK _7958_/D vssd1 vssd1 vccd1 vccd1 _7958_/Q sky130_fd_sc_hd__dfxtp_1
X_6909_ _6909_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6909_/X sky130_fd_sc_hd__and2_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7889_ _8086_/CLK _7889_/D vssd1 vssd1 vccd1 vccd1 _7889_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3860__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6716__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4822__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5971__B _5971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3772__A _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5152__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7150__28 _8160_/CLK vssd1 vssd1 vccd1 vccd1 _7527_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_32_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold290 _7567_/Q vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4889__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__A1 _4761_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3769__B2 _3767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6707__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6183__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5240_ _6933_/A _5226_/B _5259_/B1 hold595/X vssd1 vssd1 vccd1 vccd1 _5240_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5171_ hold65/X _5463_/C vssd1 vssd1 vccd1 vccd1 _5171_/X sky130_fd_sc_hd__or2_1
X_4122_ _6191_/A _6188_/A vssd1 vssd1 vccd1 vccd1 _4122_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4053_ _8505_/Q _4052_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _6094_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 i_instr_ID[12] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_1
XFILLER_0_127_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5997__A2 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6217__B _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7812_ _8332_/CLK _7812_/D vssd1 vssd1 vccd1 vccd1 _7812_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5749__A2 _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6946__A1 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7743_ _8361_/CLK _7743_/D vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
X_4955_ _8481_/Q _8413_/Q _8445_/Q _8319_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4955_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_59_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3906_ _3968_/A _3904_/Y _3905_/Y vssd1 vssd1 vccd1 vccd1 _3906_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3857__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7674_ _8343_/CLK _7674_/D vssd1 vssd1 vccd1 vccd1 _7674_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout238_A _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4886_ _4885_/X _4884_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4886_/X sky130_fd_sc_hd__mux2_1
X_3837_ _8098_/Q _7970_/Q _8034_/Q _8002_/Q _7282_/Q _3923_/B vssd1 vssd1 vccd1 vccd1
+ _3837_/X sky130_fd_sc_hd__mux4_2
XANTENNA__7048__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6625_ _6931_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6625_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6556_ _7937_/Q _7938_/Q _5183_/X vssd1 vssd1 vccd1 vccd1 _6776_/B sky130_fd_sc_hd__or3b_4
X_3768_ _3768_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _3768_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout405_A _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4804__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7246__124 _8442_/CLK vssd1 vssd1 vccd1 vccd1 _8256_/CLK sky130_fd_sc_hd__inv_2
X_5507_ _7528_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7696_/D sky130_fd_sc_hd__and3_1
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6887__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3699_ _3652_/Y _7937_/Q _5222_/B _7661_/Q _3697_/X vssd1 vssd1 vccd1 vccd1 _3705_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5134__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8226_ _8319_/CLK _8226_/D vssd1 vssd1 vccd1 vccd1 _8226_/Q sky130_fd_sc_hd__dfxtp_1
X_6487_ _6520_/A _6487_/B vssd1 vssd1 vccd1 vccd1 _6487_/X sky130_fd_sc_hd__and2_1
XFILLER_0_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5438_ _5438_/A _5470_/B _5470_/C vssd1 vssd1 vccd1 vccd1 _5438_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5369_ _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _7079_/B sky130_fd_sc_hd__and2_2
X_8157_ _8355_/CLK _8157_/D vssd1 vssd1 vccd1 vccd1 _8157_/Q sky130_fd_sc_hd__dfxtp_1
X_8088_ _8451_/CLK _8122_/D vssd1 vssd1 vccd1 vccd1 _8088_/Q sky130_fd_sc_hd__dfxtp_1
X_7108_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7108_/Y sky130_fd_sc_hd__inv_2
X_7039_ _7031_/Y _7039_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _7039_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4627__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3999__B2 _8013_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_116_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8440_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6165__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6797__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output157_A _8043_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6318__A _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6640__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6928__A1 _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3677__A _7282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3837__S1 _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _8197_/Q _8229_/Q _8293_/Q _7801_/Q _4741_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4740_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_107_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8350_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4671_ _8477_/Q _8409_/Q _8441_/Q _8315_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4671_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5892__A _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6410_ _6340_/X _6409_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6410_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7390_ _8504_/CLK _7390_/D vssd1 vssd1 vccd1 vccd1 _7390_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5364__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6341_ _6268_/X _6340_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5116__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6313__C1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6272_ _3883_/A _6414_/B1 _6398_/B1 _6259_/A _6292_/A vssd1 vssd1 vccd1 vccd1 _6272_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8011_ _8011_/CLK _8011_/D vssd1 vssd1 vccd1 vccd1 _8011_/Q sky130_fd_sc_hd__dfxtp_1
X_5223_ _5581_/A _7940_/Q vssd1 vssd1 vccd1 vccd1 _6776_/A sky130_fd_sc_hd__nand2_4
XANTENNA__4020__B _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5154_ _5154_/A1 _4407_/B _5166_/B1 _5153_/X vssd1 vssd1 vccd1 vccd1 _7389_/D sky130_fd_sc_hd__o211a_1
X_4105_ _4099_/Y _4104_/X _4045_/X vssd1 vssd1 vccd1 vccd1 _4105_/X sky130_fd_sc_hd__a21o_1
Xhold1726 _3736_/Y vssd1 vssd1 vccd1 vccd1 _6294_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_4_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1704 _7653_/Q vssd1 vssd1 vccd1 vccd1 _4314_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1715 _7648_/Q vssd1 vssd1 vccd1 vccd1 _4278_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5085_ _6977_/B _5085_/B vssd1 vssd1 vccd1 vccd1 _5085_/Y sky130_fd_sc_hd__nand2_1
Xhold1737 _5742_/X vssd1 vssd1 vccd1 vccd1 _5743_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1748 _8488_/Q vssd1 vssd1 vccd1 vccd1 _3840_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1759 _6318_/A vssd1 vssd1 vccd1 vccd1 _3723_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4036_ _7709_/Q _4081_/B vssd1 vssd1 vccd1 vccd1 _4036_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_635 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7041__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3850__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5987_ _5976_/X _5977_/Y _5986_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _5987_/X sky130_fd_sc_hd__a22o_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7059__A _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4938_ _8156_/Q _7555_/Q _7427_/Q _7587_/Q _4990_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4938_/X sky130_fd_sc_hd__mux4_1
X_7726_ _8355_/CLK _7726_/D vssd1 vssd1 vccd1 vccd1 _7726_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4869_ _4867_/X _4868_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7657_ _8501_/CLK _7657_/D vssd1 vssd1 vccd1 vccd1 _7657_/Q sky130_fd_sc_hd__dfxtp_1
X_6608_ _6847_/A _6605_/B _6607_/X vssd1 vssd1 vccd1 vccd1 _6608_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5355__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7588_ _8160_/CLK _7588_/D vssd1 vssd1 vccd1 vccd1 _7588_/Q sky130_fd_sc_hd__dfxtp_1
X_6539_ _6539_/A _6539_/B vssd1 vssd1 vccd1 vccd1 _8021_/D sky130_fd_sc_hd__and2_1
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8209_ _8431_/CLK _8209_/D vssd1 vssd1 vccd1 vccd1 _8209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6870__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7879__D _7879_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6138__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6622__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5830__A1 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5594__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4820__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5346__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5649__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3960__A _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4775__B _4775_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4085__A0 _4085_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5910_ _5908_/X _5909_/X _6302_/A vssd1 vssd1 vccd1 vccd1 _5911_/A sky130_fd_sc_hd__mux2_1
X_6890_ _7024_/A _6890_/A2 _6906_/A3 _6889_/X vssd1 vssd1 vccd1 vccd1 _6890_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_124_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5841_ _5832_/X _5840_/Y _6270_/A vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5772_ _4094_/B _3949_/Y _5772_/S vssd1 vssd1 vccd1 vccd1 _5773_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_29_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8491_ _8494_/CLK _8491_/D vssd1 vssd1 vccd1 vccd1 _8491_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7511_ _7511_/CLK _7511_/D vssd1 vssd1 vccd1 vccd1 _7511_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4723_ _8355_/Q _7831_/Q _7497_/Q _7465_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4723_/X sky130_fd_sc_hd__mux4_1
X_7186__64 _8480_/CLK vssd1 vssd1 vccd1 vccd1 _8066_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_8_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7442_ _8426_/CLK _7442_/D vssd1 vssd1 vccd1 vccd1 _7442_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4654_ _8152_/Q _7551_/Q _7423_/Q _7583_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4654_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6511__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput61 i_read_data_M[8] vssd1 vssd1 vccd1 vccd1 _6529_/B sky130_fd_sc_hd__clkbuf_1
X_7373_ _7907_/CLK _7373_/D vssd1 vssd1 vccd1 vccd1 _7373_/Q sky130_fd_sc_hd__dfxtp_1
Xhold801 _7442_/Q vssd1 vssd1 vccd1 vccd1 hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput50 i_read_data_M[27] vssd1 vssd1 vccd1 vccd1 _6548_/B sky130_fd_sc_hd__clkbuf_1
X_4585_ _4583_/X _4584_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4585_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3899__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold812 _5285_/X vssd1 vssd1 vccd1 vccd1 _7489_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3854__B _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4031__A _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 _8307_/Q vssd1 vssd1 vccd1 vccd1 hold845/X sky130_fd_sc_hd__dlygate4sd3_1
X_6324_ _6179_/X _6323_/X _6411_/S vssd1 vssd1 vccd1 vccd1 _6324_/X sky130_fd_sc_hd__mux2_1
Xhold823 _7479_/Q vssd1 vssd1 vccd1 vccd1 hold823/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold834 _5208_/X vssd1 vssd1 vccd1 vccd1 _7422_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 _6688_/X vssd1 vssd1 vccd1 vccd1 _8215_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold878 _7011_/X vssd1 vssd1 vccd1 vccd1 _8469_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 _7821_/Q vssd1 vssd1 vccd1 vccd1 hold889/X sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ _3896_/A _6414_/A2 _5927_/X _6412_/S _6254_/X vssd1 vssd1 vccd1 vccd1 _6255_/X
+ sky130_fd_sc_hd__a221o_1
Xhold867 _8209_/Q vssd1 vssd1 vccd1 vccd1 hold867/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5206_ _6941_/A _5221_/A2 _5220_/B1 hold447/X vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6186_ _6391_/A _6177_/Y _6181_/Y _6309_/A _6185_/X vssd1 vssd1 vccd1 vccd1 _6186_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__6852__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1501 _7891_/Q vssd1 vssd1 vccd1 vccd1 hold1501/X sky130_fd_sc_hd__dlygate4sd3_1
X_5137_ _5448_/A _5453_/C vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__or2_1
Xhold1523 _7069_/Y vssd1 vssd1 vccd1 vccd1 _7070_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1512 _7082_/A vssd1 vssd1 vccd1 vccd1 hold1512/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4177__S _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7061__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1534 _3729_/X vssd1 vssd1 vccd1 vccd1 _3730_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6604__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1567 _7089_/X vssd1 vssd1 vccd1 vccd1 _7090_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1556 _3917_/Y vssd1 vssd1 vccd1 vccd1 _6423_/B sky130_fd_sc_hd__buf_1
X_5068_ _7273_/A _5068_/B _5465_/B vssd1 vssd1 vccd1 vccd1 _7346_/D sky130_fd_sc_hd__or3b_1
Xhold1545 _3830_/Y vssd1 vssd1 vccd1 vccd1 _6450_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1578 _7084_/X vssd1 vssd1 vccd1 vccd1 _8516_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4019_ _4020_/A _5974_/A vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__or2_1
XANTENNA__6160__S1 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1589 _7655_/Q vssd1 vssd1 vccd1 vccd1 _4329_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6405__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7709_ _8143_/CLK _7709_/D vssd1 vssd1 vccd1 vccd1 _7709_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5040__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6421__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5328__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7252__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6315__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xcore_474 vssd1 vssd1 vccd1 vccd1 core_474/HI o_pc_IF[1] sky130_fd_sc_hd__conb_1
XFILLER_0_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5319__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4550__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 _7758_/Q vssd1 vssd1 vccd1 vccd1 _6509_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _6419_/B _4370_/B _6418_/B vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__or3b_1
Xhold119 _5661_/X vssd1 vssd1 vccd1 vccd1 _7841_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5098__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6040_ _5961_/X _6039_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6040_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6834__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7991_ _8020_/CLK _7991_/D vssd1 vssd1 vccd1 vccd1 _7991_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6942_ _7017_/A _6942_/A2 _6970_/A3 _6941_/X vssd1 vssd1 vccd1 vccd1 _6942_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3805__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6506__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4725__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5270__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6873_ _6939_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6873_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5824_ _5820_/A _5963_/S _6398_/A2 vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5022__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5755_ _6411_/S _5754_/Y _5748_/Y vssd1 vssd1 vccd1 vccd1 _5755_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__3865__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6770__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5686_ _6539_/A _5686_/B vssd1 vssd1 vccd1 vccd1 _5686_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout220_A _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8474_ _8476_/CLK _8474_/D vssd1 vssd1 vccd1 vccd1 _8474_/Q sky130_fd_sc_hd__dfxtp_1
X_4706_ _8482_/Q _8414_/Q _8446_/Q _8320_/Q _4706_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4706_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7425_ _8283_/CLK _7425_/D vssd1 vssd1 vccd1 vccd1 _7425_/Q sky130_fd_sc_hd__dfxtp_1
X_4637_ _4636_/X _4635_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold620 _6753_/X vssd1 vssd1 vccd1 vccd1 _8304_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7356_ _8011_/CLK _7356_/D vssd1 vssd1 vccd1 vccd1 _7356_/Q sky130_fd_sc_hd__dfxtp_1
X_4568_ _4567_/X _4564_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7506_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_69_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold642 _5283_/X vssd1 vssd1 vccd1 vccd1 _7487_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _8220_/Q vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6895__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold653 _8291_/Q vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _8462_/Q vssd1 vssd1 vccd1 vccd1 _7004_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 _6748_/X vssd1 vssd1 vccd1 vccd1 _8299_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _6692_/X vssd1 vssd1 vccd1 vccd1 _8219_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7287_ _8361_/CLK _7287_/D _7097_/Y vssd1 vssd1 vccd1 vccd1 _7287_/Q sky130_fd_sc_hd__dfrtp_4
X_6307_ _6307_/A _6307_/B vssd1 vssd1 vccd1 vccd1 _6307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4499_ _5154_/A1 _4262_/C _5454_/C vssd1 vssd1 vccd1 vccd1 _7299_/D sky130_fd_sc_hd__mux2_1
Xhold675 _8309_/Q vssd1 vssd1 vccd1 vccd1 hold675/X sky130_fd_sc_hd__dlygate4sd3_1
X_6238_ _6391_/A _6229_/X _6236_/X _6237_/X vssd1 vssd1 vccd1 vccd1 _6238_/X sky130_fd_sc_hd__o22a_1
X_6169_ _6157_/A _6154_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6169_/X sky130_fd_sc_hd__a21bo_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1331 _6798_/X vssd1 vssd1 vccd1 vccd1 _8336_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 _8170_/Q vssd1 vssd1 vccd1 vccd1 _6612_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1342 _8344_/Q vssd1 vssd1 vccd1 vccd1 _6814_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_96_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _8195_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1386 _7350_/Q vssd1 vssd1 vccd1 vccd1 _5544_/A sky130_fd_sc_hd__clkbuf_2
Xhold1353 _5073_/A vssd1 vssd1 vccd1 vccd1 _5543_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1375 _7355_/Q vssd1 vssd1 vccd1 vccd1 _7067_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__6589__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1364 _8377_/Q vssd1 vssd1 vccd1 vccd1 _5042_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1397 _6456_/X vssd1 vssd1 vccd1 vccd1 _7938_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4695__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3775__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6761__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8413_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6816__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_87_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _8032_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5252__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4122__A_N _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6201__A1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3870_ _3871_/A _6209_/A vssd1 vssd1 vccd1 vccd1 _3872_/A sky130_fd_sc_hd__or2_1
XANTENNA__6752__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _8354_/CLK sky130_fd_sc_hd__clkbuf_16
X_7156__34 _8431_/CLK vssd1 vssd1 vccd1 vccd1 _8036_/CLK sky130_fd_sc_hd__inv_2
X_5540_ _8259_/Q _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _7729_/D sky130_fd_sc_hd__and3_1
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5471_ _7052_/A _7090_/A vssd1 vssd1 vccd1 vccd1 _7660_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_41_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ _4422_/A _4422_/B vssd1 vssd1 vccd1 vccd1 _4422_/X sky130_fd_sc_hd__or2_1
XANTENNA__5712__A0 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8190_ _8480_/CLK _8190_/D vssd1 vssd1 vccd1 vccd1 _8190_/Q sky130_fd_sc_hd__dfxtp_1
X_4353_ _5579_/B _5060_/A1 _5470_/B vssd1 vssd1 vccd1 vccd1 _4354_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_10_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7072_ _3651_/A _7071_/A _7055_/A _7072_/B2 _7071_/Y vssd1 vssd1 vccd1 vccd1 _7073_/C
+ sky130_fd_sc_hd__a221o_1
X_8528__476 vssd1 vssd1 vccd1 vccd1 _8528_/A _8528__476/LO sky130_fd_sc_hd__conb_1
XANTENNA__6268__A1 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 _4976_/S1 vssd1 vssd1 vccd1 vccd1 _4987_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout418 _7063_/A vssd1 vssd1 vccd1 vccd1 _4983_/S0 sky130_fd_sc_hd__buf_8
Xfanout429 _7025_/A vssd1 vssd1 vccd1 vccd1 _7024_/A sky130_fd_sc_hd__buf_4
X_4284_ _8498_/Q _4285_/B vssd1 vssd1 vccd1 vccd1 _4284_/Y sky130_fd_sc_hd__nor2_1
X_6023_ _6063_/A _6023_/B _6023_/C vssd1 vssd1 vccd1 vccd1 _6023_/Y sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_78_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _8360_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5779__A0 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7974_ _8361_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 _7974_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout170_A _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6925_ _6925_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6925_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5243__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4677__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5794__A3 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6856_ _7008_/A _6856_/A2 _6845_/B _6855_/X vssd1 vssd1 vccd1 vccd1 _6856_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3999_ _7981_/Q _4079_/A2 _4079_/B1 _8013_/Q _3998_/X vssd1 vssd1 vccd1 vccd1 _3999_/X
+ sky130_fd_sc_hd__a221o_1
X_6787_ _6787_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6787_/X sky130_fd_sc_hd__and2_1
X_5807_ _5706_/X _5708_/X _5838_/A vssd1 vssd1 vccd1 vccd1 _5807_/X sky130_fd_sc_hd__mux2_1
X_5738_ _5738_/A _5738_/B vssd1 vssd1 vccd1 vccd1 _6083_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_115_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8457_ _8457_/CLK _8457_/D vssd1 vssd1 vccd1 vccd1 _8457_/Q sky130_fd_sc_hd__dfxtp_1
X_5669_ _6548_/A _5669_/B vssd1 vssd1 vccd1 vccd1 _5669_/X sky130_fd_sc_hd__and2_1
XANTENNA_hold1452_A _7284_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8388_ _8388_/CLK _8388_/D vssd1 vssd1 vccd1 vccd1 _8388_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7408_ _8355_/CLK _7408_/D vssd1 vssd1 vccd1 vccd1 _7408_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold472 _5322_/X vssd1 vssd1 vccd1 vccd1 _7553_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7339_ _8030_/CLK _7339_/D vssd1 vssd1 vccd1 vccd1 _7339_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4601__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold461 _8222_/Q vssd1 vssd1 vccd1 vccd1 hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _5252_/X vssd1 vssd1 vccd1 vccd1 _7460_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _8296_/Q vssd1 vssd1 vccd1 vccd1 hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _5468_/X vssd1 vssd1 vccd1 vccd1 _7657_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _8363_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1150 _6962_/X vssd1 vssd1 vccd1 vccd1 _8446_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 _8397_/Q vssd1 vssd1 vccd1 vccd1 _6862_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1161 _8348_/Q vssd1 vssd1 vccd1 vccd1 _6822_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1194 _6884_/X vssd1 vssd1 vccd1 vccd1 _8408_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1172 _6968_/X vssd1 vssd1 vccd1 vccd1 _8449_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5234__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4668__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6195__A0 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6734__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4840__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5924__S _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output64_A _8101_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8471_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_116_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6056__A _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5856__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4971_ _4970_/X _4967_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8257_/D sky130_fd_sc_hd__mux2_1
X_6710_ _6849_/A _6705_/B _6738_/B1 hold715/X vssd1 vssd1 vccd1 vccd1 _6710_/X sky130_fd_sc_hd__a22o_1
X_3922_ _4097_/A _3922_/B vssd1 vssd1 vccd1 vccd1 _3922_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7690_ _8427_/CLK _7690_/D vssd1 vssd1 vccd1 vccd1 _7690_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6641_ _6947_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6641_/X sky130_fd_sc_hd__and2_1
X_3853_ _4766_/B _4071_/A2 _4071_/B1 _6953_/A _3852_/X vssd1 vssd1 vccd1 vccd1 _6244_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6725__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5119__B _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8311_ _8473_/CLK _8311_/D vssd1 vssd1 vccd1 vccd1 _8311_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6572_ _6931_/A _6559_/B _6591_/B1 hold851/X vssd1 vssd1 vccd1 vccd1 _6572_/X sky130_fd_sc_hd__a22o_1
X_3784_ _4263_/A _3783_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6172_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_6_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5523_ _8242_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7712_/D sky130_fd_sc_hd__and3_1
X_8242_ _8242_/CLK _8242_/D vssd1 vssd1 vccd1 vccd1 _8242_/Q sky130_fd_sc_hd__dfxtp_1
X_5454_ _5454_/A _5503_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _5454_/X sky130_fd_sc_hd__and3_1
XFILLER_0_112_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5385_ _7067_/A _7069_/A vssd1 vssd1 vccd1 vccd1 _5385_/Y sky130_fd_sc_hd__xnor2_1
X_8173_ _8173_/CLK _8173_/D vssd1 vssd1 vccd1 vccd1 _8173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4405_ _4276_/Y _5456_/C _4404_/X _4403_/X vssd1 vssd1 vccd1 vccd1 _8375_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_100_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout204 _6411_/S vssd1 vssd1 vccd1 vccd1 _6008_/A sky130_fd_sc_hd__buf_4
X_4336_ _8491_/Q _4336_/B vssd1 vssd1 vccd1 vccd1 _4336_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout226 _5449_/C vssd1 vssd1 vccd1 vccd1 _5442_/C sky130_fd_sc_hd__clkbuf_4
Xfanout237 _5099_/B vssd1 vssd1 vccd1 vccd1 _5182_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout215 _5456_/C vssd1 vssd1 vccd1 vccd1 _5462_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout385_A _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout248 _6705_/Y vssd1 vssd1 vccd1 vccd1 _6738_/B1 sky130_fd_sc_hd__buf_6
X_7055_ _7055_/A _7055_/B _7031_/A vssd1 vssd1 vccd1 vccd1 _7071_/B sky130_fd_sc_hd__or3b_4
Xfanout259 _5299_/Y vssd1 vssd1 vccd1 vccd1 _5331_/B1 sky130_fd_sc_hd__buf_6
X_4267_ _4267_/A _4267_/B vssd1 vssd1 vccd1 vccd1 _4267_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_5_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4898__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4198_ _4198_/A _4198_/B vssd1 vssd1 vccd1 vccd1 _4198_/X sky130_fd_sc_hd__xor2_1
X_6006_ _6008_/A _5754_/Y _5955_/Y vssd1 vssd1 vccd1 vccd1 _6307_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_96_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6413__A1 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5216__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7957_ _8071_/CLK _7957_/D vssd1 vssd1 vccd1 vccd1 _7957_/Q sky130_fd_sc_hd__dfxtp_1
X_6908_ _7939_/Q _7940_/Q _6908_/C vssd1 vssd1 vccd1 vccd1 _6908_/X sky130_fd_sc_hd__or3_4
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7888_ _8463_/CLK _7888_/D vssd1 vssd1 vccd1 vccd1 _7888_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3778__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6839_ _6971_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6839_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6716__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4822__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8509_ _8510_/CLK _8509_/D vssd1 vssd1 vccd1 vccd1 _8509_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5744__S _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6024__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4586__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold280 _8136_/Q vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 _5340_/X vssd1 vssd1 vccd1 vccd1 _7567_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7260__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4889__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_64_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4823__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3769__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output102_A _7297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3947__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6707__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_79_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6977__C _7354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6340__A0 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4577__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5170_ _5170_/A1 _5067_/S _5172_/B1 _5169_/X vssd1 vssd1 vccd1 vccd1 _7397_/D sky130_fd_sc_hd__o211a_1
X_4121_ _3848_/A _4120_/X _4119_/Y vssd1 vssd1 vccd1 vccd1 _4121_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_127_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4052_ _4052_/A1 _4084_/A2 _6937_/A _4084_/B2 _4051_/X vssd1 vssd1 vccd1 vccd1 _4052_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_127_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5997__A3 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput4 i_instr_ID[13] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_2
XFILLER_0_127_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7811_ _8461_/CLK _7811_/D vssd1 vssd1 vccd1 vccd1 _7811_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5749__A3 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4954_ _8191_/Q _8223_/Q _8287_/Q _7795_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4954_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_59_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7742_ _8387_/CLK _7742_/D vssd1 vssd1 vccd1 vccd1 _7742_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6514__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3905_ _3968_/A _8516_/Q vssd1 vssd1 vccd1 vccd1 _3905_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7673_ _8473_/CLK _7673_/D vssd1 vssd1 vccd1 vccd1 _7673_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4885_ _8471_/Q _8403_/Q _8435_/Q _8309_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4885_/X sky130_fd_sc_hd__mux4_1
X_6624_ _7008_/A _6624_/A2 _6605_/B _6623_/X vssd1 vssd1 vccd1 vccd1 _6624_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _3836_/A _3836_/B vssd1 vssd1 vccd1 vccd1 _3848_/C sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3767_ _8084_/Q _3766_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _3767_/X sky130_fd_sc_hd__mux2_2
X_6555_ _5409_/A _6554_/X _7090_/A vssd1 vssd1 vccd1 vccd1 _8100_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4804__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5506_ _7527_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7695_/D sky130_fd_sc_hd__and3_1
X_3698_ _7661_/Q _5222_/B _5581_/A _7662_/Q vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__a2bb2o_1
X_6486_ _6524_/A hold25/X vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__and2_1
X_8225_ _8483_/CLK _8225_/D vssd1 vssd1 vccd1 vccd1 _8225_/Q sky130_fd_sc_hd__dfxtp_1
X_5437_ _5437_/A _5470_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _5437_/X sky130_fd_sc_hd__and3_1
X_5368_ _6971_/A _5335_/B _5368_/B1 hold711/X vssd1 vssd1 vccd1 vccd1 _5368_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6882__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8156_ _8486_/CLK _8156_/D vssd1 vssd1 vccd1 vccd1 _8156_/Q sky130_fd_sc_hd__dfxtp_1
X_5299_ _6741_/A _5299_/B vssd1 vssd1 vccd1 vccd1 _5299_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4908__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8087_ _8479_/CLK _8121_/D vssd1 vssd1 vccd1 vccd1 _8087_/Q sky130_fd_sc_hd__dfxtp_1
X_7107_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7107_/Y sky130_fd_sc_hd__inv_2
X_4319_ _4318_/Y _5050_/A1 _5465_/B vssd1 vssd1 vccd1 vccd1 _4327_/C sky130_fd_sc_hd__mux2_1
X_7038_ _7077_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7038_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6634__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3999__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4740__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6398__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7210__88 _8501_/CLK vssd1 vssd1 vccd1 vccd1 _8123_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6570__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7255__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6322__A0 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4559__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6086__C1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3722__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4731__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6334__A _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4553__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3677__B _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5600__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6053__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4670_ _8187_/Q _8219_/Q _8283_/Q _7791_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4670_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_71_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4798__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6561__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5364__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8531__472 vssd1 vssd1 vccd1 vccd1 _8531__472/HI _8531_/A sky130_fd_sc_hd__conb_1
X_6340_ _6298_/A _6281_/A _6334_/A _6318_/A _5744_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6340_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6271_ _6411_/S _6122_/X _6270_/X _5740_/B vssd1 vssd1 vccd1 vccd1 _6271_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6864__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5222_ _5296_/A _5222_/B _5183_/X vssd1 vssd1 vccd1 vccd1 _6740_/C sky130_fd_sc_hd__or3b_4
X_8010_ _8010_/CLK _8010_/D vssd1 vssd1 vccd1 vccd1 _8010_/Q sky130_fd_sc_hd__dfxtp_4
X_5153_ _5456_/A _5540_/C vssd1 vssd1 vccd1 vccd1 _5153_/X sky130_fd_sc_hd__or2_1
XANTENNA__4728__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6616__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4104_ _4092_/B _4098_/X _4103_/X _3985_/X vssd1 vssd1 vccd1 vccd1 _4104_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6509__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1705 _4314_/Y vssd1 vssd1 vccd1 vccd1 _4315_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1716 _4278_/Y vssd1 vssd1 vccd1 vccd1 _4279_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5084_ input3/X _5144_/A2 _5146_/B1 _5083_/X vssd1 vssd1 vccd1 vccd1 _7354_/D sky130_fd_sc_hd__o211a_1
Xhold1727 _8507_/Q vssd1 vssd1 vccd1 vccd1 _4221_/A sky130_fd_sc_hd__clkbuf_2
Xhold1738 _5743_/Y vssd1 vssd1 vccd1 vccd1 _7868_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1749 _3846_/A vssd1 vssd1 vccd1 vccd1 _6417_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4035_ _8076_/Q _4034_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4035_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_79_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout250_A _6669_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6244__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5986_ _5694_/Y _5985_/X _5984_/Y vssd1 vssd1 vccd1 vccd1 _5986_/X sky130_fd_sc_hd__a21bo_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5052__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7725_ _8086_/CLK _7725_/D vssd1 vssd1 vccd1 vccd1 _7725_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7059__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4937_ _8349_/Q _7825_/Q _7491_/Q _7459_/Q _4990_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4937_/X sky130_fd_sc_hd__mux4_1
X_4868_ _8146_/Q _7545_/Q _7417_/Q _7577_/Q _4997_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4868_/X sky130_fd_sc_hd__mux4_1
XANTENNA_20 _7289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7656_ _8494_/CLK hold68/X vssd1 vssd1 vccd1 vccd1 _7656_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6607_ _6911_/A _6607_/B _6661_/B vssd1 vssd1 vccd1 vccd1 _6607_/X sky130_fd_sc_hd__or3_1
X_3819_ _3819_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3819_/X sky130_fd_sc_hd__or2_1
XANTENNA__5355__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4799_ _4797_/X _4798_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__7075__A _7075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7587_ _8486_/CLK _7587_/D vssd1 vssd1 vccd1 vccd1 _7587_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6538_ _6550_/A _6538_/B vssd1 vssd1 vccd1 vccd1 _8020_/D sky130_fd_sc_hd__and2_1
X_6469_ _6552_/A hold69/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__and2_1
XFILLER_0_113_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8208_ _8462_/CLK _8208_/D vssd1 vssd1 vccd1 vccd1 _8208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8139_ _8175_/CLK _8139_/D vssd1 vssd1 vccd1 vccd1 _8139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4638__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6419__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4961__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4713__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5830__A2 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5291__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6240__C1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5594__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5993__A _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5346__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3717__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3873__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6846__A1 _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5649__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4952__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4085__A1 _4084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5282__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3832__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5840_ _5840_/A vssd1 vssd1 vccd1 vccd1 _5840_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6231__C1 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5034__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6999__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5771_ _6105_/A2 _5769_/A _5770_/X vssd1 vssd1 vccd1 vccd1 _5771_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7510_ _7510_/CLK _7510_/D vssd1 vssd1 vccd1 vccd1 _7510_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4722_ _4721_/X _4718_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7528_/D sky130_fd_sc_hd__mux2_1
X_8490_ _8501_/CLK _8490_/D vssd1 vssd1 vccd1 vccd1 _8490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5337__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7441_ _8461_/CLK _7441_/D vssd1 vssd1 vccd1 vccd1 _7441_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput40 i_read_data_M[18] vssd1 vssd1 vccd1 vccd1 _6539_/B sky130_fd_sc_hd__clkbuf_1
X_4653_ _8345_/Q _7821_/Q _7487_/Q _7455_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4653_/X sky130_fd_sc_hd__mux4_1
Xhold802 _5234_/X vssd1 vssd1 vccd1 vccd1 _7442_/D sky130_fd_sc_hd__dlygate4sd3_1
Xinput51 i_read_data_M[28] vssd1 vssd1 vccd1 vccd1 _6549_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4584_ _8142_/Q _7541_/Q _7413_/Q _7573_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4584_/X sky130_fd_sc_hd__mux4_1
X_7372_ _8507_/CLK _7372_/D vssd1 vssd1 vccd1 vccd1 _7372_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput62 i_read_data_M[9] vssd1 vssd1 vccd1 vccd1 _6530_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold835 _7815_/Q vssd1 vssd1 vccd1 vccd1 hold835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold846 _6756_/X vssd1 vssd1 vccd1 vccd1 _8307_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5127__B _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6323_ _6248_/X _6393_/B _6410_/S vssd1 vssd1 vccd1 vccd1 _6323_/X sky130_fd_sc_hd__mux2_1
Xhold824 _5275_/X vssd1 vssd1 vccd1 vccd1 _7479_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold813 _7591_/Q vssd1 vssd1 vccd1 vccd1 hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _7414_/Q vssd1 vssd1 vccd1 vccd1 hold857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 _7795_/Q vssd1 vssd1 vccd1 vccd1 hold879/X sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ _3859_/A _6414_/B1 _6398_/B1 _6242_/A _6292_/A vssd1 vssd1 vccd1 vccd1 _6254_/X
+ sky130_fd_sc_hd__a221o_1
Xhold868 _6682_/X vssd1 vssd1 vccd1 vccd1 _8209_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3870__B _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5205_ _6939_/A _5188_/B _5220_/B1 hold505/X vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout298_A _6557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6185_ _5815_/X _6128_/B _6184_/X vssd1 vssd1 vccd1 vccd1 _6185_/X sky130_fd_sc_hd__o21ba_1
Xhold1513 hold1805/X vssd1 vssd1 vccd1 vccd1 _5546_/A sky130_fd_sc_hd__buf_1
Xhold1502 _6458_/X vssd1 vssd1 vccd1 vccd1 _7940_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1524 _7070_/Y vssd1 vssd1 vccd1 vccd1 _8507_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5136_ _5136_/A1 _5085_/B _5140_/B1 _5135_/X vssd1 vssd1 vccd1 vccd1 _7380_/D sky130_fd_sc_hd__o211a_1
Xhold1535 _7635_/Q vssd1 vssd1 vccd1 vccd1 _4187_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1557 _8517_/Q vssd1 vssd1 vccd1 vccd1 _4161_/A sky130_fd_sc_hd__clkbuf_2
Xhold1546 _8495_/Q vssd1 vssd1 vccd1 vccd1 _4307_/A sky130_fd_sc_hd__buf_1
X_5067_ input25/X _5391_/A _5067_/S vssd1 vssd1 vccd1 vccd1 _5068_/B sky130_fd_sc_hd__mux2_1
Xhold1568 hold1823/X vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5273__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1579 _7640_/Q vssd1 vssd1 vccd1 vccd1 _4222_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4018_ _4752_/B _3676_/A _4082_/B1 _4011_/X _4017_/X vssd1 vssd1 vccd1 vccd1 _5974_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA_fanout465_A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5812__A2 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5969_ _5959_/X _5960_/X _5967_/X _5968_/Y vssd1 vssd1 vccd1 vccd1 _7875_/D sky130_fd_sc_hd__o31a_1
XFILLER_0_66_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6773__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7708_ _8464_/CLK _7708_/D vssd1 vssd1 vccd1 vccd1 _7708_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4921__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5328__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7639_ _8507_/CLK _7639_/D vssd1 vssd1 vccd1 vccd1 _7639_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6421__B _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1747_A _7357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6828__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3780__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4934__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5264__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5500__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3939__C _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5016__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6764__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4831__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3955__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5319__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6331__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold109 _6509_/X vssd1 vssd1 vccd1 vccd1 _7991_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5255__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7990_ _8195_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _7990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6941_ _6941_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6941_/X sky130_fd_sc_hd__and2_1
XANTENNA__3805__B2 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6872_ _7019_/A _6872_/A2 _6845_/B _6871_/X vssd1 vssd1 vccd1 vccd1 _6872_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6755__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5823_ _5823_/A _5823_/B vssd1 vssd1 vccd1 vccd1 _5823_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_76_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6204__C1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5837__S _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6522__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5754_ _5950_/S _5753_/Y _5750_/Y vssd1 vssd1 vccd1 vccd1 _5754_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8473_ _8473_/CLK _8473_/D vssd1 vssd1 vccd1 vccd1 _8473_/Q sky130_fd_sc_hd__dfxtp_1
X_5685_ _6524_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5685_/X sky130_fd_sc_hd__and2_1
X_4705_ _8192_/Q _8224_/Q _8288_/Q _7796_/Q _4706_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4705_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4042__A _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout213_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4636_ _8472_/Q _8404_/Q _8436_/Q _8310_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4636_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7424_ _8471_/CLK _7424_/D vssd1 vssd1 vccd1 vccd1 _7424_/Q sky130_fd_sc_hd__dfxtp_1
X_7355_ _8454_/CLK _7355_/D vssd1 vssd1 vccd1 vccd1 _7355_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold621 _7415_/Q vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold610 _5213_/X vssd1 vssd1 vccd1 vccd1 _7427_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4567_ _4566_/X _4565_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4567_/X sky130_fd_sc_hd__mux2_1
Xhold643 _8311_/Q vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
X_6306_ _6412_/S _6302_/Y _6305_/Y _5740_/Y _6000_/X vssd1 vssd1 vccd1 vccd1 _6306_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3881__A _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold632 _6693_/X vssd1 vssd1 vccd1 vccd1 _8220_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold654 _6736_/X vssd1 vssd1 vccd1 vccd1 _8291_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 _7480_/Q vssd1 vssd1 vccd1 vccd1 hold665/X sky130_fd_sc_hd__dlygate4sd3_1
X_7286_ _8387_/CLK _7286_/D _7096_/Y vssd1 vssd1 vccd1 vccd1 _7286_/Q sky130_fd_sc_hd__dfrtp_4
Xhold687 _8463_/Q vssd1 vssd1 vccd1 vccd1 _7005_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold676 _6758_/X vssd1 vssd1 vccd1 vccd1 _8309_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _5156_/A1 _4406_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _7300_/D sky130_fd_sc_hd__mux2_1
Xhold698 _7004_/X vssd1 vssd1 vccd1 vccd1 _8462_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ _6302_/A _6083_/A _5907_/X _5740_/Y vssd1 vssd1 vccd1 vccd1 _6237_/X sky130_fd_sc_hd__o31a_1
XANTENNA__4916__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6168_ _6391_/A _6159_/X _6167_/Y vssd1 vssd1 vccd1 vccd1 _6168_/Y sky130_fd_sc_hd__o21ai_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1310 _8176_/Q vssd1 vssd1 vccd1 vccd1 _6624_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5119_ _7074_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _5119_/X sky130_fd_sc_hd__or2_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 _6612_/X vssd1 vssd1 vccd1 vccd1 _8170_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1343 _6814_/X vssd1 vssd1 vccd1 vccd1 _8344_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1332 _8352_/Q vssd1 vssd1 vccd1 vccd1 _6830_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1365 hold883/X vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__clkbuf_2
Xhold1376 _7067_/Y vssd1 vssd1 vccd1 vccd1 _7068_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_6099_ _6035_/A _6056_/A _6075_/A _6096_/A _5782_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6099_/X sky130_fd_sc_hd__mux4_2
XANTENNA__5246__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1354 _8341_/Q vssd1 vssd1 vccd1 vccd1 _6808_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1387 _5544_/X vssd1 vssd1 vccd1 vccd1 _7733_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1398 _8368_/Q vssd1 vssd1 vccd1 vccd1 _5024_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6746__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4651__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6432__A _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5990__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7263__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3911__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6607__A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5237__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4561__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6737__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5960__A1 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5960__B2 _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3685__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5470_ _5470_/A _5470_/B _5470_/C vssd1 vssd1 vccd1 vccd1 _5470_/X sky130_fd_sc_hd__and3_1
X_4421_ _4421_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4421_/X sky130_fd_sc_hd__and2_1
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5712__A1 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7171__49 _8475_/CLK vssd1 vssd1 vccd1 vccd1 _8051_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4352_ _4352_/A _4352_/B vssd1 vssd1 vccd1 vccd1 _4352_/X sky130_fd_sc_hd__xor2_1
X_7071_ _7071_/A _7071_/B vssd1 vssd1 vccd1 vccd1 _7071_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__6268__A2 _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout419 hold1747/X vssd1 vssd1 vccd1 vccd1 _7063_/A sky130_fd_sc_hd__buf_8
Xfanout408 _7061_/A vssd1 vssd1 vccd1 vccd1 _4976_/S1 sky130_fd_sc_hd__buf_4
X_4283_ _4407_/A _4404_/B _4283_/C vssd1 vssd1 vccd1 vccd1 _4401_/A sky130_fd_sc_hd__and3_1
X_6022_ _4045_/A _6105_/A2 _6020_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _6023_/C sky130_fd_sc_hd__a22o_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6517__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4736__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7973_ _8364_/CLK _7973_/D vssd1 vssd1 vccd1 vccd1 _7973_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5779__A1 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6924_ _7026_/A _6924_/A2 _6970_/A3 _6923_/X vssd1 vssd1 vccd1 vccd1 _6924_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout163_A _5002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6855_ _6921_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6855_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6728__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3998_ _7283_/Q _7949_/Q vssd1 vssd1 vccd1 vccd1 _3998_/X sky130_fd_sc_hd__and2b_1
XANTENNA_fanout330_A _6915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5806_ _6008_/A _5806_/B vssd1 vssd1 vccd1 vccd1 _5811_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout428_A _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6786_ _7025_/A _6786_/A2 _6838_/A3 _6785_/X vssd1 vssd1 vccd1 vccd1 _6786_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_134_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7067__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5737_ _5738_/A _5738_/B vssd1 vssd1 vccd1 vccd1 _5740_/B sky130_fd_sc_hd__and2_4
XFILLER_0_72_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8456_ _8456_/CLK _8456_/D vssd1 vssd1 vccd1 vccd1 _8456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5668_ _6552_/A _5668_/B vssd1 vssd1 vccd1 vccd1 _5668_/X sky130_fd_sc_hd__and2_1
XFILLER_0_115_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7407_ _8338_/CLK _7407_/D vssd1 vssd1 vccd1 vccd1 _7407_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5599_ _6935_/A _5584_/B _5617_/B1 _5599_/B2 vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__a22o_1
X_4619_ _8147_/Q _7546_/Q _7418_/Q _7578_/Q _4696_/S0 _4737_/S1 vssd1 vssd1 vccd1
+ vccd1 _4619_/X sky130_fd_sc_hd__mux4_1
X_8387_ _8387_/CLK _8387_/D _7281_/Y vssd1 vssd1 vccd1 vccd1 _8387_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold440 _6719_/X vssd1 vssd1 vccd1 vccd1 _8274_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold451 _8211_/Q vssd1 vssd1 vccd1 vccd1 hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _6695_/X vssd1 vssd1 vccd1 vccd1 _8222_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7338_ _8033_/CLK _7338_/D vssd1 vssd1 vccd1 vccd1 _7338_/Q sky130_fd_sc_hd__dfxtp_1
Xhold484 _6745_/X vssd1 vssd1 vccd1 vccd1 _8296_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _7409_/Q vssd1 vssd1 vccd1 vccd1 hold473/X sky130_fd_sc_hd__dlygate4sd3_1
X_7269_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7269_/Y sky130_fd_sc_hd__inv_2
Xhold495 _7788_/Q vssd1 vssd1 vccd1 vccd1 hold495/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6427__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1140 _6922_/X vssd1 vssd1 vccd1 vccd1 _8426_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1151 _8429_/Q vssd1 vssd1 vccd1 vccd1 _6928_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5219__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1184 _6862_/X vssd1 vssd1 vccd1 vccd1 _8397_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 _8401_/Q vssd1 vssd1 vccd1 vccd1 _6870_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _6822_/X vssd1 vssd1 vccd1 vccd1 _8348_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1195 _8172_/Q vssd1 vssd1 vccd1 vccd1 _6616_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6719__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7258__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3786__A _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__A1 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3953__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5170__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5856__S1 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7216__94 _8500_/CLK vssd1 vssd1 vccd1 vccd1 _8129_/CLK sky130_fd_sc_hd__inv_2
X_4970_ _4969_/X _4968_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3921_ _5820_/A _5879_/S vssd1 vssd1 vccd1 vccd1 _3922_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6186__B2 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6186__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3852_ _3852_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3852_/X sky130_fd_sc_hd__or2_1
X_6640_ _7028_/A _6640_/A2 _6666_/A3 _6639_/X vssd1 vssd1 vccd1 vccd1 _6640_/X sky130_fd_sc_hd__a31o_1
X_6571_ _6929_/A _6592_/A2 _6592_/B1 hold837/X vssd1 vssd1 vccd1 vccd1 _6571_/X sky130_fd_sc_hd__a22o_1
X_8310_ _8472_/CLK _8310_/D vssd1 vssd1 vccd1 vccd1 _8310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5522_ _8241_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7711_/D sky130_fd_sc_hd__and3_1
X_3783_ _3783_/A1 _4073_/A2 _3779_/X _4073_/B2 _3782_/X vssd1 vssd1 vccd1 vccd1 _3783_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_131_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5453_ _5453_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5453_/X sky130_fd_sc_hd__and3_1
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8241_ _8241_/CLK _8241_/D vssd1 vssd1 vccd1 vccd1 _8241_/Q sky130_fd_sc_hd__dfxtp_1
X_8172_ _8462_/CLK _8172_/D vssd1 vssd1 vccd1 vccd1 _8172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5384_ _7067_/A _7069_/A _6597_/B _5382_/X vssd1 vssd1 vccd1 vccd1 _5384_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_41_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4404_ _4407_/A _4404_/B vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__or2_1
XANTENNA__5135__B _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _6250_/S vssd1 vssd1 vccd1 vccd1 _6411_/S sky130_fd_sc_hd__buf_4
X_7123_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7123_/Y sky130_fd_sc_hd__inv_2
X_4335_ _4335_/A _4336_/B vssd1 vssd1 vccd1 vccd1 _4335_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout238 _5085_/B vssd1 vssd1 vccd1 vccd1 _4448_/B sky130_fd_sc_hd__buf_4
Xfanout227 _7073_/B vssd1 vssd1 vccd1 vccd1 _5449_/C sky130_fd_sc_hd__buf_4
Xfanout216 _5456_/C vssd1 vssd1 vccd1 vccd1 _5540_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7054_ hold89/X _7069_/B vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__nand2_1
Xfanout249 _6669_/Y vssd1 vssd1 vccd1 vccd1 _6701_/B1 sky130_fd_sc_hd__buf_8
X_4266_ _4256_/Y _4260_/B _4258_/B vssd1 vssd1 vccd1 vccd1 _4267_/B sky130_fd_sc_hd__o21a_1
XANTENNA_fanout280_A _6842_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6005_ _6005_/A _6005_/B vssd1 vssd1 vccd1 vccd1 _6005_/Y sky130_fd_sc_hd__nor2_1
X_4197_ _4186_/Y _4189_/X _4188_/B vssd1 vssd1 vccd1 vccd1 _4197_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout378_A _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6964__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7956_ _8020_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 _7956_/Q sky130_fd_sc_hd__dfxtp_1
X_6907_ _7939_/Q _7940_/Q _6908_/C vssd1 vssd1 vccd1 vccd1 _6971_/B sky130_fd_sc_hd__nor3_4
X_7887_ _8419_/CLK _7887_/D vssd1 vssd1 vccd1 vccd1 _7887_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7078__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6838_ _7023_/A _6838_/A2 _6838_/A3 _6837_/X vssd1 vssd1 vccd1 vccd1 _6838_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_92_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8508_ _8519_/CLK _8508_/D vssd1 vssd1 vccd1 vccd1 _8508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6769_ _6961_/A _6773_/A2 _6773_/B1 hold933/X vssd1 vssd1 vccd1 vccd1 _6769_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6024__S1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8439_ _8475_/CLK _8439_/D vssd1 vssd1 vccd1 vccd1 _8439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4586__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold270 _7379_/Q vssd1 vssd1 vccd1 vccd1 _5446_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _6564_/X vssd1 vssd1 vccd1 vccd1 _8136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _7320_/Q vssd1 vssd1 vccd1 vccd1 _5417_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6157__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5612__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7230__108 _8332_/CLK vssd1 vssd1 vccd1 vccd1 _8240_/CLK sky130_fd_sc_hd__inv_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6168__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3926__B1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5915__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5915__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6340__A1 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7141__19 _8450_/CLK vssd1 vssd1 vccd1 vccd1 _7518_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4577__S1 _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4120_ _3818_/Y _6352_/A _3848_/C _3833_/Y _6370_/A vssd1 vssd1 vccd1 vccd1 _4120_/X
+ sky130_fd_sc_hd__o32a_1
X_4051_ _4758_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _4051_/X sky130_fd_sc_hd__and2_1
XFILLER_0_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput5 i_instr_ID[14] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5851__B1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7810_ _8428_/CLK _7810_/D vssd1 vssd1 vccd1 vccd1 _7810_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5603__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7741_ _8362_/CLK _7741_/D vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
X_4953_ _4951_/X _4952_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6946__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3904_ _3904_/A1 _4084_/A2 _6849_/A _4084_/B2 _3903_/X vssd1 vssd1 vccd1 vccd1 _3904_/Y
+ sky130_fd_sc_hd__a221oi_4
X_7672_ _8195_/CLK _7672_/D vssd1 vssd1 vccd1 vccd1 _7672_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6623_ _6929_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6623_/X sky130_fd_sc_hd__and2_1
XFILLER_0_6_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4884_ _8181_/Q _8213_/Q _8277_/Q _7785_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4884_/X sky130_fd_sc_hd__mux4_1
X_3835_ _6370_/A _6367_/A vssd1 vssd1 vccd1 vccd1 _3836_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_132_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6554_ _7079_/C _6554_/B _6554_/C _6554_/D vssd1 vssd1 vccd1 vccd1 _6554_/X sky130_fd_sc_hd__and4_1
XANTENNA__3917__B1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6530__A _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3766_ _7988_/Q _4068_/A2 _4068_/B1 _8020_/Q _3765_/X vssd1 vssd1 vccd1 vccd1 _3766_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_131_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6485_ _6520_/A hold61/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__and2_1
XANTENNA__4135__A_N _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5505_ _7526_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7694_/D sky130_fd_sc_hd__and3_1
X_3697_ _7662_/Q _7939_/Q vssd1 vssd1 vccd1 vccd1 _3697_/X sky130_fd_sc_hd__and2b_1
X_5436_ _5436_/A _5470_/B _5468_/C vssd1 vssd1 vccd1 vccd1 _5436_/X sky130_fd_sc_hd__and3_1
X_8224_ _8353_/CLK _8224_/D vssd1 vssd1 vccd1 vccd1 _8224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5134__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8155_ _8354_/CLK _8155_/D vssd1 vssd1 vccd1 vccd1 _8155_/Q sky130_fd_sc_hd__dfxtp_1
X_5367_ _6969_/A _5367_/A2 _5367_/B1 hold553/X vssd1 vssd1 vccd1 vccd1 _5367_/X sky130_fd_sc_hd__a22o_1
X_7106_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7106_/Y sky130_fd_sc_hd__inv_2
X_5298_ _6558_/A _6842_/C vssd1 vssd1 vccd1 vccd1 _5300_/B sky130_fd_sc_hd__or2_1
X_8086_ _8086_/CLK _8120_/D vssd1 vssd1 vccd1 vccd1 _8086_/Q sky130_fd_sc_hd__dfxtp_1
X_4318_ _4318_/A vssd1 vssd1 vccd1 vccd1 _4318_/Y sky130_fd_sc_hd__inv_2
X_7037_ _7031_/Y _7037_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8491_/D sky130_fd_sc_hd__a21oi_1
X_4249_ _4250_/A _7644_/Q vssd1 vssd1 vccd1 vccd1 _4249_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4740__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6705__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7939_ _8456_/CLK _7939_/D vssd1 vssd1 vccd1 vccd1 _7939_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6570__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6440__A _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4559__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6322__A1 _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7271__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6086__B1 _5732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5503__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5833__A0 _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4731__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6615__A _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4834__S _7359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6928__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3974__A _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4798__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6561__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5967__A1_N _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5364__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5116__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6270_ _6270_/A _6270_/B vssd1 vssd1 vccd1 vccd1 _6270_/X sky130_fd_sc_hd__or2_1
XANTENNA__3913__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5221_ _6971_/A _5221_/A2 _5221_/B1 hold917/X vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__a22o_1
X_5152_ _5152_/A1 _4407_/B _5166_/B1 _5151_/X vssd1 vssd1 vccd1 vccd1 _7388_/D sky130_fd_sc_hd__o211a_1
X_4103_ _3962_/X _4102_/X _4100_/Y vssd1 vssd1 vccd1 vccd1 _4103_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5413__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1717 _8502_/Q vssd1 vssd1 vccd1 vccd1 _3774_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1706 _4315_/Y vssd1 vssd1 vccd1 vccd1 _4317_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5083_ _7069_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5083_/X sky130_fd_sc_hd__or2_1
Xhold1728 _4225_/X vssd1 vssd1 vccd1 vccd1 _5561_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1739 _8511_/Q vssd1 vssd1 vccd1 vccd1 _4014_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5824__B1 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4034_ _7980_/Q _4079_/A2 _4079_/B1 _8012_/Q _4033_/X vssd1 vssd1 vccd1 vccd1 _4034_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6525__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3850__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3868__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5985_ _5703_/X _5711_/X _6028_/S vssd1 vssd1 vccd1 vccd1 _5985_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7724_ _8195_/CLK _7724_/D vssd1 vssd1 vccd1 vccd1 _7724_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout243_A _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4936_ _4935_/X _4932_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8252_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4867_ _8339_/Q _7815_/Q _7481_/Q _7449_/Q _4896_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4867_/X sky130_fd_sc_hd__mux4_1
XANTENNA_21 _7289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7655_ _8494_/CLK hold64/X vssd1 vssd1 vccd1 vccd1 _7655_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_10 _7904_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6606_ _6999_/A _6606_/A2 _6602_/X _6605_/Y vssd1 vssd1 vccd1 vccd1 _6606_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout410_A _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _6350_/A vssd1 vssd1 vccd1 vccd1 _3818_/Y sky130_fd_sc_hd__inv_2
X_7586_ _8484_/CLK _7586_/D vssd1 vssd1 vccd1 vccd1 _7586_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6260__A _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5355__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4798_ _8136_/Q _7535_/Q _7407_/Q _7567_/Q _4896_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4798_/X sky130_fd_sc_hd__mux4_1
X_6537_ _7022_/A _6537_/B vssd1 vssd1 vccd1 vccd1 _8019_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3749_ _3749_/A _3749_/B vssd1 vssd1 vccd1 vccd1 _4138_/A sky130_fd_sc_hd__and2_1
X_6468_ _6999_/A hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_63_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5419_ _5419_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5419_/X sky130_fd_sc_hd__and3_1
X_8207_ _8425_/CLK _8207_/D vssd1 vssd1 vccd1 vccd1 _8207_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput150 _8065_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[30] sky130_fd_sc_hd__buf_12
X_6399_ _3848_/A _6414_/A2 _5926_/Y _6309_/Y _6398_/X vssd1 vssd1 vccd1 vccd1 _6399_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8138_ _8154_/CLK _8138_/D vssd1 vssd1 vccd1 vccd1 _8138_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_78_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4961__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8069_ _8328_/CLK _8069_/D vssd1 vssd1 vccd1 vccd1 _8069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5291__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4713__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5830__A3 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6435__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6154__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5594__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_16_clk_A _7871_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5346__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7266__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _7871_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4952__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7236__114 _8413_/CLK vssd1 vssd1 vccd1 vccd1 _8246_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4564__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5282__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6231__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6782__A1 _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5770_ _3950_/X _6398_/A2 _6413_/B1 _5797_/S _6011_/A2 vssd1 vssd1 vccd1 vccd1 _5770_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4721_ _4720_/X _4719_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7440_ _8350_/CLK _7440_/D vssd1 vssd1 vccd1 vccd1 _7440_/Q sky130_fd_sc_hd__dfxtp_1
X_4652_ _4651_/X _4648_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7518_/D sky130_fd_sc_hd__mux2_1
Xinput30 i_instr_ID[9] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5408__B _5408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4640__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4583_ _8335_/Q _7811_/Q _7477_/Q _7445_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4583_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3899__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput63 rst vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_8
Xhold803 _8223_/Q vssd1 vssd1 vccd1 vccd1 hold803/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput52 i_read_data_M[29] vssd1 vssd1 vccd1 vccd1 _6550_/B sky130_fd_sc_hd__clkbuf_1
Xinput41 i_read_data_M[19] vssd1 vssd1 vccd1 vccd1 _6540_/B sky130_fd_sc_hd__clkbuf_1
X_7371_ _8008_/CLK _7371_/D vssd1 vssd1 vccd1 vccd1 _7371_/Q sky130_fd_sc_hd__dfxtp_1
Xhold836 _5635_/X vssd1 vssd1 vccd1 vccd1 _7815_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 _7807_/Q vssd1 vssd1 vccd1 vccd1 hold825/X sky130_fd_sc_hd__dlygate4sd3_1
X_6322_ _6298_/A _6318_/A _6262_/A _6281_/A _5772_/S _5838_/A vssd1 vssd1 vccd1 vccd1
+ _6393_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_24_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold814 _5364_/X vssd1 vssd1 vccd1 vccd1 _7591_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 _5200_/X vssd1 vssd1 vccd1 vccd1 _7414_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4739__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6253_ _6412_/S _5930_/B _6128_/X vssd1 vssd1 vccd1 vccd1 _6253_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold847 _8482_/Q vssd1 vssd1 vccd1 vccd1 _7024_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 _8156_/Q vssd1 vssd1 vccd1 vccd1 hold869/X sky130_fd_sc_hd__dlygate4sd3_1
X_5204_ _6937_/A _5221_/A2 _5221_/B1 hold751/X vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5143__B _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6184_ _3800_/C _6414_/A2 _6182_/X _6309_/A _6183_/X vssd1 vssd1 vccd1 vccd1 _6184_/X
+ sky130_fd_sc_hd__a221o_1
Xhold1514 _8329_/Q vssd1 vssd1 vccd1 vccd1 _6783_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5135_ _5447_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__or2_1
Xhold1525 hold1821/X vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__buf_1
Xhold1503 _7297_/Q vssd1 vssd1 vccd1 vccd1 _5150_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1558 _7641_/Q vssd1 vssd1 vccd1 vccd1 _4229_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1536 _4187_/Y vssd1 vssd1 vccd1 vccd1 _4188_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5066_ input24/X _5067_/S _5172_/B1 _5065_/X vssd1 vssd1 vccd1 vccd1 _7345_/D sky130_fd_sc_hd__o211a_1
Xhold1547 _4307_/Y vssd1 vssd1 vccd1 vccd1 _4308_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5273__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4017_ _7708_/Q _4081_/B vssd1 vssd1 vccd1 vccd1 _4017_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout360_A _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1569 hold1820/X vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__buf_1
XANTENNA_fanout458_A _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5968_ _3985_/B _6063_/A _7258_/A vssd1 vssd1 vccd1 vccd1 _5968_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6773__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7177__55 _8457_/CLK vssd1 vssd1 vccd1 vccd1 _8057_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_75_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7707_ _8173_/CLK _7707_/D vssd1 vssd1 vccd1 vccd1 _7707_/Q sky130_fd_sc_hd__dfxtp_1
X_4919_ _8186_/Q _8218_/Q _8282_/Q _7790_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4919_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_118_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7086__A _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5899_ _6411_/S _5899_/B vssd1 vssd1 vccd1 vccd1 _5900_/C sky130_fd_sc_hd__nor2_1
X_7638_ _8510_/CLK _7638_/D vssd1 vssd1 vccd1 vccd1 _7638_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5328__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7569_ _8461_/CLK _7569_/D vssd1 vssd1 vccd1 vccd1 _7569_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4934__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5264__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4698__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5500__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6764__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4870__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3728__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5319__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4622__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output87_A _8131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3971__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5255__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4689__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6940_ _6434_/A _6940_/A2 _6970_/A3 _6939_/X vssd1 vssd1 vccd1 vccd1 _6940_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3805__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6871_ _6937_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6871_/X sky130_fd_sc_hd__and2_1
XFILLER_0_44_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5822_ _5820_/X _5822_/B vssd1 vssd1 vccd1 vccd1 _5823_/B sky130_fd_sc_hd__and2b_1
X_5753_ _6126_/A _5838_/A _5752_/X vssd1 vssd1 vccd1 vccd1 _5753_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4861__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4704_ _4702_/X _4703_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4704_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8472_ _8472_/CLK _8472_/D vssd1 vssd1 vccd1 vccd1 _8472_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5684_ _6520_/A hold51/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__and2_1
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4635_ _8182_/Q _8214_/Q _8278_/Q _7786_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4635_/X sky130_fd_sc_hd__mux4_1
X_7423_ _8445_/CLK _7423_/D vssd1 vssd1 vccd1 vccd1 _7423_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7354_ _7907_/CLK _7354_/D vssd1 vssd1 vccd1 vccd1 _7354_/Q sky130_fd_sc_hd__dfxtp_1
X_4566_ _8462_/Q _8394_/Q _8426_/Q _8300_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4566_/X sky130_fd_sc_hd__mux4_1
Xhold611 _7782_/Q vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold600 _6766_/X vssd1 vssd1 vccd1 vccd1 _8317_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 _6760_/X vssd1 vssd1 vccd1 vccd1 _8311_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _8164_/Q vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ _6411_/S _6305_/B vssd1 vssd1 vccd1 vccd1 _6305_/Y sky130_fd_sc_hd__nand2_1
Xhold622 _5201_/X vssd1 vssd1 vccd1 vccd1 _7415_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold666 _5276_/X vssd1 vssd1 vccd1 vccd1 _7480_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7285_ _8362_/CLK _7285_/D _7095_/Y vssd1 vssd1 vccd1 vccd1 _7285_/Q sky130_fd_sc_hd__dfrtp_1
Xhold655 _7784_/Q vssd1 vssd1 vccd1 vccd1 hold655/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 _7458_/Q vssd1 vssd1 vccd1 vccd1 hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 _7005_/X vssd1 vssd1 vccd1 vccd1 _8463_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _5158_/A1 _4404_/B _5468_/C vssd1 vssd1 vccd1 vccd1 _7301_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6236_ _6411_/S _6081_/Y _6235_/Y _6412_/S vssd1 vssd1 vccd1 vccd1 _6236_/X sky130_fd_sc_hd__o211a_1
Xhold699 _7583_/Q vssd1 vssd1 vccd1 vccd1 hold699/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4916__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1300 _8434_/Q vssd1 vssd1 vccd1 vccd1 _6938_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_6167_ _6309_/A _5755_/X _6130_/A vssd1 vssd1 vccd1 vccd1 _6167_/Y sky130_fd_sc_hd__o21ai_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6691__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1311 _6624_/X vssd1 vssd1 vccd1 vccd1 _8176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 _8171_/Q vssd1 vssd1 vccd1 vccd1 _6614_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ input20/X _5067_/S _5172_/B1 _5117_/X vssd1 vssd1 vccd1 vccd1 _7371_/D sky130_fd_sc_hd__o211a_1
Xhold1333 _6830_/X vssd1 vssd1 vccd1 vccd1 _8352_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1377 _7068_/Y vssd1 vssd1 vccd1 vccd1 _8506_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6098_ _6098_/A _6098_/B vssd1 vssd1 vccd1 vccd1 _6098_/Y sky130_fd_sc_hd__xnor2_1
Xhold1344 _8342_/Q vssd1 vssd1 vccd1 vccd1 _6810_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5246__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1366 hold1511/X vssd1 vssd1 vccd1 vccd1 _7075_/A sky130_fd_sc_hd__buf_2
Xhold1355 _6808_/X vssd1 vssd1 vccd1 vccd1 _8341_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1399 _4227_/C vssd1 vssd1 vccd1 vccd1 _4504_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1388 _8382_/Q vssd1 vssd1 vccd1 vccd1 _5052_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ hold98/X _5463_/C vssd1 vssd1 vccd1 vccd1 _5049_/X sky130_fd_sc_hd__or2_1
XANTENNA__6746__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4932__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4604__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5182__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3732__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6357__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6682__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5237__A1 _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5511__B _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5003__S _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6623__A _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6737__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3966__B _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4843__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4420_ hold637/X _4425_/B _4420_/B1 _4419_/Y vssd1 vssd1 vccd1 vccd1 _8370_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4351_ _4342_/Y _4346_/B _4351_/B1 vssd1 vssd1 vccd1 vccd1 _4351_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_10_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7070_ _7071_/B _7070_/A2 _7090_/A vssd1 vssd1 vccd1 vccd1 _7070_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__6268__A3 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout409 hold1729/X vssd1 vssd1 vccd1 vccd1 _7061_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4282_ _4281_/X _5040_/A1 _5465_/B vssd1 vssd1 vccd1 vccd1 _4283_/C sky130_fd_sc_hd__mux2_1
X_6021_ _4008_/A _6398_/A2 _6413_/B1 _6013_/A vssd1 vssd1 vccd1 vccd1 _6023_/B sky130_fd_sc_hd__a22o_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5228__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5421__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7972_ _8519_/CLK _7972_/D vssd1 vssd1 vccd1 vccd1 _7972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6923_ _6923_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6923_/X sky130_fd_sc_hd__and2_1
XANTENNA__6728__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6854_ _7019_/A _6854_/A2 _6845_/B _6853_/X vssd1 vssd1 vccd1 vccd1 _6854_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3876__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3997_ _3973_/X _3974_/Y _3985_/X _3996_/X _3962_/X vssd1 vssd1 vccd1 vccd1 _4092_/B
+ sky130_fd_sc_hd__a2111o_1
X_5805_ _5952_/A _5926_/B _5803_/Y vssd1 vssd1 vccd1 vccd1 _5806_/B sky130_fd_sc_hd__a21oi_1
X_6785_ _6917_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6785_/X sky130_fd_sc_hd__and2_1
XFILLER_0_134_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5736_ _3935_/X _5728_/Y _5735_/X vssd1 vssd1 vccd1 vccd1 _5736_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7147__25 _8195_/CLK vssd1 vssd1 vccd1 vccd1 _7524_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5667_ _5667_/A _5667_/B vssd1 vssd1 vccd1 vccd1 _5667_/X sky130_fd_sc_hd__and2_1
X_8455_ _8515_/CLK _8455_/D vssd1 vssd1 vccd1 vccd1 _8455_/Q sky130_fd_sc_hd__dfxtp_1
X_7406_ _8338_/CLK _7406_/D vssd1 vssd1 vccd1 vccd1 _7406_/Q sky130_fd_sc_hd__dfxtp_1
X_4618_ _8340_/Q _7816_/Q _7482_/Q _7450_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4618_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_60_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5164__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5598_ _6933_/A _5584_/B _5617_/B1 hold611/X vssd1 vssd1 vccd1 vccd1 _5598_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_102_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8386_ _8387_/CLK _8386_/D _7280_/Y vssd1 vssd1 vccd1 vccd1 _8386_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__6900__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold463 _7533_/Q vssd1 vssd1 vccd1 vccd1 hold463/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4199__S _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 _6684_/X vssd1 vssd1 vccd1 vccd1 _8211_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 _7585_/Q vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _5249_/X vssd1 vssd1 vccd1 vccd1 _7457_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6169__B1_N _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4549_ _8137_/Q _7536_/Q _7408_/Q _7568_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4549_/X sky130_fd_sc_hd__mux4_1
X_7337_ _8382_/CLK _7337_/D vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold474 _5195_/X vssd1 vssd1 vccd1 vccd1 _7409_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _8308_/Q vssd1 vssd1 vccd1 vccd1 hold485/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _5604_/X vssd1 vssd1 vccd1 vccd1 _7788_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7268_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7268_/Y sky130_fd_sc_hd__inv_2
X_6219_ _3872_/A _6414_/B1 _6398_/B1 _3871_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6219_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_hold1605_A _7345_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1130 _6914_/X vssd1 vssd1 vccd1 vccd1 _8422_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 _8351_/Q vssd1 vssd1 vccd1 vccd1 _6828_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5219__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1152 _6928_/X vssd1 vssd1 vccd1 vccd1 _8429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1174 _6870_/X vssd1 vssd1 vccd1 vccd1 _8401_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 _8399_/Q vssd1 vssd1 vccd1 vccd1 _6866_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 _8431_/Q vssd1 vssd1 vccd1 vccd1 _6932_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1196 _6616_/X vssd1 vssd1 vccd1 vccd1 _8172_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4662__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6443__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6195__A2 _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4825__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3953__B2 _8009_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7274__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4410__B _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5506__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4837__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4130__B2 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5630__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _4014_/A _3917_/Y _3918_/Y vssd1 vssd1 vccd1 vccd1 _3920_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6072__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3851_ _8089_/Q _3850_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3851_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_132_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6570_ _6927_/A _6592_/A2 _6592_/B1 _6570_/B2 vssd1 vssd1 vccd1 vccd1 _6570_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3782_ _4762_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__and2_1
X_5521_ _8240_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7710_/D sky130_fd_sc_hd__and3_1
XANTENNA__5933__A2 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8240_ _8240_/CLK _8240_/D vssd1 vssd1 vccd1 vccd1 _8240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5452_ _5452_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5452_/X sky130_fd_sc_hd__and3_1
XANTENNA__5146__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8171_ _8461_/CLK _8171_/D vssd1 vssd1 vccd1 vccd1 _8171_/Q sky130_fd_sc_hd__dfxtp_1
X_5383_ _7065_/A _5395_/A vssd1 vssd1 vccd1 vccd1 _6597_/B sky130_fd_sc_hd__nand2_2
XANTENNA__5416__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4403_ _4403_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _4403_/X sky130_fd_sc_hd__and2_1
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7122_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7122_/Y sky130_fd_sc_hd__inv_2
X_4334_ _4383_/A _4383_/B vssd1 vssd1 vccd1 vccd1 _4334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout228 _7073_/B vssd1 vssd1 vccd1 vccd1 _7088_/B sky130_fd_sc_hd__buf_4
Xfanout206 _6250_/S vssd1 vssd1 vccd1 vccd1 _6342_/S sky130_fd_sc_hd__clkbuf_8
X_7053_ _7031_/Y _7052_/X _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8499_/D sky130_fd_sc_hd__a21oi_1
Xfanout217 _5465_/C vssd1 vssd1 vccd1 vccd1 _5463_/C sky130_fd_sc_hd__buf_4
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout239 _5099_/B vssd1 vssd1 vccd1 vccd1 _5085_/B sky130_fd_sc_hd__clkbuf_4
X_6004_ _6105_/A2 _5996_/A _6002_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6005_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_66_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4265_ _4263_/Y _4265_/B vssd1 vssd1 vccd1 vccd1 _4265_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6528__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4196_ _4194_/Y _4196_/B vssd1 vssd1 vccd1 vccd1 _4198_/A sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout273_A _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7955_ _8019_/CLK _7955_/D vssd1 vssd1 vccd1 vccd1 _7955_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6906_ _7026_/A _6906_/A2 _6906_/A3 _6905_/X vssd1 vssd1 vccd1 vccd1 _6906_/X sky130_fd_sc_hd__a31o_1
X_7886_ _8427_/CLK _7886_/D vssd1 vssd1 vccd1 vccd1 _7886_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout440_A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6837_ _6969_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6837_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4807__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8507_ _8507_/CLK _8507_/D vssd1 vssd1 vccd1 vccd1 _8507_/Q sky130_fd_sc_hd__dfxtp_1
X_6768_ _6959_/A _6773_/A2 _6773_/B1 hold477/X vssd1 vssd1 vccd1 vccd1 _6768_/X sky130_fd_sc_hd__a22o_1
X_5719_ _5711_/X _5718_/X _6028_/S vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__mux2_2
X_6699_ _6965_/A _6701_/A2 _6701_/B1 hold569/X vssd1 vssd1 vccd1 vccd1 _6699_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3826__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8438_ _8476_/CLK _8438_/D vssd1 vssd1 vccd1 vccd1 _8438_/Q sky130_fd_sc_hd__dfxtp_1
X_8369_ _8369_/CLK _8369_/D _7263_/Y vssd1 vssd1 vccd1 vccd1 _8369_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold260 _7772_/Q vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _5446_/X vssd1 vssd1 vccd1 vccd1 _7635_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _5417_/X vssd1 vssd1 vccd1 vccd1 _7606_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _7374_/Q vssd1 vssd1 vccd1 vccd1 _5441_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6652__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5061__B _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7062__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3797__A _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5612__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7269__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6173__A _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6901__A _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3926__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5128__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6340__A2 _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4567__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4050_ _4758_/B _3676_/A _4082_/B1 _4048_/X _4049_/X vssd1 vssd1 vccd1 vccd1 _6096_/A
+ sky130_fd_sc_hd__o221a_4
Xinput6 i_instr_ID[15] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__7053__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5603__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7740_ _8364_/CLK _7740_/D vssd1 vssd1 vccd1 vccd1 _7740_/Q sky130_fd_sc_hd__dfxtp_1
X_4952_ _8158_/Q _7557_/Q _7429_/Q _7589_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4952_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7671_ _8328_/CLK _7671_/D vssd1 vssd1 vccd1 vccd1 _7671_/Q sky130_fd_sc_hd__dfxtp_1
X_3903_ hold5/X _4083_/B vssd1 vssd1 vccd1 vccd1 _3903_/X sky130_fd_sc_hd__and2_1
XFILLER_0_74_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4883_ _4881_/X _4882_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__mux2_1
X_6622_ _7007_/A _6622_/A2 _6605_/B _6621_/X vssd1 vssd1 vccd1 vccd1 _6622_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_86_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3834_ _6370_/A _6367_/A vssd1 vssd1 vccd1 vccd1 _3836_/A sky130_fd_sc_hd__or2_1
XANTENNA__5367__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6811__A _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6553_ _6553_/A _6553_/B vssd1 vssd1 vccd1 vccd1 _6554_/D sky130_fd_sc_hd__nand2_1
XANTENNA__3917__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3765_ _4067_/A_N _7956_/Q vssd1 vssd1 vccd1 vccd1 _3765_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3696_ _3696_/A _3696_/B _3696_/C vssd1 vssd1 vccd1 vccd1 _3696_/Y sky130_fd_sc_hd__nor3_1
X_5504_ _7525_/Q _5538_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7693_/D sky130_fd_sc_hd__and3_1
X_6484_ _6524_/A _6484_/B vssd1 vssd1 vccd1 vccd1 _6484_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8223_ _8319_/CLK _8223_/D vssd1 vssd1 vccd1 vccd1 _8223_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5435_ _5435_/A _5465_/B _5463_/C vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__and3_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8154_ _8154_/CLK _8154_/D vssd1 vssd1 vccd1 vccd1 _8154_/Q sky130_fd_sc_hd__dfxtp_1
X_5366_ _6967_/A _5367_/A2 _5367_/B1 hold769/X vssd1 vssd1 vccd1 vccd1 _5366_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6882__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5297_ _6558_/A _6842_/C vssd1 vssd1 vccd1 vccd1 _5297_/Y sky130_fd_sc_hd__nor2_2
X_7105_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7105_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8085_ _8463_/CLK _8085_/D vssd1 vssd1 vccd1 vccd1 _8085_/Q sky130_fd_sc_hd__dfxtp_1
X_4317_ _4317_/A _4317_/B vssd1 vssd1 vccd1 vccd1 _4318_/A sky130_fd_sc_hd__xnor2_1
X_7036_ _7076_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7036_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6634__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4248_ _4419_/A _4415_/B vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__and2_1
XFILLER_0_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4179_ _4174_/Y _4176_/B _4174_/B vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__o21a_1
XANTENNA__3853__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6705__B _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6398__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7938_ _8456_/CLK _7938_/D vssd1 vssd1 vccd1 vccd1 _7938_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5358__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7869_ _8464_/CLK _7869_/D vssd1 vssd1 vccd1 vccd1 _7869_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6570__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6322__A2 _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5833__A1 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7035__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6615__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5597__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5349__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7201__79 _8080_/CLK vssd1 vssd1 vccd1 vccd1 _8114_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6010__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6631__A _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6561__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6010__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3974__B _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6350__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5220_ _6969_/A _5188_/B _5220_/B1 hold735/X vssd1 vssd1 vccd1 vccd1 _5220_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6864__A3 _6842_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5151_ _5455_/A _5540_/C vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__or2_1
XANTENNA__6616__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5082_ input2/X _4448_/B _5140_/B1 _5081_/X vssd1 vssd1 vccd1 vccd1 _7353_/D sky130_fd_sc_hd__o211a_1
X_4102_ _6198_/S _5870_/A _3996_/X _4101_/Y vssd1 vssd1 vccd1 vccd1 _4102_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5413__C _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1707 _4318_/A vssd1 vssd1 vccd1 vccd1 _5574_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4033_ _3923_/B _7948_/Q vssd1 vssd1 vccd1 vccd1 _4033_/X sky130_fd_sc_hd__and2b_1
Xhold1718 _8490_/Q vssd1 vssd1 vccd1 vccd1 _3831_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_47_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1729 _7358_/Q vssd1 vssd1 vccd1 vccd1 hold1729/X sky130_fd_sc_hd__clkbuf_4
X_5984_ _6028_/S _5982_/X _5983_/Y _5740_/B vssd1 vssd1 vccd1 vccd1 _5984_/Y sky130_fd_sc_hd__o211ai_1
XANTENNA__5052__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7723_ _8355_/CLK _7723_/D vssd1 vssd1 vccd1 vccd1 _7723_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4935_ _4934_/X _4933_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__mux2_1
X_4866_ _4865_/X _4862_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8242_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout236_A _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 _8024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6541__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7654_ _8033_/CLK hold66/X vssd1 vssd1 vccd1 vccd1 _7654_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_22 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6605_ _6845_/A _6605_/B vssd1 vssd1 vccd1 vccd1 _6605_/Y sky130_fd_sc_hd__nor2_1
X_4797_ _8329_/Q _7805_/Q _7471_/Q _7439_/Q _4896_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4797_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4012__B1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7585_ _8283_/CLK _7585_/D vssd1 vssd1 vccd1 vccd1 _7585_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3817_ _4335_/A _3816_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6350_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout403_A _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7075__C _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ _6334_/A _6331_/A vssd1 vssd1 vccd1 vccd1 _3749_/B sky130_fd_sc_hd__nand2_1
X_6536_ _7022_/A _6536_/B vssd1 vssd1 vccd1 vccd1 _8018_/D sky130_fd_sc_hd__and2_1
XFILLER_0_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6467_ _6534_/A hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__and2_1
XFILLER_0_101_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3679_ _7282_/Q _3923_/B vssd1 vssd1 vccd1 vccd1 _3679_/X sky130_fd_sc_hd__and2_1
XFILLER_0_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5418_ _5418_/A _5453_/B _5449_/C vssd1 vssd1 vccd1 vccd1 _5418_/X sky130_fd_sc_hd__and3_1
X_8206_ _8270_/CLK _8206_/D vssd1 vssd1 vccd1 vccd1 _8206_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5391__C_N _5408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6398_ _3811_/A _6398_/A2 _6398_/B1 _6386_/A _5734_/X vssd1 vssd1 vccd1 vccd1 _6398_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput151 _8066_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[31] sky130_fd_sc_hd__buf_12
Xoutput140 _8056_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[21] sky130_fd_sc_hd__buf_12
X_5349_ _6933_/A _5335_/B _5368_/B1 _5349_/B2 vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8137_ _8355_/CLK _8137_/D vssd1 vssd1 vccd1 vccd1 _8137_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4000__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4079__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8068_ _8519_/CLK _8102_/D vssd1 vssd1 vccd1 vccd1 _8068_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5620__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7019_ _7019_/A _7019_/B vssd1 vssd1 vccd1 vccd1 _7019_/X sky130_fd_sc_hd__and2_1
XANTENNA__4935__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5291__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6435__B _6435_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4236__A _8505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8388_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6451__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3794__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5751__A0 _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6846__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4845__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5282__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5034__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_41_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _8136_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6361__A _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4720_ _8484_/Q _8416_/Q _8448_/Q _8322_/Q _4720_/S0 _4741_/S1 vssd1 vssd1 vccd1
+ vccd1 _4720_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_17_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4651_ _4650_/X _4649_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4651_/X sky130_fd_sc_hd__mux2_1
Xinput31 i_read_data_M[0] vssd1 vssd1 vccd1 vccd1 _6521_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput20 i_instr_ID[29] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_1
Xinput53 i_read_data_M[2] vssd1 vssd1 vccd1 vccd1 _6523_/B sky130_fd_sc_hd__clkbuf_1
Xinput42 i_read_data_M[1] vssd1 vssd1 vccd1 vccd1 _6522_/B sky130_fd_sc_hd__clkbuf_1
X_4582_ _4581_/X _4578_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7508_/D sky130_fd_sc_hd__mux2_1
X_7370_ _8154_/CLK _7370_/D vssd1 vssd1 vccd1 vccd1 _7370_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4640__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold837 _8143_/Q vssd1 vssd1 vccd1 vccd1 hold837/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold826 _5627_/X vssd1 vssd1 vccd1 vccd1 _7807_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6321_ _6083_/A _6027_/Y _6128_/X vssd1 vssd1 vccd1 vccd1 _6321_/X sky130_fd_sc_hd__o21a_1
Xhold804 _6696_/X vssd1 vssd1 vccd1 vccd1 _8223_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold815 _7491_/Q vssd1 vssd1 vccd1 vccd1 hold815/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6252_ _6251_/A _5936_/Y _6251_/Y _6083_/A vssd1 vssd1 vccd1 vccd1 _6252_/X sky130_fd_sc_hd__a211o_1
Xhold848 _7024_/X vssd1 vssd1 vccd1 vccd1 _8482_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold859 _7440_/Q vssd1 vssd1 vccd1 vccd1 hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5203_ _4080_/X _5221_/A2 _5221_/B1 hold931/X vssd1 vssd1 vccd1 vccd1 _5203_/X sky130_fd_sc_hd__a22o_1
X_6183_ _3787_/B _6414_/B1 _6398_/B1 _6172_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6183_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5424__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5134_ _5134_/A1 _4448_/B _5140_/B1 _5133_/X vssd1 vssd1 vccd1 vccd1 _7379_/D sky130_fd_sc_hd__o211a_1
Xhold1515 _6784_/X vssd1 vssd1 vccd1 vccd1 _8329_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1526 _4157_/Y vssd1 vssd1 vccd1 vccd1 _4159_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1504 _7366_/Q vssd1 vssd1 vccd1 vccd1 _7044_/A sky130_fd_sc_hd__buf_2
Xhold1559 _4229_/Y vssd1 vssd1 vccd1 vccd1 _4230_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1537 _4197_/X vssd1 vssd1 vccd1 vccd1 _4198_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5065_ _5404_/A _5465_/C vssd1 vssd1 vccd1 vccd1 _5065_/X sky130_fd_sc_hd__or2_1
Xhold1548 _4308_/Y vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5273__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4016_ _4014_/A _4013_/Y _4014_/Y vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5967_ _5734_/A _5949_/X _5966_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _5967_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6773__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8466_/CLK sky130_fd_sc_hd__clkbuf_16
X_7706_ _8143_/CLK _7706_/D vssd1 vssd1 vccd1 vccd1 _7706_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5981__A0 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4918_ _4916_/X _4917_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4918_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7637_ _8365_/CLK _7637_/D vssd1 vssd1 vccd1 vccd1 _7637_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7086__B _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _5952_/A _5898_/B vssd1 vssd1 vccd1 vccd1 _5899_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4849_ _8176_/Q _8208_/Q _8272_/Q _7780_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4849_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7568_ _8160_/CLK _7568_/D vssd1 vssd1 vccd1 vccd1 _7568_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7499_ _8451_/CLK _7499_/D vssd1 vssd1 vccd1 vccd1 _7499_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6519_ _6539_/A _6519_/B vssd1 vssd1 vccd1 vccd1 _6519_/X sky130_fd_sc_hd__and2_1
XFILLER_0_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6828__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_99_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _8503_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4665__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6446__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5264__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4698__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5016__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6764__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6213__B2 _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8283_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__7277__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4870__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5509__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4622__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4575__S _7365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4689__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_62_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6870_ _7029_/A _6870_/A2 _6845_/B _6869_/X vssd1 vssd1 vccd1 vccd1 _6870_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6755__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6803__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5821_ _5820_/B _5820_/C _5820_/A vssd1 vssd1 vccd1 vccd1 _5822_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_9_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5752_ _5804_/A _5752_/B vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__and2_1
XANTENNA__4861__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5419__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_14_clk _7871_/CLK vssd1 vssd1 vccd1 vccd1 _8487_/CLK sky130_fd_sc_hd__clkbuf_16
X_4703_ _8159_/Q _7558_/Q _7430_/Q _7590_/Q _4734_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4703_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_127_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_77_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5683_ _6524_/A _5683_/B vssd1 vssd1 vccd1 vccd1 _5683_/X sky130_fd_sc_hd__and2_1
X_8471_ _8471_/CLK _8471_/D vssd1 vssd1 vccd1 vccd1 _8471_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4634_ _4632_/X _4633_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5715__A0 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7422_ _8218_/CLK _7422_/D vssd1 vssd1 vccd1 vccd1 _7422_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold612 _5598_/X vssd1 vssd1 vccd1 vccd1 _7782_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _8172_/Q _8204_/Q _8268_/Q _7776_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4565_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5191__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7353_ _7977_/CLK _7353_/D vssd1 vssd1 vccd1 vccd1 _7353_/Q sky130_fd_sc_hd__dfxtp_1
Xhold601 _8276_/Q vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold623 _7570_/Q vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 _6592_/X vssd1 vssd1 vccd1 vccd1 _8164_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ _6233_/X _6303_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6305_/B sky130_fd_sc_hd__mux2_1
Xhold645 _8162_/Q vssd1 vssd1 vccd1 vccd1 hold645/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold667 _7410_/Q vssd1 vssd1 vccd1 vccd1 hold667/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold656 _5600_/X vssd1 vssd1 vccd1 vccd1 _7784_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7284_ _8363_/CLK _7284_/D _6494_/A vssd1 vssd1 vccd1 vccd1 _7284_/Q sky130_fd_sc_hd__dfrtp_4
Xhold678 _5250_/X vssd1 vssd1 vccd1 vccd1 _7458_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4496_ _5160_/A1 _4496_/A1 _5465_/C vssd1 vssd1 vccd1 vccd1 _7302_/D sky130_fd_sc_hd__mux2_1
Xhold689 _7801_/Q vssd1 vssd1 vccd1 vccd1 hold689/X sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ _6411_/S _6235_/B vssd1 vssd1 vccd1 vccd1 _6235_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_15_clk_A _7871_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6166_ _5760_/Y _6130_/B _6159_/A _6414_/A2 _6165_/X vssd1 vssd1 vccd1 vccd1 _6166_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6691__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1312 _8391_/Q vssd1 vssd1 vccd1 vccd1 _6850_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1323 _6614_/X vssd1 vssd1 vccd1 vccd1 _8171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6097_ _6097_/A _6097_/B vssd1 vssd1 vccd1 vccd1 _6098_/B sky130_fd_sc_hd__nand2_1
Xhold1301 _6938_/X vssd1 vssd1 vccd1 vccd1 _8434_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4485__S _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1334 _8189_/Q vssd1 vssd1 vccd1 vccd1 _6650_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5117_ _7075_/A _5465_/C vssd1 vssd1 vccd1 vccd1 _5117_/X sky130_fd_sc_hd__or2_1
Xhold1345 _6810_/X vssd1 vssd1 vccd1 vccd1 _8342_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1356 _8448_/Q vssd1 vssd1 vccd1 vccd1 _6966_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1367 _7034_/Y vssd1 vssd1 vccd1 vccd1 _7035_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5246__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5048_ _4389_/A _5067_/S _5166_/B1 _5047_/X vssd1 vssd1 vccd1 vccd1 _7336_/D sky130_fd_sc_hd__o211a_1
Xhold1389 _8366_/Q vssd1 vssd1 vccd1 vccd1 _5020_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1378 _8386_/Q vssd1 vssd1 vccd1 vccd1 _5060_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6746__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6999_ _6999_/A _6999_/B vssd1 vssd1 vccd1 vccd1 _6999_/X sky130_fd_sc_hd__and2_1
Xclkbuf_4_8_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_8_0_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__7097__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5706__A0 _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4604__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3732__A2 _6445_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6357__S1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6682__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6607__C _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5237__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5511__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output118_A _7312_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6623__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6737__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4843__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ _4350_/A _4350_/B vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4281_ _4281_/A _4281_/B vssd1 vssd1 vccd1 vccd1 _4281_/X sky130_fd_sc_hd__xor2_1
XANTENNA__6673__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6020_ _5806_/B _6362_/C _6019_/X _5881_/C vssd1 vssd1 vccd1 vccd1 _6020_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_3_clk clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _8467_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5421__C _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7971_ _8519_/CLK _7971_/D vssd1 vssd1 vccd1 vccd1 _7971_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4531__S0 _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6922_ _7008_/A _6922_/A2 _6943_/B _6921_/X vssd1 vssd1 vccd1 vccd1 _6922_/X sky130_fd_sc_hd__a31o_1
X_6853_ _6853_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6853_/X sky130_fd_sc_hd__and2_1
XANTENNA__6728__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6284__S0 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5804_ _5804_/A _5804_/B vssd1 vssd1 vccd1 vccd1 _5926_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6784_ _6849_/A _6779_/B _6783_/X vssd1 vssd1 vccd1 vccd1 _6784_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_119_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3996_ _3996_/A _3996_/B vssd1 vssd1 vccd1 vccd1 _3996_/X sky130_fd_sc_hd__and2_1
XFILLER_0_85_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5735_ _3935_/B _6398_/A2 _6413_/B1 _5789_/S _6011_/A2 vssd1 vssd1 vccd1 vccd1 _5735_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout316_A _5186_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5666_ _6534_/A hold85/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__and2_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8454_ _8454_/CLK _8454_/D vssd1 vssd1 vccd1 vccd1 _8454_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7405_ _8136_/CLK _7405_/D vssd1 vssd1 vccd1 vccd1 _7405_/Q sky130_fd_sc_hd__dfxtp_1
X_4617_ _4616_/X _4613_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7513_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4598__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold420 _5244_/X vssd1 vssd1 vccd1 vccd1 _7452_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8385_ _8385_/CLK _8385_/D _7279_/Y vssd1 vssd1 vccd1 vccd1 _8385_/Q sky130_fd_sc_hd__dfrtp_1
X_5597_ _6931_/A _5616_/A2 _5616_/B1 hold765/X vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold431 _7814_/Q vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 _5358_/X vssd1 vssd1 vccd1 vccd1 _7585_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7336_ _8091_/CLK _7336_/D vssd1 vssd1 vccd1 vccd1 _7336_/Q sky130_fd_sc_hd__dfxtp_1
Xhold453 _7463_/Q vssd1 vssd1 vccd1 vccd1 hold453/X sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _8330_/Q _7806_/Q _7472_/Q _7440_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4548_/X sky130_fd_sc_hd__mux4_1
X_4479_ _7008_/A _7908_/Q vssd1 vssd1 vccd1 vccd1 _8040_/D sky130_fd_sc_hd__and2_1
Xhold464 _5302_/X vssd1 vssd1 vccd1 vccd1 _7533_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _6757_/X vssd1 vssd1 vccd1 vccd1 _8308_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _8218_/Q vssd1 vssd1 vccd1 vccd1 hold475/X sky130_fd_sc_hd__dlygate4sd3_1
X_7267_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7267_/Y sky130_fd_sc_hd__inv_2
Xhold497 _7823_/Q vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
X_6218_ _6342_/S _6066_/B _6214_/X _6217_/X vssd1 vssd1 vccd1 vccd1 _6218_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6664__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1131 _8428_/Q vssd1 vssd1 vccd1 vccd1 _6926_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1120 _6952_/X vssd1 vssd1 vccd1 vccd1 _8441_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _6828_/X vssd1 vssd1 vccd1 vccd1 _8351_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ _3800_/A _6414_/A2 _6130_/B _5719_/X _6148_/X vssd1 vssd1 vccd1 vccd1 _6149_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5219__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1153 _7783_/Q vssd1 vssd1 vccd1 vccd1 _5599_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 _8180_/Q vssd1 vssd1 vccd1 vccd1 _6632_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 _6866_/X vssd1 vssd1 vccd1 vccd1 _8399_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1186 _6932_/X vssd1 vssd1 vccd1 vccd1 _8431_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4943__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1197 _8415_/Q vssd1 vssd1 vccd1 vccd1 _6898_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6443__B _6443_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6719__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6195__A3 _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5059__B _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__S1 _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3953__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5075__A _5544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5506__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6104__B1 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5522__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4419__A _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4130__A2 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5630__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3850_ _7993_/Q _4068_/A2 _4068_/B1 _8025_/Q _3849_/X vssd1 vssd1 vccd1 vccd1 _3850_/X
+ sky130_fd_sc_hd__a221o_1
X_3781_ _4762_/B _4071_/A2 _4071_/B1 _6945_/A _3780_/X vssd1 vssd1 vccd1 vccd1 _6175_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_6_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6591__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5520_ _8239_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7709_/D sky130_fd_sc_hd__and3_1
XFILLER_0_41_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5451_ _5451_/A _7073_/A _5451_/C vssd1 vssd1 vccd1 vccd1 _5451_/X sky130_fd_sc_hd__and3_1
XFILLER_0_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5382_ _6977_/B _5382_/B vssd1 vssd1 vccd1 vccd1 _5382_/X sky130_fd_sc_hd__or2_1
XANTENNA__6894__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8170_ _8460_/CLK _8170_/D vssd1 vssd1 vccd1 vccd1 _8170_/Q sky130_fd_sc_hd__dfxtp_1
X_4402_ _5040_/A1 _5182_/A2 _4400_/X _4401_/Y vssd1 vssd1 vccd1 vccd1 _8376_/D sky130_fd_sc_hd__a22o_1
XANTENNA__6809__A _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4333_ _5576_/B _4382_/A _5470_/B vssd1 vssd1 vccd1 vccd1 _4383_/B sky130_fd_sc_hd__mux2_2
X_7121_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7121_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout229 _7073_/B vssd1 vssd1 vccd1 vccd1 _5546_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__6646__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout207 _3906_/X vssd1 vssd1 vccd1 vccd1 _6250_/S sky130_fd_sc_hd__clkbuf_4
X_7052_ _7052_/A _7079_/C vssd1 vssd1 vccd1 vccd1 _7052_/X sky130_fd_sc_hd__or2_1
Xfanout218 _5456_/C vssd1 vssd1 vccd1 vccd1 _5465_/C sky130_fd_sc_hd__buf_4
X_4264_ _8501_/Q _4264_/B vssd1 vssd1 vccd1 vccd1 _4264_/Y sky130_fd_sc_hd__nand2_1
X_6003_ _4044_/A _6398_/A2 _6413_/B1 _5990_/A _6011_/A2 vssd1 vssd1 vccd1 vccd1 _6005_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5854__C1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5432__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4195_ _8511_/Q _7636_/Q vssd1 vssd1 vccd1 vccd1 _4196_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3880__A1 _6444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5859__S _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6544__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7954_ _8090_/CLK hold40/X vssd1 vssd1 vccd1 vccd1 _7954_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5082__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3887__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6905_ _6971_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6905_/X sky130_fd_sc_hd__and2_1
X_7207__85 _8319_/CLK vssd1 vssd1 vccd1 vccd1 _8120_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7885_ _8270_/CLK _7885_/D vssd1 vssd1 vccd1 vccd1 _7885_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7078__C _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout433_A _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6836_ _7025_/A _6836_/A2 _6838_/A3 _6835_/X vssd1 vssd1 vccd1 vccd1 _6836_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_135_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6031__C1 _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6582__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4807__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6767_ _6891_/A _6773_/A2 _6773_/B1 hold939/X vssd1 vssd1 vccd1 vccd1 _6767_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_135_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8506_ _8513_/CLK _8506_/D vssd1 vssd1 vccd1 vccd1 _8506_/Q sky130_fd_sc_hd__dfxtp_1
X_5718_ _5714_/X _5874_/B _5950_/S vssd1 vssd1 vccd1 vccd1 _5718_/X sky130_fd_sc_hd__mux2_1
X_3979_ _4751_/B _3676_/A _4082_/B1 _3977_/X _3978_/X vssd1 vssd1 vccd1 vccd1 _5946_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_18_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6698_ _6963_/A _6701_/A2 _6701_/B1 hold971/X vssd1 vssd1 vccd1 vccd1 _6698_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_103_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8437_ _8473_/CLK _8437_/D vssd1 vssd1 vccd1 vccd1 _8437_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5649_ _6963_/A _5652_/A2 _5652_/B1 hold887/X vssd1 vssd1 vccd1 vccd1 _5649_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_32_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8368_ _8368_/CLK _8368_/D _7262_/Y vssd1 vssd1 vccd1 vccd1 _8368_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold261 _5588_/X vssd1 vssd1 vccd1 vccd1 _7772_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7319_ _8363_/CLK _7319_/D vssd1 vssd1 vccd1 vccd1 _7319_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold250 _7394_/Q vssd1 vssd1 vccd1 vccd1 _5461_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _7385_/Q vssd1 vssd1 vccd1 vccd1 _5452_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _7322_/Q vssd1 vssd1 vccd1 vccd1 _5419_/A sky130_fd_sc_hd__dlygate4sd3_1
X_8299_ _8425_/CLK _8299_/D vssd1 vssd1 vccd1 vccd1 _8299_/Q sky130_fd_sc_hd__dfxtp_1
Xhold283 _5441_/X vssd1 vssd1 vccd1 vccd1 _7630_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6454__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4673__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7062__A1 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5612__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6573__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3726__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6901__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3926__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4421__B _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6876__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4848__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6340__A3 _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6628__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4982__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4734__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 i_instr_ID[16] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
XFILLER_0_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3862__A1 _3861_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5064__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5603__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6800__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4951_ _8351_/Q _7827_/Q _7493_/Q _7461_/Q _4997_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4951_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7670_ _8328_/CLK _7670_/D vssd1 vssd1 vccd1 vccd1 _7670_/Q sky130_fd_sc_hd__dfxtp_1
X_3902_ hold5/X _3676_/A _4082_/B1 _6849_/A _3901_/X vssd1 vssd1 vccd1 vccd1 _5846_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_86_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4882_ _8148_/Q _7547_/Q _7419_/Q _7579_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4882_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_117_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6621_ _6927_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6621_/X sky130_fd_sc_hd__and2_1
X_3833_ _6367_/A vssd1 vssd1 vccd1 vccd1 _3833_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5367__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6811__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6552_ _6552_/A _6552_/B vssd1 vssd1 vccd1 vccd1 _8034_/D sky130_fd_sc_hd__and2_1
XANTENNA__3917__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3764_ _3764_/A _3764_/B vssd1 vssd1 vccd1 vccd1 _3800_/A sky130_fd_sc_hd__and2_1
XFILLER_0_55_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3695_ _7661_/Q _3653_/Y _3687_/Y _3689_/Y _7902_/Q vssd1 vssd1 vccd1 vccd1 _3696_/C
+ sky130_fd_sc_hd__o2111ai_1
X_6483_ _6524_/A hold33/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__and2_1
XFILLER_0_15_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5503_ _7524_/Q _5503_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _7692_/D sky130_fd_sc_hd__and3_1
XANTENNA__5427__B _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5434_ hold98/X _5465_/B _5463_/C vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__and3_1
X_8222_ _8460_/CLK _8222_/D vssd1 vssd1 vccd1 vccd1 _8222_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8153_ _8218_/CLK _8153_/D vssd1 vssd1 vccd1 vccd1 _8153_/Q sky130_fd_sc_hd__dfxtp_1
X_7104_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7104_/Y sky130_fd_sc_hd__inv_2
X_5365_ _6965_/A _5367_/A2 _5367_/B1 hold789/X vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4973__S0 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6539__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5296_ _5296_/A _7938_/Q _5183_/X vssd1 vssd1 vccd1 vccd1 _6842_/C sky130_fd_sc_hd__or3b_4
X_8084_ _8510_/CLK _8118_/D vssd1 vssd1 vccd1 vccd1 _8084_/Q sky130_fd_sc_hd__dfxtp_1
X_4316_ _4310_/A _4310_/B _4308_/B vssd1 vssd1 vccd1 vccd1 _4317_/B sky130_fd_sc_hd__o21a_1
XANTENNA_fanout383_A _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7035_ _7031_/Y _7035_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _7035_/Y sky130_fd_sc_hd__a21oi_1
X_4247_ _5564_/B _5030_/A1 _5503_/B vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__mux2_1
X_4178_ _4171_/Y _4178_/B vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__3853__B2 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7937_ _8080_/CLK _7937_/D vssd1 vssd1 vccd1 vccd1 _7937_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_96_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7868_ _8080_/CLK _7868_/D vssd1 vssd1 vccd1 vccd1 _7868_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold1498_A _7288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5358__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6819_ _6951_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6819_/X sky130_fd_sc_hd__and2_1
XFILLER_0_65_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6555__B1 _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7799_ _8350_/CLK _7799_/D vssd1 vssd1 vccd1 vccd1 _7799_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_135_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6858__A1 _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6322__A3 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6449__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6086__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4716__S0 _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5833__A2 _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5294__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5046__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5597__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4416__B _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output100_A _7295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7198__76 _8388_/CLK vssd1 vssd1 vccd1 vccd1 _8111_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6631__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6123__S _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5263__A _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4578__S _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4955__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5150_ _5150_/A1 _4416_/B _5166_/B1 _5149_/X vssd1 vssd1 vccd1 vccd1 _7387_/D sky130_fd_sc_hd__o211a_1
X_5081_ _5081_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__or2_1
X_4101_ _5892_/A _5889_/A vssd1 vssd1 vccd1 vccd1 _4101_/Y sky130_fd_sc_hd__nand2b_1
Xhold1708 _7694_/Q vssd1 vssd1 vccd1 vccd1 _3721_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4032_ _4032_/A _4032_/B vssd1 vssd1 vccd1 vccd1 _4109_/A sky130_fd_sc_hd__and2_1
Xhold1719 _7673_/Q vssd1 vssd1 vccd1 vccd1 _3992_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5285__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5588__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ _5879_/S _4095_/A _6028_/S vssd1 vssd1 vccd1 vccd1 _5983_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7722_ _8478_/CLK _7722_/D vssd1 vssd1 vccd1 vccd1 _7722_/Q sky130_fd_sc_hd__dfxtp_1
X_4934_ _8478_/Q _8410_/Q _8442_/Q _8316_/Q _4983_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4934_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4865_ _4864_/X _4863_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 _7597_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _6436_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7653_ _8091_/CLK _7653_/D vssd1 vssd1 vccd1 vccd1 _7653_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout229_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6604_ _6999_/A _6604_/A2 _6605_/B _6603_/X vssd1 vssd1 vccd1 vccd1 _6604_/X sky130_fd_sc_hd__a31o_1
X_4796_ _4795_/X _4792_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8232_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4012__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3816_ _3816_/A1 _4073_/A2 _6965_/A _4073_/B2 _3815_/X vssd1 vssd1 vccd1 vccd1 _3816_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_7_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7584_ _8471_/CLK _7584_/D vssd1 vssd1 vccd1 vccd1 _7584_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6535_ _6548_/A _6535_/B vssd1 vssd1 vccd1 vccd1 _8017_/D sky130_fd_sc_hd__and2_1
XANTENNA__5760__A1 _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3747_ _6334_/A _6331_/A vssd1 vssd1 vccd1 vccd1 _3749_/A sky130_fd_sc_hd__or2_1
XFILLER_0_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6466_ _6498_/A hold83/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__and2_1
X_3678_ _7282_/Q _3923_/B vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__or2_2
X_8205_ _8427_/CLK _8205_/D vssd1 vssd1 vccd1 vccd1 _8205_/Q sky130_fd_sc_hd__dfxtp_1
Xoutput141 _8057_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[22] sky130_fd_sc_hd__buf_12
Xoutput130 _8047_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[12] sky130_fd_sc_hd__buf_12
X_5417_ _5417_/A _7073_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5417_/X sky130_fd_sc_hd__and3_1
X_6397_ _6307_/A _6107_/Y _6128_/X vssd1 vssd1 vccd1 vccd1 _6397_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput152 _8038_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[3] sky130_fd_sc_hd__buf_12
X_8136_ _8136_/CLK _8136_/D vssd1 vssd1 vccd1 vccd1 _8136_/Q sky130_fd_sc_hd__dfxtp_1
X_5348_ _6931_/A _5367_/A2 _5367_/B1 hold557/X vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_694 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8067_ _8507_/CLK _8067_/D vssd1 vssd1 vccd1 vccd1 _8067_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5276__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7018_ _7018_/A _7018_/B vssd1 vssd1 vccd1 vccd1 _7018_/X sky130_fd_sc_hd__and2_1
X_5279_ _6939_/A _5294_/A2 _5294_/B1 hold629/X vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5620__B _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5028__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6240__A2 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5200__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5751__A1 _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5782__S _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5083__A _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4937__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6700__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5514__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout390 hold1641/X vssd1 vssd1 vccd1 vccd1 _4720_/S0 sky130_fd_sc_hd__buf_4
XANTENNA__3817__A1 _3816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5530__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6231__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6767__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6782__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4650_ _8474_/Q _8406_/Q _8438_/Q _8312_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4650_/X sky130_fd_sc_hd__mux4_1
Xinput21 i_instr_ID[2] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput10 i_instr_ID[19] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
X_4581_ _4580_/X _4579_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _4581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput32 i_read_data_M[10] vssd1 vssd1 vccd1 vccd1 _6531_/B sky130_fd_sc_hd__buf_1
X_6320_ _6320_/A _6320_/B vssd1 vssd1 vccd1 vccd1 _6320_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput43 i_read_data_M[20] vssd1 vssd1 vccd1 vccd1 _6541_/B sky130_fd_sc_hd__buf_1
XANTENNA__3753__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput54 i_read_data_M[30] vssd1 vssd1 vccd1 vccd1 _6551_/B sky130_fd_sc_hd__clkbuf_1
Xhold805 _7868_/Q vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__buf_1
Xhold827 _8472_/Q vssd1 vssd1 vccd1 vccd1 _7014_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold816 _5287_/X vssd1 vssd1 vccd1 vccd1 _7491_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold838 _6571_/X vssd1 vssd1 vccd1 vccd1 _8143_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6251_ _6251_/A _6251_/B vssd1 vssd1 vccd1 vccd1 _6251_/Y sky130_fd_sc_hd__nor2_1
Xhold849 _7426_/Q vssd1 vssd1 vccd1 vccd1 hold849/X sky130_fd_sc_hd__dlygate4sd3_1
X_5202_ _6933_/A _5221_/A2 _5221_/B1 hold669/X vssd1 vssd1 vccd1 vccd1 _5202_/X sky130_fd_sc_hd__a22o_1
X_6182_ _6126_/A _5881_/C _5792_/Y _5793_/Y vssd1 vssd1 vccd1 vccd1 _6182_/X sky130_fd_sc_hd__a22o_1
X_5133_ _5446_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5133_/X sky130_fd_sc_hd__or2_1
Xhold1516 hold1809/X vssd1 vssd1 vccd1 vccd1 _5545_/A sky130_fd_sc_hd__buf_1
Xhold1505 _7044_/Y vssd1 vssd1 vccd1 vccd1 _7045_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6817__A _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5258__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5064_ input21/X _4425_/B _5146_/B1 _5063_/X vssd1 vssd1 vccd1 vccd1 _7344_/D sky130_fd_sc_hd__o211a_1
Xhold1538 _4198_/X vssd1 vssd1 vccd1 vccd1 _5557_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 _4159_/Y vssd1 vssd1 vccd1 vccd1 _5552_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3808__A1 _3807_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1549 _4310_/X vssd1 vssd1 vccd1 vccd1 _5573_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4015_ _4014_/A _4013_/Y _4014_/Y vssd1 vssd1 vccd1 vccd1 _5971_/A sky130_fd_sc_hd__o21a_1
XANTENNA__5440__B _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A hold1510/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6758__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6552__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A _3966_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5966_ _5793_/Y _5962_/X _5965_/X _5694_/Y vssd1 vssd1 vccd1 vccd1 _5966_/X sky130_fd_sc_hd__a22o_1
X_7705_ _8473_/CLK _7705_/D vssd1 vssd1 vccd1 vccd1 _7705_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5981__A1 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5897_ _6270_/A _5897_/B vssd1 vssd1 vccd1 vccd1 _5900_/B sky130_fd_sc_hd__nor2_1
X_4917_ _8153_/Q _7552_/Q _7424_/Q _7584_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4917_/X sky130_fd_sc_hd__mux4_1
X_4848_ _4846_/X _4847_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3992__B1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7636_ _8364_/CLK _7636_/D vssd1 vssd1 vccd1 vccd1 _7636_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4779_ _8166_/Q _8198_/Q _8262_/Q _7770_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4779_/X sky130_fd_sc_hd__mux4_1
X_7567_ _8338_/CLK _7567_/D vssd1 vssd1 vccd1 vccd1 _7567_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6518_ _6524_/A _6518_/B vssd1 vssd1 vccd1 vccd1 _6518_/X sky130_fd_sc_hd__and2_1
X_7498_ _8467_/CLK _7498_/D vssd1 vssd1 vccd1 vccd1 _7498_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6289__A2 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4919__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6449_ _7028_/A _6449_/B vssd1 vssd1 vccd1 vccd1 _7931_/D sky130_fd_sc_hd__and2_1
XANTENNA__4011__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8119_ _8119_/CLK _8119_/D vssd1 vssd1 vccd1 vccd1 _8119_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5249__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4946__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6446__B _6446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6749__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6462__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7168__46 _8471_/CLK vssd1 vssd1 vccd1 vccd1 _8048_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5509__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3735__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5525__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7242__120 _8478_/CLK vssd1 vssd1 vccd1 vccd1 _8252_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_0_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6637__A _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6204__A2 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5820_ _5820_/A _5820_/B _5820_/C vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__and3_1
XFILLER_0_69_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5751_ _6388_/A _6370_/A _5772_/S vssd1 vssd1 vccd1 vccd1 _5752_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_84_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8470_ _8477_/CLK _8470_/D vssd1 vssd1 vccd1 vccd1 _8470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4702_ _8352_/Q _7828_/Q _7494_/Q _7462_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4702_/X sky130_fd_sc_hd__mux4_1
X_7421_ _8343_/CLK _7421_/D vssd1 vssd1 vccd1 vccd1 _7421_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5682_ _6551_/A hold79/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__and2_1
XFILLER_0_114_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4633_ _8149_/Q _7548_/Q _7420_/Q _7580_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4633_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5715__A1 _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7352_ _7907_/CLK _7352_/D vssd1 vssd1 vccd1 vccd1 _7352_/Q sky130_fd_sc_hd__dfxtp_1
X_4564_ _4562_/X _4563_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold602 _6721_/X vssd1 vssd1 vccd1 vccd1 _8276_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7182__60 _8010_/CLK vssd1 vssd1 vccd1 vccd1 _8062_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold624 _5343_/X vssd1 vssd1 vccd1 vccd1 _7570_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7283_ _8507_/CLK _7283_/D vssd1 vssd1 vccd1 vccd1 _7283_/Q sky130_fd_sc_hd__dfxtp_4
Xhold635 _8293_/Q vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
X_6303_ _6298_/A _6281_/A _6262_/A _6244_/A _5744_/S _5859_/S vssd1 vssd1 vccd1 vccd1
+ _6303_/X sky130_fd_sc_hd__mux4_1
Xhold613 _7830_/Q vssd1 vssd1 vccd1 vccd1 hold613/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5435__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold668 _5196_/X vssd1 vssd1 vccd1 vccd1 _7410_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6234_ _6160_/X _6233_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6235_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_69_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold657 _8316_/Q vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 _6590_/X vssd1 vssd1 vccd1 vccd1 _8162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 _7492_/Q vssd1 vssd1 vccd1 vccd1 hold679/X sky130_fd_sc_hd__dlygate4sd3_1
X_4495_ _5162_/A1 _4397_/B _5463_/C vssd1 vssd1 vccd1 vccd1 _7303_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6547__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6165_ _3775_/X _6414_/B1 _6398_/B1 _6154_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6165_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6691__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1313 _6850_/X vssd1 vssd1 vccd1 vccd1 _8391_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5116_ input19/X _5099_/B _5148_/B1 _5115_/X vssd1 vssd1 vccd1 vccd1 _7370_/D sky130_fd_sc_hd__o211a_1
X_6096_ _6096_/A _6096_/B vssd1 vssd1 vccd1 vccd1 _6097_/B sky130_fd_sc_hd__or2_1
Xhold1324 _8185_/Q vssd1 vssd1 vccd1 vccd1 _6642_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _8330_/Q vssd1 vssd1 vccd1 vccd1 _6786_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5877__S1 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1357 _6966_/X vssd1 vssd1 vccd1 vccd1 _8448_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1368 _7035_/Y vssd1 vssd1 vccd1 vccd1 _8490_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1335 _6650_/X vssd1 vssd1 vccd1 vccd1 _8189_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5047_ _5433_/A _5465_/C vssd1 vssd1 vccd1 vccd1 _5047_/X sky130_fd_sc_hd__or2_1
Xhold1346 _8355_/Q vssd1 vssd1 vccd1 vccd1 _6836_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1379 hold1800/X vssd1 vssd1 vccd1 vccd1 _5034_/A1 sky130_fd_sc_hd__buf_1
XANTENNA__5651__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout463_A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6998_ _6999_/A _6998_/B vssd1 vssd1 vccd1 vccd1 _6998_/X sky130_fd_sc_hd__and2_1
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5949_ _5949_/A _5949_/B vssd1 vssd1 vccd1 vccd1 _5949_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_48_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5706__A1 _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7619_ _8373_/CLK _7619_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
X_7226__104 _8175_/CLK vssd1 vssd1 vccd1 vccd1 _8236_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__5182__A2 _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6682__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4676__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5642__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3956__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4280_ _4270_/Y _4274_/B _4272_/B vssd1 vssd1 vccd1 vccd1 _4281_/B sky130_fd_sc_hd__o21a_1
X_7970_ _8363_/CLK _7970_/D vssd1 vssd1 vccd1 vccd1 _7970_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5633__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4531__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6921_ _6921_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6921_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6852_ _7024_/A _6852_/A2 _6906_/A3 _6851_/X vssd1 vssd1 vccd1 vccd1 _6852_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6284__S1 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5803_ _5952_/A _5803_/B vssd1 vssd1 vccd1 vccd1 _5803_/Y sky130_fd_sc_hd__nor2_1
X_6783_ _6911_/A _6783_/B _6839_/B vssd1 vssd1 vccd1 vccd1 _6783_/X sky130_fd_sc_hd__or3_1
X_3995_ _5892_/A _5889_/A vssd1 vssd1 vccd1 vccd1 _3996_/B sky130_fd_sc_hd__nand2_1
X_5734_ _5734_/A _6380_/A _5734_/C vssd1 vssd1 vccd1 vccd1 _5734_/X sky130_fd_sc_hd__and3_2
XFILLER_0_57_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5665_ _6498_/A _5665_/B vssd1 vssd1 vccd1 vccd1 _5665_/X sky130_fd_sc_hd__and2_1
X_8453_ _8515_/CLK _8453_/D vssd1 vssd1 vccd1 vccd1 _8453_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7404_ _8136_/CLK _7404_/D vssd1 vssd1 vccd1 vccd1 _7404_/Q sky130_fd_sc_hd__dfxtp_1
X_4616_ _4615_/X _4614_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4616_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8384_ _8387_/CLK _8384_/D _7278_/Y vssd1 vssd1 vccd1 vccd1 _8384_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5164__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5596_ _6929_/A _5584_/B _5617_/B1 hold785/X vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_115_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5795__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6900__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold410 _7561_/Q vssd1 vssd1 vccd1 vccd1 hold410/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7335_ _8379_/CLK _7335_/D vssd1 vssd1 vccd1 vccd1 _7335_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4598__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 _7803_/Q vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _4546_/X _4543_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7503_/D sky130_fd_sc_hd__mux2_1
Xhold432 _5634_/X vssd1 vssd1 vccd1 vccd1 _7814_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 _7540_/Q vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _5255_/X vssd1 vssd1 vccd1 vccd1 _7463_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _7008_/A _7909_/Q vssd1 vssd1 vccd1 vccd1 _8041_/D sky130_fd_sc_hd__and2_1
Xhold487 _7563_/Q vssd1 vssd1 vccd1 vccd1 hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 _7790_/Q vssd1 vssd1 vccd1 vccd1 hold465/X sky130_fd_sc_hd__dlygate4sd3_1
X_7266_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7266_/Y sky130_fd_sc_hd__inv_2
Xhold476 _6691_/X vssd1 vssd1 vccd1 vccd1 _8218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 _5643_/X vssd1 vssd1 vccd1 vccd1 _7823_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ _6302_/A _6309_/A _6217_/C vssd1 vssd1 vccd1 vccd1 _6217_/X sky130_fd_sc_hd__or3_1
XANTENNA__4496__S _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6148_ _3764_/A _6414_/B1 _6398_/B1 _6137_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6148_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 _8327_/Q vssd1 vssd1 vccd1 vccd1 _6780_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1132 _6926_/X vssd1 vssd1 vccd1 vccd1 _8428_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _6902_/X vssd1 vssd1 vccd1 vccd1 _8417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 _8394_/Q vssd1 vssd1 vccd1 vccd1 _6856_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5624__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1154 _5599_/X vssd1 vssd1 vccd1 vccd1 _7783_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6079_ _6016_/A _6035_/A _6056_/A _6075_/A _5782_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6079_/X sky130_fd_sc_hd__mux4_1
Xhold1176 _6632_/X vssd1 vssd1 vccd1 vccd1 _8180_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 _8404_/Q vssd1 vssd1 vccd1 vccd1 _6876_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 _8369_/Q vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1198 _6898_/X vssd1 vssd1 vccd1 vccd1 _8415_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1695_A _3958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7138__16 _8450_/CLK vssd1 vssd1 vccd1 vccd1 _7515_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_91_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5075__B _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_61_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5522__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__A _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4419__B _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6915__A _6915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5615__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6958__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6591__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3780_ _3780_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3780_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_14_clk_A _7871_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5450_ _5450_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__and3_1
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5146__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5777__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6343__B2 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4401_ _4401_/A _4407_/B vssd1 vssd1 vccd1 vccd1 _4401_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_29_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5381_ _7069_/A _5386_/B vssd1 vssd1 vccd1 vccd1 _5382_/B sky130_fd_sc_hd__nand2_1
X_7152__30 _8463_/CLK vssd1 vssd1 vccd1 vccd1 _7529_/CLK sky130_fd_sc_hd__inv_2
X_4332_ _4332_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__xor2_1
X_7120_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7120_/Y sky130_fd_sc_hd__inv_2
Xfanout208 _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6292_/A sky130_fd_sc_hd__buf_4
XANTENNA__6809__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7051_ _7031_/Y _7051_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8498_/D sky130_fd_sc_hd__a21oi_1
Xfanout219 _7073_/B vssd1 vssd1 vccd1 vccd1 _5456_/C sky130_fd_sc_hd__clkbuf_4
X_4263_ _4263_/A _4264_/B vssd1 vssd1 vccd1 vccd1 _4263_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5854__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6002_ _5694_/Y _6001_/X _6000_/X vssd1 vssd1 vccd1 vccd1 _6002_/X sky130_fd_sc_hd__a21bo_1
Xclkbuf_4_7_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_7_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_4194_ _8511_/Q _7636_/Q vssd1 vssd1 vccd1 vccd1 _4194_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5606__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6825__A _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4409__A1 _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7953_ _8034_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _7953_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6904_ _6434_/A _6904_/A2 _6906_/A3 _6903_/X vssd1 vssd1 vccd1 vccd1 _6904_/X sky130_fd_sc_hd__a31o_1
X_7884_ _8086_/CLK _7884_/D vssd1 vssd1 vccd1 vccd1 _7884_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout259_A _5299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout161_A _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4064__B _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6835_ _6967_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6835_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6560__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout426_A _7283_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6582__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3978_ _3978_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3978_/X sky130_fd_sc_hd__or2_1
X_6766_ _6955_/A _6773_/A2 _6773_/B1 hold599/X vssd1 vssd1 vccd1 vccd1 _6766_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8505_ _8513_/CLK _8505_/D vssd1 vssd1 vccd1 vccd1 _8505_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5717_ _5715_/X _5804_/B _5838_/A vssd1 vssd1 vccd1 vccd1 _5874_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6697_ _6961_/A _6701_/A2 _6701_/B1 hold571/X vssd1 vssd1 vccd1 vccd1 _6697_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8436_ _8472_/CLK _8436_/D vssd1 vssd1 vccd1 vccd1 _8436_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5648_ _6961_/A _5652_/A2 _5652_/B1 hold354/X vssd1 vssd1 vccd1 vccd1 _5648_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_130_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8367_ _8368_/CLK _8367_/D _7261_/Y vssd1 vssd1 vccd1 vccd1 _8367_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5579_ _6520_/A _5579_/B vssd1 vssd1 vccd1 vccd1 _7768_/D sky130_fd_sc_hd__and2_1
XFILLER_0_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold262 _8263_/Q vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold240 _7771_/Q vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
X_7318_ _7977_/CLK _7318_/D vssd1 vssd1 vccd1 vccd1 _7318_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8298_ _8460_/CLK _8298_/D vssd1 vssd1 vccd1 vccd1 _8298_/Q sky130_fd_sc_hd__dfxtp_1
Xhold251 _5461_/X vssd1 vssd1 vccd1 vccd1 _7650_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _7407_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 _5452_/X vssd1 vssd1 vccd1 vccd1 _7641_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _5419_/X vssd1 vssd1 vccd1 vccd1 _7608_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6248__S1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5517__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5128__A2 _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6325__B2 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6629__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4982__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5533__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4734__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 i_instr_ID[17] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6645__A _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _4949_/X _4946_/X _7057_/A vssd1 vssd1 vccd1 vccd1 _8254_/D sky130_fd_sc_hd__mux2_1
X_3901_ _7703_/Q _4081_/B vssd1 vssd1 vccd1 vccd1 _3901_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4881_ _8341_/Q _7817_/Q _7483_/Q _7451_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4881_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6564__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6620_ _4775_/A _6620_/A2 _6605_/B _6619_/X vssd1 vssd1 vccd1 vccd1 _6620_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6380__A _6380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3832_ _3968_/A _3830_/Y _3831_/Y vssd1 vssd1 vccd1 vccd1 _6367_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__5367__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6551_ _6551_/A _6551_/B vssd1 vssd1 vccd1 vccd1 _8033_/D sky130_fd_sc_hd__and2_1
XANTENNA__4670__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3763_ _6137_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3764_/B sky130_fd_sc_hd__nand2_1
X_5502_ _7523_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7691_/D sky130_fd_sc_hd__and3_1
XFILLER_0_27_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3694_ _3692_/Y _3693_/X _3690_/Y vssd1 vssd1 vccd1 vccd1 _3696_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6482_ _6524_/A hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5433_ _5433_/A _5465_/B _5465_/C vssd1 vssd1 vccd1 vccd1 _5433_/X sky130_fd_sc_hd__and3_1
X_8221_ _8353_/CLK _8221_/D vssd1 vssd1 vccd1 vccd1 _8221_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8152_ _8445_/CLK _8152_/D vssd1 vssd1 vccd1 vccd1 _8152_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5364_ _6963_/A _5367_/A2 _5367_/B1 hold813/X vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__a22o_1
X_7103_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7103_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5443__B _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4973__S1 _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4315_ _4315_/A _4315_/B vssd1 vssd1 vccd1 vccd1 _4315_/Y sky130_fd_sc_hd__nand2_1
X_5295_ _6971_/A _5262_/B _5295_/B1 hold861/X vssd1 vssd1 vccd1 vccd1 _5295_/X sky130_fd_sc_hd__a22o_1
X_8083_ _8086_/CLK _8117_/D vssd1 vssd1 vccd1 vccd1 _8083_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7034_ _7075_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7034_/Y sky130_fd_sc_hd__nand2_1
X_4246_ _4246_/A _4246_/B vssd1 vssd1 vccd1 vccd1 _4246_/X sky130_fd_sc_hd__xor2_1
X_4177_ _5554_/B _4442_/A _7082_/A vssd1 vssd1 vccd1 vccd1 _4178_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3853__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout376_A _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7936_ _8388_/CLK _7936_/D vssd1 vssd1 vccd1 vccd1 _7936_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4075__A _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7867_ _8500_/CLK _7867_/D vssd1 vssd1 vccd1 vccd1 _7867_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5358__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6818_ _6434_/A _6818_/A2 _6838_/A3 _6817_/X vssd1 vssd1 vccd1 vccd1 _6818_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_65_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7798_ _8319_/CLK _7798_/D vssd1 vssd1 vccd1 vccd1 _7798_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6749_ _6921_/A _6741_/B _6774_/B1 hold425/X vssd1 vssd1 vccd1 vccd1 _6749_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4661__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1658_A _3816_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8419_ _8419_/CLK _8419_/D vssd1 vssd1 vccd1 vccd1 _8419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4949__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4716__S1 _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6465__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5833__A3 _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5294__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6794__A1 _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5597__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5349__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4360__A1_N _7052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4859__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5544__A _5544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4955__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5080_ input1/X _5144_/A2 _5146_/B1 _5079_/X vssd1 vssd1 vccd1 vccd1 _7352_/D sky130_fd_sc_hd__o211a_1
X_4100_ _5921_/A _5918_/A vssd1 vssd1 vccd1 vccd1 _4100_/Y sky130_fd_sc_hd__nand2b_1
X_4031_ _6035_/A _6032_/A vssd1 vssd1 vccd1 vccd1 _4032_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5285__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1709 _8515_/Q vssd1 vssd1 vccd1 vccd1 _3968_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_37_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6094__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5982_ _5877_/X _5981_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _5982_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7721_ _8481_/CLK _7721_/D vssd1 vssd1 vccd1 vccd1 _7721_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4933_ _8188_/Q _8220_/Q _8284_/Q _7792_/Q _5089_/A _4969_/S1 vssd1 vssd1 vccd1 vccd1
+ _4933_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4891__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4864_ _8468_/Q _8400_/Q _8432_/Q _8306_/Q _4896_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4864_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_62_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 _7597_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7652_ _8382_/CLK _7652_/D vssd1 vssd1 vccd1 vccd1 _7652_/Q sky130_fd_sc_hd__dfxtp_1
X_4795_ _4794_/X _4793_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__mux2_1
X_6603_ _6777_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6603_/X sky130_fd_sc_hd__and2_1
XANTENNA__4012__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7583_ _8445_/CLK _7583_/D vssd1 vssd1 vccd1 vccd1 _7583_/Q sky130_fd_sc_hd__dfxtp_1
X_3815_ _4772_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3815_/X sky130_fd_sc_hd__and2_1
XANTENNA__5438__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_24 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6534_ _6534_/A _6534_/B vssd1 vssd1 vccd1 vccd1 _8016_/D sky130_fd_sc_hd__and2_1
XANTENNA__4643__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3746_ _3968_/A _6448_/B _3745_/Y vssd1 vssd1 vccd1 vccd1 _6331_/A sky130_fd_sc_hd__o21ai_2
X_6465_ _6498_/A _6465_/B vssd1 vssd1 vccd1 vccd1 _6465_/X sky130_fd_sc_hd__and2_1
XFILLER_0_70_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8204_ _8462_/CLK _8204_/D vssd1 vssd1 vccd1 vccd1 _8204_/Q sky130_fd_sc_hd__dfxtp_1
X_3677_ _7282_/Q _3923_/B vssd1 vssd1 vccd1 vccd1 _3677_/Y sky130_fd_sc_hd__nor2_1
X_5416_ _5416_/A _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5416_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput120 _7285_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[3] sky130_fd_sc_hd__buf_12
X_6396_ _6412_/S _6101_/X _6395_/X _5740_/B vssd1 vssd1 vccd1 vccd1 _6396_/X sky130_fd_sc_hd__o211a_1
XANTENNA__6170__C1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput142 _8058_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[23] sky130_fd_sc_hd__buf_12
Xoutput131 _8048_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[13] sky130_fd_sc_hd__buf_12
Xoutput153 _8039_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[4] sky130_fd_sc_hd__buf_12
X_8135_ _8136_/CLK _8135_/D vssd1 vssd1 vccd1 vccd1 _8135_/Q sky130_fd_sc_hd__dfxtp_1
X_5347_ _6929_/A _5335_/B _5368_/B1 hold899/X vssd1 vssd1 vccd1 vccd1 _5347_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5278_ _6937_/A _5262_/B _5295_/B1 hold923/X vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__a22o_1
X_8066_ _8066_/CLK _8066_/D vssd1 vssd1 vccd1 vccd1 _8066_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4079__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4229_ _8506_/Q _4229_/B vssd1 vssd1 vccd1 vccd1 _4229_/Y sky130_fd_sc_hd__nand2_1
X_7017_ _7017_/A _7017_/B vssd1 vssd1 vccd1 vccd1 _7017_/X sky130_fd_sc_hd__and2_1
XFILLER_0_97_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7919_ _8475_/CLK _7919_/D vssd1 vssd1 vccd1 vccd1 _7919_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5984__C1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4882__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5200__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4679__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4937__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6700__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5267__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout391 _7362_/Q vssd1 vssd1 vccd1 vccd1 _4727_/S0 sky130_fd_sc_hd__buf_8
Xfanout380 _7050_/A vssd1 vssd1 vccd1 vccd1 _4727_/S1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5530__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6923__A _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6767__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4580_ _8464_/Q _8396_/Q _8428_/Q _8302_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4580_/X sky130_fd_sc_hd__mux4_1
Xinput22 i_instr_ID[30] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_2
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput11 i_instr_ID[20] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_1
XANTENNA__4625__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput44 i_read_data_M[21] vssd1 vssd1 vccd1 vccd1 _6542_/B sky130_fd_sc_hd__clkbuf_1
Xinput33 i_read_data_M[11] vssd1 vssd1 vccd1 vccd1 _6532_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__4589__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput55 i_read_data_M[31] vssd1 vssd1 vccd1 vccd1 _6552_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold806 _8101_/D vssd1 vssd1 vccd1 vccd1 _8067_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _7014_/X vssd1 vssd1 vccd1 vccd1 _8472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 _8301_/Q vssd1 vssd1 vccd1 vccd1 hold817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7904__D _7904_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6250_ _6100_/X _6249_/X _6250_/S vssd1 vssd1 vccd1 vccd1 _6251_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_40_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold839 _8216_/Q vssd1 vssd1 vccd1 vccd1 hold839/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6181_ _5740_/B _6180_/X _5811_/X vssd1 vssd1 vccd1 vccd1 _6181_/Y sky130_fd_sc_hd__a21boi_1
X_5201_ _6931_/A _5188_/B _5220_/B1 hold621/X vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__a22o_1
X_5132_ _5132_/A1 _4448_/B _5140_/B1 _5131_/X vssd1 vssd1 vccd1 vccd1 _7378_/D sky130_fd_sc_hd__o211a_1
Xhold1517 _8358_/Q vssd1 vssd1 vccd1 vccd1 _5003_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1506 _7597_/Q vssd1 vssd1 vccd1 vccd1 hold1506/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6817__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5258__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5063_ _5404_/B _5451_/C vssd1 vssd1 vccd1 vccd1 _5063_/X sky130_fd_sc_hd__or2_1
Xhold1528 hold1797/X vssd1 vssd1 vccd1 vccd1 _4752_/B sky130_fd_sc_hd__clkbuf_2
Xhold1539 _4200_/B vssd1 vssd1 vccd1 vccd1 _4508_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_4014_ _4014_/A _4014_/B vssd1 vssd1 vccd1 vccd1 _4014_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5440__C _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6833__A _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6758__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4864__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5965_ _5963_/X _5964_/X _6028_/S vssd1 vssd1 vccd1 vccd1 _5965_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout241_A _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5981__A2 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5896_ _5746_/X _5750_/B _5950_/S vssd1 vssd1 vccd1 vccd1 _5897_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4916_ _8346_/Q _7822_/Q _7488_/Q _7456_/Q _5089_/A _4990_/S1 vssd1 vssd1 vccd1 vccd1
+ _4916_/X sky130_fd_sc_hd__mux4_1
X_7704_ _8195_/CLK _7704_/D vssd1 vssd1 vccd1 vccd1 _7704_/Q sky130_fd_sc_hd__dfxtp_1
X_4847_ _8143_/Q _7542_/Q _7414_/Q _7574_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4847_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3992__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7635_ _8358_/CLK _7635_/D vssd1 vssd1 vccd1 vccd1 _7635_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4072__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5194__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6930__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4778_ _4776_/X _4777_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__mux2_1
X_7566_ _8136_/CLK _7566_/D vssd1 vssd1 vccd1 vccd1 _7566_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3744__A1 _4771_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6517_ _6520_/A hold87/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__and2_1
XFILLER_0_43_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3729_ _3729_/A1 _4073_/A2 _6891_/A _4073_/B2 vssd1 vssd1 vccd1 vccd1 _3729_/X sky130_fd_sc_hd__a22o_1
X_7497_ _8355_/CLK _7497_/D vssd1 vssd1 vccd1 vccd1 _7497_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4919__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6448_ _7267_/A _6448_/B vssd1 vssd1 vccd1 vccd1 _7930_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_30_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6379_ _3836_/A _6414_/B1 _6398_/B1 _6367_/A _6292_/A vssd1 vssd1 vccd1 vccd1 _6379_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6694__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8118_ _8118_/CLK _8118_/D vssd1 vssd1 vccd1 vccd1 _8118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5249__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6997__A1 _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8049_ _8049_/CLK _8049_/D vssd1 vssd1 vccd1 vccd1 _8049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6749__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6213__A3 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4607__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3735__B2 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5525__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_100_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _8463_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6685__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6637__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5541__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4872__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6653__A _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4846__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5750_ _5950_/S _5750_/B vssd1 vssd1 vccd1 vccd1 _5750_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4701_ _4700_/X _4697_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7525_/D sky130_fd_sc_hd__mux2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _6524_/A _5681_/B vssd1 vssd1 vccd1 vccd1 _5681_/X sky130_fd_sc_hd__and2_1
XFILLER_0_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7420_ _8402_/CLK _7420_/D vssd1 vssd1 vccd1 vccd1 _7420_/Q sky130_fd_sc_hd__dfxtp_1
X_4632_ _8342_/Q _7818_/Q _7484_/Q _7452_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4632_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5176__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6912__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7351_ _8456_/CLK _7351_/D vssd1 vssd1 vccd1 vccd1 _7351_/Q sky130_fd_sc_hd__dfxtp_1
X_4563_ _8139_/Q _7538_/Q _7410_/Q _7570_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4563_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_8_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold603 _7428_/Q vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
X_7282_ _8507_/CLK _7282_/D vssd1 vssd1 vccd1 vccd1 _7282_/Q sky130_fd_sc_hd__dfxtp_2
Xhold636 _6738_/X vssd1 vssd1 vccd1 vccd1 _8293_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6302_ _6302_/A _6302_/B vssd1 vssd1 vccd1 vccd1 _6302_/Y sky130_fd_sc_hd__nand2_1
Xhold614 _5650_/X vssd1 vssd1 vccd1 vccd1 _7830_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold625 _8280_/Q vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _5164_/A1 _4395_/B _5462_/C vssd1 vssd1 vccd1 vccd1 _7304_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6676__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold669 _7416_/Q vssd1 vssd1 vccd1 vccd1 hold669/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold647 _8133_/Q vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap355 _6406_/B vssd1 vssd1 vccd1 vccd1 _5971_/B sky130_fd_sc_hd__buf_4
X_6233_ _6175_/A _6191_/A _6209_/A _6226_/A _5782_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6233_/X sky130_fd_sc_hd__mux4_1
Xhold658 _6765_/X vssd1 vssd1 vccd1 vccd1 _8316_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6164_ _6163_/A _6162_/X _6163_/Y _5740_/B vssd1 vssd1 vccd1 vccd1 _6164_/X sky130_fd_sc_hd__o211a_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__B _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A _5716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5115_ _7076_/A _5542_/C vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__or2_1
X_6095_ _6096_/A _6096_/B vssd1 vssd1 vccd1 vccd1 _6097_/A sky130_fd_sc_hd__nand2_1
Xhold1325 _6642_/X vssd1 vssd1 vccd1 vccd1 _8185_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1314 _8447_/Q vssd1 vssd1 vccd1 vccd1 _6964_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1303 _6786_/X vssd1 vssd1 vccd1 vccd1 _8330_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1358 _8331_/Q vssd1 vssd1 vccd1 vccd1 _6788_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5100__B1 _5002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_A _6703_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4067__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5046_ _5046_/A1 _4416_/B _5166_/B1 _5045_/X vssd1 vssd1 vccd1 vccd1 _7335_/D sky130_fd_sc_hd__o211a_1
Xhold1336 _8184_/Q vssd1 vssd1 vccd1 vccd1 _6640_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1347 _6836_/X vssd1 vssd1 vccd1 vccd1 _8355_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4782__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5878__S _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1369 _8439_/Q vssd1 vssd1 vccd1 vccd1 _6948_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5651__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout456_A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6997_ _7074_/A _6990_/S _6996_/Y _7079_/B vssd1 vssd1 vccd1 vccd1 _8455_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4083__A _4757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5948_ _5923_/A _5922_/A _5920_/Y vssd1 vssd1 vccd1 vccd1 _5949_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5879_ _5696_/X _5699_/X _5879_/S vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7618_ _8020_/CLK _7618_/D vssd1 vssd1 vccd1 vccd1 _7618_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7549_ _8339_/CLK _7549_/D vssd1 vssd1 vccd1 vccd1 _7549_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4957__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5642__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4828__S0 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5089__A _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3956__B2 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6412__S _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5158__B1 _5002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5536__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5552__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6367__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5330__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4436__A2 _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__S _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5633__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6920_ _6853_/A _6963_/B _6919_/X _7015_/A vssd1 vssd1 vccd1 vccd1 _6920_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6851_ _6917_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6851_/X sky130_fd_sc_hd__and2_1
XANTENNA__4819__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5802_ _5713_/X _5715_/X _5838_/A vssd1 vssd1 vccd1 vccd1 _5803_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6782_ _6706_/A _6782_/A2 _6779_/B _6781_/X vssd1 vssd1 vccd1 vccd1 _6782_/X sky130_fd_sc_hd__a31o_1
X_3994_ _5892_/A _5889_/A vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__or2_1
XFILLER_0_71_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5733_ _6413_/B1 _5786_/B _5733_/C _5733_/D vssd1 vssd1 vccd1 vccd1 _5734_/C sky130_fd_sc_hd__and4b_1
X_7249__127 _8463_/CLK vssd1 vssd1 vccd1 vccd1 _8259_/CLK sky130_fd_sc_hd__inv_2
X_8452_ _8507_/CLK _8452_/D vssd1 vssd1 vccd1 vccd1 _8452_/Q sky130_fd_sc_hd__dfxtp_1
X_5664_ _6498_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5664_/X sky130_fd_sc_hd__and2_1
XFILLER_0_60_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5595_ _6927_/A _5584_/B _5617_/B1 hold513/X vssd1 vssd1 vccd1 vccd1 _5595_/X sky130_fd_sc_hd__a22o_1
X_4615_ _8469_/Q _8401_/Q _8433_/Q _8307_/Q _4741_/S0 _4737_/S1 vssd1 vssd1 vccd1
+ vccd1 _4615_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5446__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7403_ _8360_/CLK _7403_/D vssd1 vssd1 vccd1 vccd1 _7403_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8383_ _8385_/CLK _8383_/D _7277_/Y vssd1 vssd1 vccd1 vccd1 _8383_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4546_ _4545_/X _4544_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4546_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold411 _5330_/X vssd1 vssd1 vccd1 vccd1 _7561_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7334_ _8379_/CLK _7334_/D vssd1 vssd1 vccd1 vccd1 _7334_/Q sky130_fd_sc_hd__dfxtp_1
Xhold400 _7820_/Q vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold444 _5623_/X vssd1 vssd1 vccd1 vccd1 _7803_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _5309_/X vssd1 vssd1 vccd1 vccd1 _7540_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold433 _8298_/Q vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold477 _8319_/Q vssd1 vssd1 vccd1 vccd1 hold477/X sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _6545_/A _7910_/Q vssd1 vssd1 vccd1 vccd1 _8042_/D sky130_fd_sc_hd__and2_1
Xhold466 _5606_/X vssd1 vssd1 vccd1 vccd1 _7790_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7265_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7265_/Y sky130_fd_sc_hd__inv_2
Xhold455 _8160_/Q vssd1 vssd1 vccd1 vccd1 hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 _5332_/X vssd1 vssd1 vccd1 vccd1 _7563_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6216_ _6143_/X _6215_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6217_/C sky130_fd_sc_hd__mux2_1
Xhold499 _7391_/Q vssd1 vssd1 vccd1 vccd1 _5458_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5321__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6664__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1100 _6910_/X vssd1 vssd1 vccd1 vccd1 _8420_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6147_ _6163_/A _6145_/X _6146_/X _5740_/B vssd1 vssd1 vccd1 vccd1 _6147_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5181__B _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _6780_/X vssd1 vssd1 vccd1 vccd1 _8327_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1111 _7598_/Q vssd1 vssd1 vccd1 vccd1 _6419_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1133 _8413_/Q vssd1 vssd1 vccd1 vccd1 _6894_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1155 _8389_/Q vssd1 vssd1 vccd1 vccd1 _6846_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 _6856_/X vssd1 vssd1 vccd1 vccd1 _8394_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5624__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6078_ _6078_/A _6078_/B vssd1 vssd1 vccd1 vccd1 _6078_/X sky130_fd_sc_hd__xor2_1
Xhold1144 _6876_/X vssd1 vssd1 vccd1 vccd1 _8404_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 _8400_/Q vssd1 vssd1 vccd1 vccd1 _6868_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 _5026_/X vssd1 vssd1 vccd1 vccd1 _7325_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1177 _8182_/Q vssd1 vssd1 vccd1 vccd1 _6636_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5029_ _5424_/A _5454_/C vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__or2_1
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold1688_A _3709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4060__A0 _4221_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3856__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6468__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5372__A _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4687__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5312__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5863__A1 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__B _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3874__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6915__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5615__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output123_A _7288_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6931__A _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6591__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5547__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4400_ _4410_/A _4406_/B _4404_/B _4496_/A1 vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5380_ _7065_/A _5395_/A vssd1 vssd1 vccd1 vccd1 _5386_/B sky130_fd_sc_hd__and2b_1
XANTENNA__6894__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4331_ _4325_/A _4322_/Y _4323_/Y vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__o21a_1
XANTENNA__6646__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout209 _5734_/X vssd1 vssd1 vccd1 vccd1 _6417_/A2 sky130_fd_sc_hd__clkbuf_8
X_7050_ _7050_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7050_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4262_ _4416_/A _4413_/B _4262_/C vssd1 vssd1 vccd1 vccd1 _4410_/A sky130_fd_sc_hd__and3_1
X_6001_ _5748_/B _5784_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6001_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_66_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4193_ _4440_/A _4193_/B _4193_/C vssd1 vssd1 vccd1 vccd1 _4435_/B sky130_fd_sc_hd__or3_1
XANTENNA__7056__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6825__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5606__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7952_ _8034_/CLK _7952_/D vssd1 vssd1 vccd1 vccd1 _7952_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5082__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7002__A _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6903_ _6969_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6903_/X sky130_fd_sc_hd__and2_1
XFILLER_0_77_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7883_ _8419_/CLK _7883_/D vssd1 vssd1 vccd1 vccd1 _7883_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6834_ _7026_/A _6834_/A2 _6838_/A3 _6833_/X vssd1 vssd1 vccd1 vccd1 _6834_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_92_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6582__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3977_ _8074_/Q _3976_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6765_ _6953_/A _6773_/A2 _6773_/B1 hold657/X vssd1 vssd1 vccd1 vccd1 _6765_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_134_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout321_A _4035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5716_ _6388_/A _6126_/A _5716_/S vssd1 vssd1 vccd1 vccd1 _5804_/B sky130_fd_sc_hd__mux2_1
X_8504_ _8504_/CLK _8504_/D vssd1 vssd1 vccd1 vccd1 _8504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6696_ _6959_/A _6701_/A2 _6701_/B1 hold803/X vssd1 vssd1 vccd1 vccd1 _6696_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout419_A hold1747/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8435_ _8471_/CLK _8435_/D vssd1 vssd1 vccd1 vccd1 _8435_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5647_ _6959_/A _5620_/B _5653_/B1 hold396/X vssd1 vssd1 vccd1 vccd1 _5647_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8366_ _8369_/CLK _8366_/D _7260_/Y vssd1 vssd1 vccd1 vccd1 _8366_/Q sky130_fd_sc_hd__dfrtp_1
X_5578_ _6539_/A _5578_/B vssd1 vssd1 vccd1 vccd1 _7767_/D sky130_fd_sc_hd__and2_1
Xhold241 _5587_/X vssd1 vssd1 vccd1 vccd1 _7771_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _8200_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
X_8297_ _8338_/CLK _8297_/D vssd1 vssd1 vccd1 vccd1 _8297_/Q sky130_fd_sc_hd__dfxtp_1
Xhold230 _7471_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4527_/X _4528_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _4529_/X sky130_fd_sc_hd__mux2_1
X_7317_ _8360_/CLK _7317_/D vssd1 vssd1 vccd1 vccd1 _7317_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold263 _6708_/X vssd1 vssd1 vccd1 vccd1 _8263_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _8198_/Q vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 _5193_/X vssd1 vssd1 vccd1 vccd1 _7407_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold296 _7336_/Q vssd1 vssd1 vccd1 vccd1 _5433_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5920__A _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7047__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4970__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_80_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _8096_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6573__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6022__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5781__A0 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4271__A _8500_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6876__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6628__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5533__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6645__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 i_instr_ID[18] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__5064__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5695__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6800__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3900_ _8070_/Q _3899_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _6915_/A sky130_fd_sc_hd__mux2_2
X_4880_ _4879_/X _4876_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8244_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4880__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_71_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _8358_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6661__A _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3831_ _3968_/A _3831_/B vssd1 vssd1 vccd1 vccd1 _3831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3762_ _6137_/A _6140_/A vssd1 vssd1 vccd1 vccd1 _3764_/A sky130_fd_sc_hd__or2_1
X_6550_ _6550_/A _6550_/B vssd1 vssd1 vccd1 vccd1 _8032_/D sky130_fd_sc_hd__and2_1
XFILLER_0_6_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7212__90 _8091_/CLK vssd1 vssd1 vccd1 vccd1 _8125_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4670__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5501_ _7522_/Q _5541_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7690_/D sky130_fd_sc_hd__and3_1
XFILLER_0_6_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3693_ _7663_/Q _7837_/Q vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__or2_1
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6481_ _6550_/A hold31/X vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__and2_1
XFILLER_0_70_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8220_ _8442_/CLK _8220_/D vssd1 vssd1 vccd1 vccd1 _8220_/Q sky130_fd_sc_hd__dfxtp_1
X_5432_ _5432_/A _5503_/B _5462_/C vssd1 vssd1 vccd1 vccd1 _5432_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8151_ _8450_/CLK _8151_/D vssd1 vssd1 vccd1 vccd1 _8151_/Q sky130_fd_sc_hd__dfxtp_1
X_5363_ _6961_/A _5367_/A2 _5367_/B1 hold559/X vssd1 vssd1 vccd1 vccd1 _5363_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7102_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7102_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5443__C _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4314_ _8494_/Q _4314_/B vssd1 vssd1 vccd1 vccd1 _4314_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5827__A1 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8082_ _8484_/CLK _8116_/D vssd1 vssd1 vccd1 vccd1 _8082_/Q sky130_fd_sc_hd__dfxtp_1
X_5294_ _6969_/A _5294_/A2 _5294_/B1 hold519/X vssd1 vssd1 vccd1 vccd1 _5294_/X sky130_fd_sc_hd__a22o_1
X_4245_ _4235_/Y _4238_/X _4237_/B vssd1 vssd1 vccd1 vccd1 _4246_/B sky130_fd_sc_hd__o21a_2
X_7033_ _7031_/Y _7033_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _7033_/Y sky130_fd_sc_hd__a21oi_1
X_4176_ _4176_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _4176_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_93_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout271_A _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A _7083_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6252__A1 _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7935_ _8010_/CLK _7935_/D vssd1 vssd1 vccd1 vccd1 _7935_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_60_clk_A clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _8369_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6004__A1 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7866_ _8030_/CLK _7866_/D vssd1 vssd1 vccd1 vccd1 _7866_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6004__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6817_ _6949_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6817_/X sky130_fd_sc_hd__and2_1
XFILLER_0_133_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7797_ _8483_/CLK _7797_/D vssd1 vssd1 vccd1 vccd1 _7797_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6748_ _6853_/A _6741_/B _6774_/B1 hold663/X vssd1 vssd1 vccd1 vccd1 _6748_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_116_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6679_ _6925_/A _6669_/B _6702_/B1 hold366/X vssd1 vssd1 vccd1 vccd1 _6679_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_75_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4661__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6858__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8418_ _8450_/CLK _8418_/D vssd1 vssd1 vccd1 vccd1 _8418_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8349_ _8353_/CLK _8349_/D vssd1 vssd1 vccd1 vccd1 _8349_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3829__B1 _3826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5294__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5046__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_53_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8456_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_28_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6481__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5528__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_6_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_6_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5544__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5560__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4030_ _6035_/A _6032_/A vssd1 vssd1 vccd1 vccd1 _4032_/A sky130_fd_sc_hd__or2_1
XANTENNA__5285__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5981_ _5921_/A _5892_/A _5974_/A _5946_/A _5716_/S _5804_/A vssd1 vssd1 vccd1 vccd1
+ _5981_/X sky130_fd_sc_hd__mux4_1
Xclkbuf_leaf_44_clk _7871_/CLK vssd1 vssd1 vccd1 vccd1 _8270_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6391__A _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4932_ _4930_/X _4931_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4932_/X sky130_fd_sc_hd__mux2_1
X_7720_ _8450_/CLK _7720_/D vssd1 vssd1 vccd1 vccd1 _7720_/Q sky130_fd_sc_hd__dfxtp_1
X_7189__67 _8519_/CLK vssd1 vssd1 vccd1 vccd1 _8102_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_86_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4891__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7651_ _8379_/CLK _7651_/D vssd1 vssd1 vccd1 vccd1 _7651_/Q sky130_fd_sc_hd__dfxtp_1
X_4863_ _8178_/Q _8210_/Q _8274_/Q _7782_/Q _4896_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4863_/X sky130_fd_sc_hd__mux4_1
X_6602_ _6704_/B _6776_/B vssd1 vssd1 vccd1 vccd1 _6602_/X sky130_fd_sc_hd__or2_2
XFILLER_0_74_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5745__A0 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 _7597_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4794_ _8458_/Q _8390_/Q _8422_/Q _8296_/Q _5475_/A _4867_/S1 vssd1 vssd1 vccd1 vccd1
+ _4794_/X sky130_fd_sc_hd__mux4_1
X_3814_ _8095_/Q _3813_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3814_/X sky130_fd_sc_hd__mux2_2
XANTENNA__5438__C _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7582_ _8218_/CLK _7582_/D vssd1 vssd1 vccd1 vccd1 _7582_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_25 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3954__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6533_ _6548_/A _6533_/B vssd1 vssd1 vccd1 vccd1 _8015_/D sky130_fd_sc_hd__and2_1
XANTENNA__4643__S1 _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3745_ _3968_/A _3745_/B vssd1 vssd1 vccd1 vccd1 _3745_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6464_ _6494_/A hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__and2_1
X_3676_ _3676_/A _3676_/B vssd1 vssd1 vccd1 vccd1 _3676_/Y sky130_fd_sc_hd__nand2_2
X_8203_ _8283_/CLK _8203_/D vssd1 vssd1 vccd1 vccd1 _8203_/Q sky130_fd_sc_hd__dfxtp_1
X_5415_ _5415_/A _7073_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5415_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput110 _7305_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[23] sky130_fd_sc_hd__buf_12
XANTENNA__5454__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput143 _8059_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[24] sky130_fd_sc_hd__buf_12
XFILLER_0_113_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6395_ _6270_/A _6249_/X _6393_/X _6394_/X _6309_/A vssd1 vssd1 vccd1 vccd1 _6395_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput132 _8049_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[14] sky130_fd_sc_hd__buf_12
XFILLER_0_2_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput121 _7286_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[4] sky130_fd_sc_hd__buf_12
XFILLER_0_11_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput154 _8040_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[5] sky130_fd_sc_hd__buf_12
X_8134_ _8428_/CLK _8134_/D vssd1 vssd1 vccd1 vccd1 _8134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5346_ _6927_/A _5335_/B _5368_/B1 hold415/X vssd1 vssd1 vccd1 vccd1 _5346_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4785__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5277_ _6935_/A _5262_/B _5295_/B1 hold979/X vssd1 vssd1 vccd1 vccd1 _5277_/X sky130_fd_sc_hd__a22o_1
X_8065_ _8065_/CLK _8065_/D vssd1 vssd1 vccd1 vccd1 _8065_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5276__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4228_ _8506_/Q _4229_/B vssd1 vssd1 vccd1 vccd1 _4228_/Y sky130_fd_sc_hd__nor2_1
X_7016_ _7028_/A _7016_/B vssd1 vssd1 vccd1 vccd1 _7016_/X sky130_fd_sc_hd__and2_1
XFILLER_0_128_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5028__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4159_ _4159_/A _4159_/B vssd1 vssd1 vccd1 vccd1 _4159_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7918_ _8440_/CLK _7918_/D vssd1 vssd1 vccd1 vccd1 _7918_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_35_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _8338_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4882__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7849_ _8034_/CLK _7849_/D vssd1 vssd1 vccd1 vccd1 _7849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5200__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5831__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6700__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6476__A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout381 _4737_/S1 vssd1 vssd1 vccd1 vccd1 _4740_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout392 _7072_/B2 vssd1 vssd1 vccd1 vccd1 _4696_/S0 sky130_fd_sc_hd__buf_8
Xfanout370 _7048_/A vssd1 vssd1 vccd1 vccd1 _5103_/A sky130_fd_sc_hd__buf_8
XANTENNA__4570__S0 _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6923__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6767__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8343_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__7100__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5539__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput12 i_instr_ID[21] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__4625__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput23 i_instr_ID[31] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_2
Xinput34 i_read_data_M[12] vssd1 vssd1 vccd1 vccd1 _6533_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__5555__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput45 i_read_data_M[22] vssd1 vssd1 vccd1 vccd1 _6543_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__3753__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold807 _7581_/Q vssd1 vssd1 vccd1 vccd1 hold807/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput56 i_read_data_M[3] vssd1 vssd1 vccd1 vccd1 _6524_/B sky130_fd_sc_hd__clkbuf_1
Xhold818 _6750_/X vssd1 vssd1 vccd1 vccd1 _8301_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold829 _7818_/Q vssd1 vssd1 vccd1 vccd1 hold829/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6152__B1 _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5200_ _6929_/A _5221_/A2 _5221_/B1 hold857/X vssd1 vssd1 vccd1 vccd1 _5200_/X sky130_fd_sc_hd__a22o_1
X_6180_ _6026_/B _6179_/X _6411_/S vssd1 vssd1 vccd1 vccd1 _6180_/X sky130_fd_sc_hd__mux2_1
X_5131_ _5445_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5131_/X sky130_fd_sc_hd__or2_1
Xhold1507 _6455_/X vssd1 vssd1 vccd1 vccd1 _7937_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5062_ _5062_/A1 _5182_/A2 _5182_/B1 _5061_/X vssd1 vssd1 vccd1 vccd1 _7343_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5258__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1518 _8421_/Q vssd1 vssd1 vccd1 vccd1 _6911_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1529 _8388_/Q vssd1 vssd1 vccd1 vccd1 _6843_/B sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ _4752_/B _3966_/B _4012_/X vssd1 vssd1 vccd1 vccd1 _4013_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_35_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6833__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6758__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7010__A _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5449__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7703_ _8328_/CLK _7703_/D vssd1 vssd1 vccd1 vccd1 _7703_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_17_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8473_/CLK sky130_fd_sc_hd__clkbuf_16
X_5964_ _5830_/X _5860_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _5964_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4864__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5895_ _5895_/A _5895_/B vssd1 vssd1 vccd1 vccd1 _5895_/X sky130_fd_sc_hd__xor2_1
XANTENNA__5981__A3 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4915_ _4914_/X _4911_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8249_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4846_ _8336_/Q _7812_/Q _7478_/Q _7446_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4846_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3992__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7634_ _8362_/CLK _7634_/D vssd1 vssd1 vccd1 vccd1 _7634_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout234_A _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7565_ _7805_/CLK _7565_/D vssd1 vssd1 vccd1 vccd1 _7565_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5194__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4777_ _8133_/Q _7532_/Q _7404_/Q _7564_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4777_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout401_A _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6516_ _6524_/A _6516_/B vssd1 vssd1 vccd1 vccd1 _6516_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3744__A2 _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7496_ _8354_/CLK _7496_/D vssd1 vssd1 vccd1 vccd1 _7496_/Q sky130_fd_sc_hd__dfxtp_1
X_3728_ _8091_/Q _3727_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _6957_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3659_ _7664_/Q vssd1 vssd1 vccd1 vccd1 _3659_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_113_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6143__A0 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6447_ _7022_/A _6447_/B vssd1 vssd1 vccd1 vccd1 _7929_/D sky130_fd_sc_hd__and2_1
X_6378_ _6412_/S _6088_/X _6128_/X vssd1 vssd1 vccd1 vccd1 _6378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6694__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8117_ _8117_/CLK _8117_/D vssd1 vssd1 vccd1 vccd1 _8117_/Q sky130_fd_sc_hd__dfxtp_2
X_5329_ _3814_/X _5299_/B _5331_/B1 hold985/X vssd1 vssd1 vccd1 vccd1 _5329_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6296__A _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5249__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3713__A _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8048_ _8048_/CLK _8048_/D vssd1 vssd1 vccd1 vccd1 _8048_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4552__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6749__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5709__A0 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4607__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5375__A _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3735__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6134__B1 _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6685__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4791__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5541__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6653__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4454__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4846__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7159__37 _7907_/CLK vssd1 vssd1 vccd1 vccd1 _8039_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_127_532 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4700_ _4699_/X _4698_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__mux2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _6551_/A _5680_/B vssd1 vssd1 vccd1 vccd1 _5680_/X sky130_fd_sc_hd__and2_1
XFILLER_0_127_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4631_ _4630_/X _4627_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7515_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6912__A2 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7350_ _8468_/CLK _7350_/D vssd1 vssd1 vccd1 vccd1 _7350_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4562_ _8332_/Q _7808_/Q _7474_/Q _7442_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4562_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_40_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold615 _7589_/Q vssd1 vssd1 vccd1 vccd1 hold615/X sky130_fd_sc_hd__dlygate4sd3_1
X_7281_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7281_/Y sky130_fd_sc_hd__inv_2
X_6301_ _6301_/A _6301_/B vssd1 vssd1 vccd1 vccd1 _6301_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_52_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold626 _6725_/X vssd1 vssd1 vccd1 vccd1 _8280_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _5166_/A1 _4392_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _7305_/D sky130_fd_sc_hd__mux2_1
Xhold604 _5214_/X vssd1 vssd1 vccd1 vccd1 _7428_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold659 _7808_/Q vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6676__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold637 _8370_/Q vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 _6561_/X vssd1 vssd1 vccd1 vccd1 _8133_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _8472_/CLK sky130_fd_sc_hd__clkbuf_16
X_6232_ _6414_/A2 _6229_/A _6231_/X vssd1 vssd1 vccd1 vccd1 _6232_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6163_ _6163_/A _6163_/B vssd1 vssd1 vccd1 vccd1 _6163_/Y sky130_fd_sc_hd__nand2_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7005__A _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5114_ input18/X _5144_/A2 _5146_/B1 _5113_/X vssd1 vssd1 vccd1 vccd1 _7369_/D sky130_fd_sc_hd__o211a_1
XANTENNA__5451__C _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1304 _8183_/Q vssd1 vssd1 vccd1 vccd1 _6638_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6094_ _6094_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6096_/B sky130_fd_sc_hd__xnor2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1315 _6964_/X vssd1 vssd1 vccd1 vccd1 _8447_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1348 _8332_/Q vssd1 vssd1 vccd1 vccd1 _6790_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4534__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1359 _6788_/X vssd1 vssd1 vccd1 vccd1 _8331_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 _8354_/Q vssd1 vssd1 vccd1 vccd1 _6834_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5045_ _5432_/A _5462_/C vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__or2_1
Xhold1337 _6640_/X vssd1 vssd1 vccd1 vccd1 _8184_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5651__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout449_A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4364__A _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6996_ _6981_/Y _6995_/Y _6990_/S vssd1 vssd1 vccd1 vccd1 _6996_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4083__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5947_ _5947_/A _5947_/B vssd1 vssd1 vccd1 vccd1 _5949_/A sky130_fd_sc_hd__nor2_1
XANTENNA__5179__B _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6039__S0 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5878_ _4095_/Y _5877_/X _6393_/A vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__mux2_1
X_7617_ _8504_/CLK _7617_/D vssd1 vssd1 vccd1 vccd1 _7617_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3708__A _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6364__B1 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4829_ _8463_/Q _8395_/Q _8427_/Q _8301_/Q _7063_/A _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4829_/X sky130_fd_sc_hd__mux4_1
X_7173__51 _8457_/CLK vssd1 vssd1 vccd1 vccd1 _8053_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7548_ _8413_/CLK _7548_/D vssd1 vssd1 vccd1 vccd1 _7548_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7479_ _8467_/CLK _7479_/D vssd1 vssd1 vccd1 vccd1 _7479_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5642__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4828__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5089__B _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3956__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4213__S _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5536__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6929__A _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6658__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output78_A _8123_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5330__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7083__B2 _7083_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4883__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5094__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6830__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5633__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6850_ _7010_/A _6850_/A2 _6842_/X _6849_/X vssd1 vssd1 vccd1 vccd1 _6850_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4819__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6781_ _6847_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6781_/X sky130_fd_sc_hd__and2_1
X_5801_ _5792_/Y _5793_/Y _5800_/X _5694_/Y vssd1 vssd1 vccd1 vccd1 _5801_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3993_ _3993_/A0 _6426_/B _4085_/S vssd1 vssd1 vccd1 vccd1 _5889_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_85_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5732_ _8453_/Q _4148_/B _5732_/C _5732_/D vssd1 vssd1 vccd1 vccd1 _5732_/X sky130_fd_sc_hd__and4bb_2
XFILLER_0_57_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5663_ _6494_/A _5663_/B vssd1 vssd1 vccd1 vccd1 _5663_/X sky130_fd_sc_hd__and2_1
X_8451_ _8451_/CLK _8451_/D vssd1 vssd1 vccd1 vccd1 _8451_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5594_ _6925_/A _5584_/B _5617_/B1 hold651/X vssd1 vssd1 vccd1 vccd1 _5594_/X sky130_fd_sc_hd__a22o_1
X_4614_ _8179_/Q _8211_/Q _8275_/Q _7783_/Q _4741_/S0 _4737_/S1 vssd1 vssd1 vccd1
+ vccd1 _4614_/X sky130_fd_sc_hd__mux4_1
X_7402_ _8030_/CLK _7402_/D vssd1 vssd1 vccd1 vccd1 _7402_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8382_ _8382_/CLK _8382_/D _7276_/Y vssd1 vssd1 vccd1 vccd1 _8382_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4545_ _8459_/Q _8391_/Q _8423_/Q _8297_/Q _4640_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4545_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_53_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold401 _5640_/X vssd1 vssd1 vccd1 vccd1 _7820_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7333_ _8504_/CLK _7333_/D vssd1 vssd1 vccd1 vccd1 _7333_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6839__A _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 _8315_/Q vssd1 vssd1 vccd1 vccd1 hold445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 hold412/A vssd1 vssd1 vccd1 vccd1 _4751_/B sky130_fd_sc_hd__clkbuf_2
Xhold434 _6747_/X vssd1 vssd1 vccd1 vccd1 _8298_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold423 _7588_/Q vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7264_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7264_/Y sky130_fd_sc_hd__inv_2
X_4476_ _7015_/A _7911_/Q vssd1 vssd1 vccd1 vccd1 _8043_/D sky130_fd_sc_hd__and2_1
Xhold478 _6768_/X vssd1 vssd1 vccd1 vccd1 _8319_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5462__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold467 _7431_/Q vssd1 vssd1 vccd1 vccd1 hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _6588_/X vssd1 vssd1 vccd1 vccd1 _8160_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4359__A _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold489 _7450_/Q vssd1 vssd1 vccd1 vccd1 hold489/X sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6157_/A _6175_/A _6191_/A _6209_/A _5782_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6215_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5321__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6146_ _6342_/S _6144_/S _4095_/Y _6198_/S vssd1 vssd1 vccd1 vccd1 _6146_/X sky130_fd_sc_hd__a31o_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1123 _8326_/Q vssd1 vssd1 vccd1 vccd1 _6778_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 _6419_/X vssd1 vssd1 vccd1 vccd1 _7901_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1101 _8283_/Q vssd1 vssd1 vccd1 vccd1 _6728_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1156 _6846_/X vssd1 vssd1 vccd1 vccd1 _8389_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5624__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1145 _8146_/Q vssd1 vssd1 vccd1 vccd1 _6574_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_6077_ _6058_/A _6057_/A _6055_/Y vssd1 vssd1 vccd1 vccd1 _6078_/B sky130_fd_sc_hd__a21o_1
Xhold1134 _6894_/X vssd1 vssd1 vccd1 vccd1 _8413_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 _7539_/Q vssd1 vssd1 vccd1 vccd1 _5308_/B2 sky130_fd_sc_hd__dlygate4sd3_1
X_5028_ hold637/X _4425_/B _5148_/B1 _5027_/X vssd1 vssd1 vccd1 vccd1 _5028_/X sky130_fd_sc_hd__o211a_1
Xhold1178 _6636_/X vssd1 vssd1 vccd1 vccd1 _8182_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 _8190_/Q vssd1 vssd1 vccd1 vccd1 _6652_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4094__A _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7232__110 _8143_/CLK vssd1 vssd1 vccd1 vccd1 _8242_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold1583_A _7368_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6979_ _6977_/B _6597_/B _5547_/B _6974_/A vssd1 vssd1 vccd1 vccd1 _6979_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_83_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6585__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6888__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4994__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5372__B _7344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold990 _5235_/X vssd1 vssd1 vccd1 vccd1 _7443_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5312__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6812__A1 _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6273__C1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6484__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5615__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1690 _7676_/Q vssd1 vssd1 vccd1 vccd1 _4012_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output116_A _7311_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6931__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6576__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3929__A2 _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5563__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6659__A _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4330_ _4328_/Y _4330_/B vssd1 vssd1 vccd1 vccd1 _4330_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5303__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4737__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4261_ _5566_/B _5034_/A1 _5503_/B vssd1 vssd1 vccd1 vccd1 _4262_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5854__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6000_ _6302_/A _5774_/B _5999_/Y _6083_/A vssd1 vssd1 vccd1 vccd1 _6000_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_66_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4192_ _4192_/A vssd1 vssd1 vccd1 vccd1 _4193_/C sky130_fd_sc_hd__inv_2
XANTENNA__5606__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7951_ _8011_/CLK hold70/X vssd1 vssd1 vccd1 vccd1 _7951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7882_ _8469_/CLK _7882_/D vssd1 vssd1 vccd1 vccd1 _7882_/Q sky130_fd_sc_hd__dfxtp_1
X_6902_ _7027_/A _6902_/A2 _6845_/B _6901_/X vssd1 vssd1 vccd1 vccd1 _6902_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_82_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6833_ _6965_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6833_/X sky130_fd_sc_hd__and2_1
XANTENNA__6567__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6031__A2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6764_ _6951_/A _6741_/B _6774_/B1 hold445/X vssd1 vssd1 vccd1 vccd1 _6764_/X sky130_fd_sc_hd__a22o_1
X_3976_ _7978_/Q _4079_/A2 _4079_/B1 _8010_/Q _3975_/X vssd1 vssd1 vccd1 vccd1 _3976_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5790__A1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5715_ _6352_/A _6370_/A _5716_/S vssd1 vssd1 vccd1 vccd1 _5715_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8503_ _8503_/CLK _8503_/D vssd1 vssd1 vccd1 vccd1 _8503_/Q sky130_fd_sc_hd__dfxtp_1
X_6695_ _6891_/A _6701_/A2 _6701_/B1 hold461/X vssd1 vssd1 vccd1 vccd1 _6695_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5457__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8434_ _8477_/CLK _8434_/D vssd1 vssd1 vccd1 vccd1 _8434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5646_ _6891_/A _5652_/A2 _5652_/B1 hold871/X vssd1 vssd1 vccd1 vccd1 _5646_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4788__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5473__A _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8365_ _8365_/CLK _8365_/D _7259_/Y vssd1 vssd1 vccd1 vccd1 _8365_/Q sky130_fd_sc_hd__dfrtp_1
X_5577_ _6520_/A _5577_/B vssd1 vssd1 vccd1 vccd1 _7766_/D sky130_fd_sc_hd__and2_1
XANTENNA__4976__S0 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 _7759_/Q vssd1 vssd1 vccd1 vccd1 _6510_/B sky130_fd_sc_hd__dlygate4sd3_1
X_7143__21 _8218_/CLK vssd1 vssd1 vccd1 vccd1 _7520_/CLK sky130_fd_sc_hd__inv_2
Xhold242 _8295_/Q vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _6673_/X vssd1 vssd1 vccd1 vccd1 _8200_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8296_ _8468_/CLK _8296_/D vssd1 vssd1 vccd1 vccd1 _8296_/Q sky130_fd_sc_hd__dfxtp_1
Xhold231 _5267_/X vssd1 vssd1 vccd1 vccd1 _7471_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ _8134_/Q _7533_/Q _7405_/Q _7565_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4528_/X sky130_fd_sc_hd__mux4_1
X_7316_ _8360_/CLK _7316_/D vssd1 vssd1 vccd1 vccd1 _7316_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold275 _6671_/X vssd1 vssd1 vccd1 vccd1 _8198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _7406_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _7532_/Q vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _6551_/A _7928_/Q vssd1 vssd1 vccd1 vccd1 _8060_/D sky130_fd_sc_hd__and2_1
Xhold297 _5433_/X vssd1 vssd1 vccd1 vccd1 _7622_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1429_A _7304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3856__A1 _3855_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6129_ _6309_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _6130_/B sky130_fd_sc_hd__nor2_2
XANTENNA__5058__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6022__A2 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5230__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5781__A1 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5383__A _7065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6730__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6479__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4719__S0 _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7103__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5695__S1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5558__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6661__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4462__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5221__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4024__A1 _4023_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3830_ _4773_/B _4072_/B _3829_/X vssd1 vssd1 vccd1 vccd1 _3830_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3761_ _4760_/B _4071_/A2 _4071_/B1 _3754_/X _3760_/X vssd1 vssd1 vccd1 vccd1 _6140_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5500_ _7521_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7689_/D sky130_fd_sc_hd__and3_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3692_ _7663_/Q _7837_/Q vssd1 vssd1 vccd1 vccd1 _3692_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_113_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6480_ _6545_/A hold73/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__and2_1
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6721__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7923__D _7923_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4958__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5431_ _5431_/A _5503_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _5431_/X sky130_fd_sc_hd__and3_1
X_8150_ _8339_/CLK _8150_/D vssd1 vssd1 vccd1 vccd1 _8150_/Q sky130_fd_sc_hd__dfxtp_1
X_5362_ _6959_/A _5335_/B _5368_/B1 hold615/X vssd1 vssd1 vccd1 vccd1 _5362_/X sky130_fd_sc_hd__a22o_1
X_7101_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7101_/Y sky130_fd_sc_hd__inv_2
X_8081_ _8469_/CLK _8115_/D vssd1 vssd1 vccd1 vccd1 _8081_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4313_ _8494_/Q _4314_/B vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__or2_1
X_7032_ _7074_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7032_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5288__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5293_ _6967_/A _5294_/A2 _5294_/B1 _5293_/B2 vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__a22o_1
X_4244_ _4242_/Y _4244_/B vssd1 vssd1 vccd1 vccd1 _4244_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__5740__B _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4175_ _4169_/A _4166_/Y _4168_/B vssd1 vssd1 vccd1 vccd1 _4176_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_93_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7013__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout264_A _5226_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7934_ _8480_/CLK _7934_/D vssd1 vssd1 vccd1 vccd1 _7934_/Q sky130_fd_sc_hd__dfxtp_1
X_7865_ _8385_/CLK _7865_/D vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
X_6816_ _7017_/A _6816_/A2 _6838_/A3 _6815_/X vssd1 vssd1 vccd1 vccd1 _6816_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7796_ _8479_/CLK _7796_/D vssd1 vssd1 vccd1 vccd1 _7796_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout431_A _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5212__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6747_ _6917_/A _6773_/A2 _6773_/B1 hold433/X vssd1 vssd1 vccd1 vccd1 _6747_/X sky130_fd_sc_hd__a22o_1
X_3959_ _4180_/A _3958_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _5918_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6678_ _6923_/A _6701_/A2 _6701_/B1 hold925/X vssd1 vssd1 vccd1 vccd1 _6678_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6712__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5629_ _6923_/A _5652_/A2 _5652_/B1 _5629_/B2 vssd1 vssd1 vccd1 vccd1 _5629_/X sky130_fd_sc_hd__a22o_1
X_8417_ _8485_/CLK _8417_/D vssd1 vssd1 vccd1 vccd1 _8417_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_115_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8348_ _8442_/CLK _8348_/D vssd1 vssd1 vccd1 vccd1 _8348_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4311__S _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8279_ _8461_/CLK _8279_/D vssd1 vssd1 vccd1 vccd1 _8279_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5279__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3829__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4981__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6794__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5203__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__B _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6937__A _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4457__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6219__C1 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5980_ _4045_/B _6105_/A2 _5978_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _5980_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_87_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4931_ _8155_/Q _7554_/Q _7426_/Q _7586_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4931_/X sky130_fd_sc_hd__mux4_1
X_4862_ _4860_/X _4861_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7650_ _8373_/CLK _7650_/D vssd1 vssd1 vccd1 vccd1 _7650_/Q sky130_fd_sc_hd__dfxtp_1
X_6601_ _6704_/B _6776_/B vssd1 vssd1 vccd1 vccd1 _6601_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _7999_/Q _4068_/A2 _4068_/B1 _8031_/Q _3812_/X vssd1 vssd1 vccd1 vccd1 _3813_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4793_ _8168_/Q _8200_/Q _8264_/Q _7772_/Q _5475_/A _4896_/S1 vssd1 vssd1 vccd1 vccd1
+ _4793_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7581_ _8343_/CLK _7581_/D vssd1 vssd1 vccd1 vccd1 _7581_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5745__A1 _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_15 _3757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6532_ _7008_/A _6532_/B vssd1 vssd1 vccd1 vccd1 _8014_/D sky130_fd_sc_hd__and2_1
XFILLER_0_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3756__B1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3744_ _4771_/B _4072_/B _3743_/X vssd1 vssd1 vccd1 vccd1 _6448_/B sky130_fd_sc_hd__a21oi_4
X_3675_ _3675_/A _3675_/B _3675_/C vssd1 vssd1 vccd1 vccd1 _3676_/B sky130_fd_sc_hd__and3_1
X_6463_ _6498_/A _6463_/B vssd1 vssd1 vccd1 vccd1 _6463_/X sky130_fd_sc_hd__and2_1
XFILLER_0_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7008__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput100 _7295_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[13] sky130_fd_sc_hd__buf_12
X_5414_ _5414_/A _7030_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _5414_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8202_ _8350_/CLK _8202_/D vssd1 vssd1 vccd1 vccd1 _8202_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8133_ _8428_/CLK _8133_/D vssd1 vssd1 vccd1 vccd1 _8133_/Q sky130_fd_sc_hd__dfxtp_1
X_7125__3 _8328_/CLK vssd1 vssd1 vccd1 vccd1 _7502_/CLK sky130_fd_sc_hd__inv_2
Xoutput122 _7287_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[5] sky130_fd_sc_hd__buf_12
X_6394_ _5952_/A _6392_/X _6008_/A vssd1 vssd1 vccd1 vccd1 _6394_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput133 _8050_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[15] sky130_fd_sc_hd__buf_12
XFILLER_0_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput111 _7306_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[24] sky130_fd_sc_hd__buf_12
Xoutput155 _8041_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[6] sky130_fd_sc_hd__buf_12
XANTENNA__6847__A _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5345_ _6925_/A _5335_/B _5368_/B1 _5345_/B2 vssd1 vssd1 vccd1 vccd1 _5345_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput144 _8060_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[25] sky130_fd_sc_hd__buf_12
X_5276_ _6933_/A _5262_/B _5295_/B1 hold665/X vssd1 vssd1 vccd1 vccd1 _5276_/X sky130_fd_sc_hd__a22o_1
X_8064_ _8064_/CLK _8064_/D vssd1 vssd1 vccd1 vccd1 _8064_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout381_A _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4227_ _4427_/A _4227_/B _4227_/C vssd1 vssd1 vccd1 vccd1 _4422_/A sky130_fd_sc_hd__and3_1
X_7015_ _7015_/A _7015_/B vssd1 vssd1 vccd1 vccd1 _7015_/X sky130_fd_sc_hd__and2_1
XANTENNA__5470__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4158_ _4161_/A _4161_/B _4158_/C vssd1 vssd1 vccd1 vccd1 _4159_/B sky130_fd_sc_hd__and3_1
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4089_ _4089_/A _4089_/B vssd1 vssd1 vccd1 vccd1 _4090_/D sky130_fd_sc_hd__and2_1
XFILLER_0_78_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7917_ _8010_/CLK _7917_/D vssd1 vssd1 vccd1 vccd1 _7917_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7848_ _8368_/CLK _7848_/D vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7779_ _8465_/CLK _7779_/D vssd1 vssd1 vccd1 vccd1 _7779_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1663_A _4028_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5831__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5661__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3880__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout382 _4737_/S1 vssd1 vssd1 vccd1 vccd1 _4639_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout393 _7072_/B2 vssd1 vssd1 vccd1 vccd1 _4741_/S0 sky130_fd_sc_hd__clkbuf_4
Xfanout360 _4079_/A2 vssd1 vssd1 vccd1 vccd1 _4068_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout371 _7048_/A vssd1 vssd1 vccd1 vccd1 _4735_/S sky130_fd_sc_hd__buf_4
XFILLER_0_17_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4570__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6492__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5539__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 i_instr_ID[22] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
Xinput35 i_read_data_M[13] vssd1 vssd1 vccd1 vccd1 _6534_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput46 i_read_data_M[23] vssd1 vssd1 vccd1 vccd1 _6544_/B sky130_fd_sc_hd__clkbuf_1
Xinput24 i_instr_ID[3] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold808 _5354_/X vssd1 vssd1 vccd1 vccd1 _7581_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput57 i_read_data_M[4] vssd1 vssd1 vccd1 vccd1 _6525_/B sky130_fd_sc_hd__buf_1
Xhold819 _7817_/Q vssd1 vssd1 vccd1 vccd1 hold819/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4886__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5571__A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5130_ _5130_/A1 _4448_/B _5140_/B1 _5129_/X vssd1 vssd1 vccd1 vccd1 _7377_/D sky130_fd_sc_hd__o211a_1
X_5061_ _5440_/A _7030_/C vssd1 vssd1 vccd1 vccd1 _5061_/X sky130_fd_sc_hd__or2_1
XANTENNA__6386__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1508 hold1815/X vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__buf_1
Xhold1519 _6912_/X vssd1 vssd1 vccd1 vccd1 _8421_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4012_ _4012_/A1 _4084_/A2 _6925_/A _4084_/B2 vssd1 vssd1 vccd1 vccd1 _4012_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_74_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5963_ _5857_/X _5859_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5963_/X sky130_fd_sc_hd__mux2_1
X_7702_ _8328_/CLK _7702_/D vssd1 vssd1 vccd1 vccd1 _7702_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4914_ _4913_/X _4912_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5449__C _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5894_ _5872_/A _5871_/A _5869_/Y vssd1 vssd1 vccd1 vccd1 _5895_/B sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_89_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4845_ _4844_/X _4841_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8239_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7633_ _8363_/CLK _7633_/D vssd1 vssd1 vccd1 vccd1 _7633_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3965__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4776_ _8326_/Q _7802_/Q _7468_/Q _7436_/Q _5475_/A _5476_/A vssd1 vssd1 vccd1 vccd1
+ _4776_/X sky130_fd_sc_hd__mux4_1
X_7564_ _7805_/CLK _7564_/D vssd1 vssd1 vccd1 vccd1 _7564_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5194__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3729__B1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6930__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout227_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3727_ _7995_/Q _4068_/A2 _4068_/B1 _8027_/Q _3726_/X vssd1 vssd1 vccd1 vccd1 _3727_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5465__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6515_ _6551_/A hold41/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__and2_1
XFILLER_0_130_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7495_ _8353_/CLK _7495_/D vssd1 vssd1 vccd1 vccd1 _7495_/Q sky130_fd_sc_hd__dfxtp_1
X_3658_ _7665_/Q vssd1 vssd1 vccd1 vccd1 _3658_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_70_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6446_ _6551_/A _6446_/B vssd1 vssd1 vccd1 vccd1 _7928_/D sky130_fd_sc_hd__and2_1
XANTENNA__4796__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6377_ _6309_/A _6376_/X _6083_/X _5740_/Y vssd1 vssd1 vccd1 vccd1 _6377_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6694__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_27_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8116_ _8116_/CLK _8116_/D vssd1 vssd1 vccd1 vccd1 _8116_/Q sky130_fd_sc_hd__dfxtp_2
X_5328_ _6963_/A _5299_/B _5331_/B1 hold897/X vssd1 vssd1 vccd1 vccd1 _5328_/X sky130_fd_sc_hd__a22o_1
X_8047_ _8047_/CLK _8047_/D vssd1 vssd1 vccd1 vccd1 _8047_/Q sky130_fd_sc_hd__dfxtp_1
X_5259_ _6971_/A _5226_/B _5259_/B1 hold967/X vssd1 vssd1 vccd1 vccd1 _5259_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_4_5_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_5_0_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__4552__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1780_A _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5709__A1 _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3875__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5656__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6382__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6685__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6487__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5391__A _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4791__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5645__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _5789_/S vssd1 vssd1 vccd1 vccd1 _5744_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7111__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5176__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4470__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4630_ _4629_/X _4628_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4630_/X sky130_fd_sc_hd__mux2_1
X_4561_ _4560_/X _4557_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7505_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6300_ _6283_/A _6282_/B _6280_/Y vssd1 vssd1 vccd1 vccd1 _6301_/B sky130_fd_sc_hd__a21o_1
Xhold616 _5362_/X vssd1 vssd1 vccd1 vccd1 _7589_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6125__B2 _5739_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6125__A1 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7280_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7280_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_40_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4492_ _5168_/A1 _4390_/B _5465_/C vssd1 vssd1 vccd1 vccd1 _7306_/D sky130_fd_sc_hd__mux2_1
Xhold627 _7550_/Q vssd1 vssd1 vccd1 vccd1 hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold605 _7831_/Q vssd1 vssd1 vccd1 vccd1 hold605/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6676__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold638 _5028_/X vssd1 vssd1 vccd1 vccd1 _7326_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ _3895_/A _6414_/B1 _6398_/B1 _6223_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6231_/X
+ sky130_fd_sc_hd__a221o_1
Xhold649 _7447_/Q vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6162_ _5999_/B _6302_/B _6342_/S vssd1 vssd1 vccd1 vccd1 _6162_/X sky130_fd_sc_hd__mux2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5113_ _7077_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5113_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 _8339_/Q vssd1 vssd1 vccd1 vccd1 _6804_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1305 _6638_/X vssd1 vssd1 vccd1 vccd1 _8183_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6093_ _6074_/Y _6078_/B _6076_/B vssd1 vssd1 vccd1 vccd1 _6098_/A sky130_fd_sc_hd__a21o_1
XANTENNA__5636__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1349 _6790_/X vssd1 vssd1 vccd1 vccd1 _8332_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4534__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1338 _8197_/Q vssd1 vssd1 vccd1 vccd1 _6666_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1327 _6834_/X vssd1 vssd1 vccd1 vccd1 _8354_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5044_ _4394_/A _4416_/B _5166_/B1 _5043_/X vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5100__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_A _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7021__A _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6061__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6995_ _5384_/X _6994_/X _6983_/B vssd1 vssd1 vccd1 vccd1 _6995_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_48_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5946_ _5946_/A _5946_/B vssd1 vssd1 vccd1 vccd1 _5947_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout344_A _3717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5877_ _5846_/A _5765_/A _5870_/A _5820_/A _5797_/S _5772_/S vssd1 vssd1 vccd1 vccd1
+ _5877_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6039__S1 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5476__A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _8173_/Q _8205_/Q _8269_/Q _7777_/Q _7063_/A _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4828_/X sky130_fd_sc_hd__mux4_1
X_7616_ _8071_/CLK _7616_/D vssd1 vssd1 vccd1 vccd1 _7616_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4759_ _7023_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _8116_/D sky130_fd_sc_hd__and2_1
X_7547_ _8467_/CLK _7547_/D vssd1 vssd1 vccd1 vccd1 _7547_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7478_ _8332_/CLK _7478_/D vssd1 vssd1 vccd1 vccd1 _7478_/Q sky130_fd_sc_hd__dfxtp_1
X_6429_ _6741_/A _6429_/B vssd1 vssd1 vccd1 vccd1 _7911_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3724__A _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5627__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5158__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6977__A_N _7356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6929__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7106__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5961__S0 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5330__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6945__A _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7219__97 _8454_/CLK vssd1 vssd1 vccd1 vccd1 _8132_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4465__A _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6780_ _7010_/A _6780_/A2 _6779_/B _6779_/Y vssd1 vssd1 vccd1 vccd1 _6780_/X sky130_fd_sc_hd__a31o_1
X_3992_ _3992_/A1 _4084_/A2 _6853_/A _4084_/B2 _3991_/X vssd1 vssd1 vccd1 vccd1 _6426_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6594__A1 _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5397__A2 _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5800_ _5796_/X _5799_/X _6302_/A vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__mux2_1
X_5731_ _5731_/A _5733_/D vssd1 vssd1 vccd1 vccd1 _5731_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3809__A _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5662_ _6498_/A _5662_/B vssd1 vssd1 vccd1 vccd1 _5662_/X sky130_fd_sc_hd__and2_1
XANTENNA__6346__B2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8450_ _8450_/CLK _8450_/D vssd1 vssd1 vccd1 vccd1 _8450_/Q sky130_fd_sc_hd__dfxtp_1
X_4613_ _4611_/X _4612_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4613_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_53_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5593_ _6923_/A _5616_/A2 _5616_/B1 hold929/X vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__a22o_1
X_7401_ _8501_/CLK _7401_/D vssd1 vssd1 vccd1 vccd1 _7401_/Q sky130_fd_sc_hd__dfxtp_1
X_8381_ _8382_/CLK _8381_/D _7275_/Y vssd1 vssd1 vccd1 vccd1 _8381_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4544_ _8169_/Q _8201_/Q _8265_/Q _7773_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4544_/X sky130_fd_sc_hd__mux4_1
Xhold402 _7580_/Q vssd1 vssd1 vccd1 vccd1 hold402/X sky130_fd_sc_hd__dlygate4sd3_1
X_7332_ _8091_/CLK _7332_/D vssd1 vssd1 vccd1 vccd1 _7332_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_123_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7263_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7263_/Y sky130_fd_sc_hd__inv_2
Xhold413 _7542_/Q vssd1 vssd1 vccd1 vccd1 hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _8267_/Q vssd1 vssd1 vccd1 vccd1 hold435/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6839__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold424 _5361_/X vssd1 vssd1 vccd1 vccd1 _7588_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _7007_/A _7912_/Q vssd1 vssd1 vccd1 vccd1 _8044_/D sky130_fd_sc_hd__and2_1
XANTENNA__5857__A0 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold446 _6764_/X vssd1 vssd1 vccd1 vccd1 _8315_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6214_ _5793_/Y _5878_/X _5739_/Y vssd1 vssd1 vccd1 vccd1 _6214_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_40_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold457 _7785_/Q vssd1 vssd1 vccd1 vccd1 hold457/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7016__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold468 _5217_/X vssd1 vssd1 vccd1 vccd1 _7431_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold479 _7466_/Q vssd1 vssd1 vccd1 vccd1 hold479/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5321__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6855__A _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6145_ _5982_/X _6144_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6145_/X sky130_fd_sc_hd__mux2_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1124 _6778_/X vssd1 vssd1 vccd1 vccd1 _8326_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6076_ _6076_/A _6076_/B vssd1 vssd1 vccd1 vccd1 _6078_/A sky130_fd_sc_hd__nor2_1
Xhold1102 _6728_/X vssd1 vssd1 vccd1 vccd1 _8283_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 _8427_/Q vssd1 vssd1 vccd1 vccd1 _6924_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5609__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5423_/A _5453_/C vssd1 vssd1 vccd1 vccd1 _5027_/X sky130_fd_sc_hd__or2_1
Xhold1146 _6574_/X vssd1 vssd1 vccd1 vccd1 _8146_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1135 _8393_/Q vssd1 vssd1 vccd1 vccd1 _6854_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1157 _8407_/Q vssd1 vssd1 vccd1 vccd1 _6882_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout461_A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1168 _5308_/X vssd1 vssd1 vccd1 vccd1 _7539_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _8375_/Q vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__dlygate4sd3_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6585__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5918__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6978_ _7355_/Q _6976_/B _6976_/Y _8527_/Z _6977_/X vssd1 vssd1 vccd1 vccd1 _6978_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1576_A _7365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5929_ _6008_/A _5928_/Y _5925_/X vssd1 vssd1 vccd1 vccd1 _5930_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4691__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4994__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold980 _5277_/X vssd1 vssd1 vccd1 vccd1 _7481_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5312__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold991 _8157_/Q vssd1 vssd1 vccd1 vccd1 hold991/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4984__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3874__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3901__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1680 _3795_/X vssd1 vssd1 vccd1 vccd1 _6440_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1691 _4013_/Y vssd1 vssd1 vccd1 vccd1 _6429_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6576__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output109_A _7304_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4682__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6328__A1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6659__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4737__S1 _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5934__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4260_ _4260_/A _4260_/B vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__xor2_1
X_4191_ _4190_/X _4437_/A _7082_/A vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__mux2_1
XANTENNA__4894__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7056__A2 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5067__A1 _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7950_ _8079_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 _7950_/Q sky130_fd_sc_hd__dfxtp_1
X_7881_ _8270_/CLK _7881_/D vssd1 vssd1 vccd1 vccd1 _7881_/Q sky130_fd_sc_hd__dfxtp_1
X_6901_ _6967_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6901_/X sky130_fd_sc_hd__and2_1
X_6832_ _7025_/A _6832_/A2 _6838_/A3 _6831_/X vssd1 vssd1 vccd1 vccd1 _6832_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6567__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3975_ _3923_/B _7946_/Q vssd1 vssd1 vccd1 vccd1 _3975_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_57_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6763_ _6949_/A _6773_/A2 _6773_/B1 hold378/X vssd1 vssd1 vccd1 vccd1 _6763_/X sky130_fd_sc_hd__a22o_1
X_5714_ _5712_/X _5713_/X _5838_/A vssd1 vssd1 vccd1 vccd1 _5714_/X sky130_fd_sc_hd__mux2_1
X_8502_ _8503_/CLK _8502_/D vssd1 vssd1 vccd1 vccd1 _8502_/Q sky130_fd_sc_hd__dfxtp_1
X_6694_ _6955_/A _6701_/A2 _6701_/B1 hold527/X vssd1 vssd1 vccd1 vccd1 _6694_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8433_ _8469_/CLK _8433_/D vssd1 vssd1 vccd1 vccd1 _8433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5645_ _6955_/A _5652_/A2 _5652_/B1 hold661/X vssd1 vssd1 vccd1 vccd1 _5645_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5473__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8364_ _8364_/CLK _8364_/D _7258_/Y vssd1 vssd1 vccd1 vccd1 _8364_/Q sky130_fd_sc_hd__dfrtp_1
Xhold210 _7605_/Q vssd1 vssd1 vccd1 vccd1 _5663_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5576_ _6524_/A _5576_/B vssd1 vssd1 vccd1 vccd1 _7765_/D sky130_fd_sc_hd__and2_1
XANTENNA_fanout307_A _5333_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4976__S1 _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold243 _6744_/X vssd1 vssd1 vccd1 vccd1 _8295_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8295_ _8456_/CLK _8295_/D vssd1 vssd1 vccd1 vccd1 _8295_/Q sky130_fd_sc_hd__dfxtp_1
X_4527_ _8327_/Q _7803_/Q _7469_/Q _7437_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4527_/X sky130_fd_sc_hd__mux4_1
X_7315_ _8361_/CLK _7315_/D vssd1 vssd1 vccd1 vccd1 _7315_/Q sky130_fd_sc_hd__dfxtp_1
Xhold232 _8361_/Q vssd1 vssd1 vccd1 vccd1 _4442_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6178__S0 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold221 _6510_/X vssd1 vssd1 vccd1 vccd1 _7992_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _7439_/Q vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _7805_/Q vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 _5192_/X vssd1 vssd1 vccd1 vccd1 _7406_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold265 _5301_/X vssd1 vssd1 vccd1 vccd1 _7532_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4458_ _7018_/A _7929_/Q vssd1 vssd1 vccd1 vccd1 _8061_/D sky130_fd_sc_hd__and2_1
Xhold298 _8294_/Q vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
X_6128_ _6128_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _6128_/X sky130_fd_sc_hd__or2_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4389_ _4389_/A _5067_/S vssd1 vssd1 vccd1 vccd1 _4389_/X sky130_fd_sc_hd__and2_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ _6008_/A _5875_/X _5955_/Y vssd1 vssd1 vccd1 vccd1 _6361_/B sky130_fd_sc_hd__a21oi_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1693_A _3967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5230__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4664__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5664__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6730__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4719__S1 _4741_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6495__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7239__117 _8445_/CLK vssd1 vssd1 vccd1 vccd1 _8249_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_99_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5221__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3760_ _3760_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3760_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3783__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3691_ _3652_/Y _7834_/Q _3653_/Y _7661_/Q _3688_/X vssd1 vssd1 vccd1 vccd1 _3696_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5574__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5430_ _5430_/A _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _5430_/X sky130_fd_sc_hd__and3_1
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6721__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4958__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3806__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5361_ _6891_/A _5367_/A2 _5367_/B1 hold423/X vssd1 vssd1 vccd1 vccd1 _5361_/X sky130_fd_sc_hd__a22o_1
X_8080_ _8080_/CLK _8114_/D vssd1 vssd1 vccd1 vccd1 _8080_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7100_ _7258_/A vssd1 vssd1 vccd1 vccd1 _7100_/Y sky130_fd_sc_hd__inv_2
X_5292_ _6965_/A _5294_/A2 _5294_/B1 hold747/X vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4312_ _4390_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__nand2_1
X_7031_ _7031_/A _7079_/C vssd1 vssd1 vccd1 vccd1 _7031_/Y sky130_fd_sc_hd__nand2_4
XANTENNA__5288__A1 _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4243_ _8504_/Q _4243_/B vssd1 vssd1 vccd1 vccd1 _4243_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_93_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4174_ _4174_/A _4174_/B vssd1 vssd1 vccd1 vccd1 _4174_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6788__A1 _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7933_ _8360_/CLK _7933_/D vssd1 vssd1 vccd1 vccd1 _7933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7864_ _8387_/CLK hold52/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout257_A _5335_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7795_ _8445_/CLK _7795_/D vssd1 vssd1 vccd1 vccd1 _7795_/Q sky130_fd_sc_hd__dfxtp_1
X_6815_ _6815_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6815_/X sky130_fd_sc_hd__and2_1
XFILLER_0_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5468__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5212__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6746_ _6849_/A _6741_/B _6774_/B1 hold891/X vssd1 vssd1 vccd1 vccd1 _6746_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_107_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_A hold1747/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7203__81 _8484_/CLK vssd1 vssd1 vccd1 vccd1 _8116_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4646__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4799__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3958_ _3958_/A1 _4084_/A2 _3954_/X _4084_/B2 _3957_/X vssd1 vssd1 vccd1 vccd1 _3958_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__6960__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3774__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6677_ _6921_/A _6669_/B _6702_/B1 hold417/X vssd1 vssd1 vccd1 vccd1 _6677_/X sky130_fd_sc_hd__a22o_1
X_3889_ _4765_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _3889_/X sky130_fd_sc_hd__and2_1
XFILLER_0_61_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6712__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5628_ _6921_/A _5620_/B _5653_/B1 hold659/X vssd1 vssd1 vccd1 vccd1 _5628_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_115_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8416_ _8448_/CLK _8416_/D vssd1 vssd1 vccd1 vccd1 _8416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5559_ _6534_/A _5559_/B vssd1 vssd1 vccd1 vccd1 _7748_/D sky130_fd_sc_hd__and2_1
X_8347_ _8413_/CLK _8347_/D vssd1 vssd1 vccd1 vccd1 _8347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1441_A _7295_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8278_ _8477_/CLK _8278_/D vssd1 vssd1 vccd1 vccd1 _8278_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5279__A1 _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3829__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5659__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4885__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5203__A1 _4080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6400__B1 _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4502__S _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6164__C1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6937__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7114__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6219__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6953__A _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5569__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4473__A _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4930_ _8348_/Q _7824_/Q _7490_/Q _7458_/Q _4987_/S0 _4976_/S1 vssd1 vssd1 vccd1
+ vccd1 _4930_/X sky130_fd_sc_hd__mux4_1
X_4861_ _8145_/Q _7544_/Q _7416_/Q _7576_/Q _4896_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4861_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6600_ _6600_/A _6600_/B _6600_/C vssd1 vssd1 vccd1 vccd1 _8165_/D sky130_fd_sc_hd__and3_1
X_3812_ _4067_/A_N _7967_/Q vssd1 vssd1 vccd1 vccd1 _3812_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4628__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4792_ _4790_/X _4791_/X _7359_/Q vssd1 vssd1 vccd1 vccd1 _4792_/X sky130_fd_sc_hd__mux2_1
X_7580_ _8402_/CLK _7580_/D vssd1 vssd1 vccd1 vccd1 _7580_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6942__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5745__A2 _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 _3757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6531_ _7007_/A _6531_/B vssd1 vssd1 vccd1 vccd1 _8013_/D sky130_fd_sc_hd__and2_1
XFILLER_0_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3756__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3743_ _3743_/A1 _4073_/A2 _6963_/A _4073_/B2 vssd1 vssd1 vccd1 vccd1 _3743_/X sky130_fd_sc_hd__a22o_1
X_3674_ _5222_/B _7665_/Q _3663_/X _7936_/Q vssd1 vssd1 vccd1 vccd1 _3675_/C sky130_fd_sc_hd__o211a_1
X_6462_ _6539_/A _6462_/B vssd1 vssd1 vccd1 vccd1 _6462_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput101 _7296_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[14] sky130_fd_sc_hd__buf_12
X_8201_ _8338_/CLK _8201_/D vssd1 vssd1 vccd1 vccd1 _8201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6393_ _6393_/A _6393_/B vssd1 vssd1 vccd1 vccd1 _6393_/X sky130_fd_sc_hd__or2_1
X_5413_ _5413_/A _5470_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _5413_/X sky130_fd_sc_hd__and3_1
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4800__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8132_ _8132_/CLK _8132_/D vssd1 vssd1 vccd1 vccd1 _8132_/Q sky130_fd_sc_hd__dfxtp_2
X_5344_ _6923_/A _5367_/A2 _5367_/B1 hold959/X vssd1 vssd1 vccd1 vccd1 _5344_/X sky130_fd_sc_hd__a22o_1
Xoutput134 _8051_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[16] sky130_fd_sc_hd__buf_12
Xoutput123 _7288_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[6] sky130_fd_sc_hd__buf_12
XFILLER_0_2_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput112 _7307_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[25] sky130_fd_sc_hd__buf_12
XANTENNA__6847__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput145 _8061_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[26] sky130_fd_sc_hd__buf_12
Xoutput156 _8042_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[7] sky130_fd_sc_hd__buf_12
X_5275_ _6931_/A _5294_/A2 _5294_/B1 hold823/X vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__a22o_1
X_8063_ _8063_/CLK _8063_/D vssd1 vssd1 vccd1 vccd1 _8063_/Q sky130_fd_sc_hd__dfxtp_1
X_4226_ _4225_/X _5024_/A1 _5453_/B vssd1 vssd1 vccd1 vccd1 _4227_/C sky130_fd_sc_hd__mux2_1
XANTENNA__5130__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7014_ _7017_/A _7014_/B vssd1 vssd1 vccd1 vccd1 _7014_/X sky130_fd_sc_hd__and2_1
XANTENNA__5470__C _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7024__A _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6863__A _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4157_ _8517_/Q _4161_/B _4158_/C vssd1 vssd1 vccd1 vccd1 _4157_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout374_A _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4867__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4088_ _6075_/A _6072_/A vssd1 vssd1 vccd1 vccd1 _4089_/B sky130_fd_sc_hd__nand2_1
X_7916_ _8471_/CLK _7916_/D vssd1 vssd1 vccd1 vccd1 _7916_/Q sky130_fd_sc_hd__dfxtp_1
X_7847_ _7907_/CLK _7847_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__8005__D _8005_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4619__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5197__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7778_ _8428_/CLK _7778_/D vssd1 vssd1 vccd1 vccd1 _7778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6729_ _6953_/A _6737_/A2 _6737_/B1 hold793/X vssd1 vssd1 vccd1 vccd1 _6729_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold1656_A _3890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_112_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8486_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6697__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout350 _5732_/X vssd1 vssd1 vccd1 vccd1 _6413_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout383 _4737_/S1 vssd1 vssd1 vccd1 vccd1 _4640_/S1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout361 _3679_/X vssd1 vssd1 vccd1 vccd1 _4079_/A2 sky130_fd_sc_hd__buf_8
Xfanout372 hold1637/X vssd1 vssd1 vccd1 vccd1 _7048_/A sky130_fd_sc_hd__buf_6
XFILLER_0_17_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout394 _7072_/B2 vssd1 vssd1 vccd1 vccd1 _4640_/S0 sky130_fd_sc_hd__buf_8
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6924__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7194__72 _8143_/CLK vssd1 vssd1 vccd1 vccd1 _8107_/CLK sky130_fd_sc_hd__inv_2
Xinput36 i_read_data_M[14] vssd1 vssd1 vccd1 vccd1 _6535_/B sky130_fd_sc_hd__clkbuf_1
Xinput14 i_instr_ID[23] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__buf_1
XFILLER_0_64_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_103_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _8478_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput25 i_instr_ID[4] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__7109__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6688__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold809 _7421_/Q vssd1 vssd1 vccd1 vccd1 hold809/X sky130_fd_sc_hd__dlygate4sd3_1
Xinput47 i_read_data_M[24] vssd1 vssd1 vccd1 vccd1 _6545_/B sky130_fd_sc_hd__clkbuf_1
Xinput58 i_read_data_M[5] vssd1 vssd1 vccd1 vccd1 _6526_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6152__A2 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5360__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4468__A _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5060_ _5060_/A1 _5069_/S _5182_/B1 _5059_/X vssd1 vssd1 vccd1 vccd1 _7342_/D sky130_fd_sc_hd__o211a_1
X_4011_ _8075_/Q _4010_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4011_/X sky130_fd_sc_hd__mux2_2
Xhold1509 _7737_/Q vssd1 vssd1 vccd1 vccd1 _4155_/B1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7929__D _7929_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4849__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5299__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5962_ _5853_/C _5961_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _5962_/X sky130_fd_sc_hd__mux2_1
X_7701_ _8464_/CLK _7701_/D vssd1 vssd1 vccd1 vccd1 _7701_/Q sky130_fd_sc_hd__dfxtp_1
X_4913_ _8475_/Q _8407_/Q _8439_/Q _8313_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4913_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_114_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5893_ _5893_/A _5893_/B vssd1 vssd1 vccd1 vccd1 _5895_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_74_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4844_ _4843_/X _4842_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7632_ _8387_/CLK _7632_/D vssd1 vssd1 vccd1 vccd1 _7632_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7563_ _8487_/CLK _7563_/D vssd1 vssd1 vccd1 vccd1 _7563_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4775_ _4775_/A _4775_/B vssd1 vssd1 vccd1 vccd1 _8132_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3729__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7019__A _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6514_ _6524_/A hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__and2_1
X_3726_ _4067_/A_N _7963_/Q vssd1 vssd1 vccd1 vccd1 _3726_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5465__C _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6679__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7494_ _8353_/CLK _7494_/D vssd1 vssd1 vccd1 vccd1 _7494_/Q sky130_fd_sc_hd__dfxtp_1
X_6445_ _7258_/A _6445_/B vssd1 vssd1 vccd1 vccd1 _7927_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_113_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5762__A _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6143__A2 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3657_ _3968_/A vssd1 vssd1 vccd1 vccd1 _3657_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5351__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6376_ _6235_/B _6375_/X _6411_/S vssd1 vssd1 vccd1 vccd1 _6376_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5481__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8115_ _8115_/CLK _8115_/D vssd1 vssd1 vccd1 vccd1 _8115_/Q sky130_fd_sc_hd__dfxtp_1
X_5327_ _6961_/A _5299_/B _5331_/B1 hold949/X vssd1 vssd1 vccd1 vccd1 _5327_/X sky130_fd_sc_hd__a22o_1
X_8046_ _8046_/CLK _8046_/D vssd1 vssd1 vccd1 vccd1 _8046_/Q sky130_fd_sc_hd__dfxtp_1
X_5258_ _6969_/A _5258_/A2 _5258_/B1 hold479/X vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__a22o_1
X_5189_ _6706_/A _5189_/B vssd1 vssd1 vccd1 vccd1 _5189_/Y sky130_fd_sc_hd__nand2_1
X_4209_ _8509_/Q _4209_/B vssd1 vssd1 vccd1 vccd1 _4209_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5701__S _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5002__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6906__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5590__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6134__A2 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3891__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5342__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5645__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 _5716_/S vssd1 vssd1 vccd1 vccd1 _5789_/S sky130_fd_sc_hd__clkbuf_8
Xfanout180 _6251_/A vssd1 vssd1 vccd1 vccd1 _6309_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__3959__A1 _3958_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6070__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6070__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4751__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4559_/X _4558_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4560_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_123_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4897__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold617 _8325_/Q vssd1 vssd1 vccd1 vccd1 hold617/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4491_ _5170_/A1 _4387_/B _5465_/C vssd1 vssd1 vccd1 vccd1 _7307_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold606 _5651_/X vssd1 vssd1 vccd1 vccd1 _7831_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold639 _7425_/Q vssd1 vssd1 vccd1 vccd1 hold639/X sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ _6309_/A _5902_/Y _6130_/A vssd1 vssd1 vccd1 vccd1 _6230_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4136__B2 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold628 _5319_/X vssd1 vssd1 vccd1 vccd1 _7550_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6161_ _6079_/X _6160_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6302_/B sky130_fd_sc_hd__mux2_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5112_ input17/X _5099_/B _5148_/B1 _5111_/X vssd1 vssd1 vccd1 vccd1 _7368_/D sky130_fd_sc_hd__o211a_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ _6086_/X _6087_/X _6090_/X _6091_/Y vssd1 vssd1 vccd1 vccd1 _6092_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5636__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3752__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1306 _8188_/Q vssd1 vssd1 vccd1 vccd1 _6648_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1317 _6804_/X vssd1 vssd1 vccd1 vccd1 _8339_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1339 _6666_/X vssd1 vssd1 vccd1 vccd1 _8197_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5431_/A _5454_/C vssd1 vssd1 vccd1 vccd1 _5043_/X sky130_fd_sc_hd__or2_1
Xhold1328 _8193_/Q vssd1 vssd1 vccd1 vccd1 _6658_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_7_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6994_ _7074_/A _6593_/X _6993_/X _5397_/Y vssd1 vssd1 vccd1 vccd1 _6994_/X sky130_fd_sc_hd__a2bb2o_1
X_5945_ _5946_/A _5946_/B vssd1 vssd1 vccd1 vccd1 _5945_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5876_ _5873_/X _5875_/X _6270_/A vssd1 vssd1 vccd1 vccd1 _5876_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5476__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4827_ _4825_/X _4826_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__mux2_1
X_7615_ _8379_/CLK _7615_/D vssd1 vssd1 vccd1 vccd1 _7615_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6364__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7546_ _8473_/CLK _7546_/D vssd1 vssd1 vccd1 vccd1 _7546_/Q sky130_fd_sc_hd__dfxtp_1
X_4758_ _7029_/A _4758_/B vssd1 vssd1 vccd1 vccd1 _8115_/D sky130_fd_sc_hd__and2_1
XFILLER_0_71_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7477_ _8461_/CLK _7477_/D vssd1 vssd1 vccd1 vccd1 _7477_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3709_ _3683_/X _4073_/B2 _4073_/A2 _3709_/B2 _3707_/X vssd1 vssd1 vccd1 vccd1 _3709_/X
+ sky130_fd_sc_hd__a221o_2
X_4689_ _8157_/Q _7556_/Q _7428_/Q _7588_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4689_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5324__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6428_ _6545_/A _6428_/B vssd1 vssd1 vccd1 vccd1 _7910_/D sky130_fd_sc_hd__and2_1
XANTENNA__5875__A1 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6359_ _6217_/C _6358_/X _6411_/S vssd1 vssd1 vccd1 vccd1 _6359_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5627__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8029_ _8029_/CLK _8029_/D vssd1 vssd1 vccd1 vccd1 _8029_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_98_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4063__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3886__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5667__A _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7164__42 _8426_/CLK vssd1 vssd1 vccd1 vccd1 _8044_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6498__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_73_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5315__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6658__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7068__B1 _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5961__S1 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3877__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6945__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_88_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4746__A _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5094__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7122__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6830__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6961__A _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3991_ hold55/X _4083_/B vssd1 vssd1 vccd1 vccd1 _3991_/X sky130_fd_sc_hd__and2_1
XANTENNA__6594__A2 _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5730_ _5730_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _5733_/D sky130_fd_sc_hd__or2_1
XANTENNA__4481__A _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5577__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5661_ _6539_/A _5661_/B vssd1 vssd1 vccd1 vccd1 _5661_/X sky130_fd_sc_hd__and2_1
XFILLER_0_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7400_ _8385_/CLK _7400_/D vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_127_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5592_ _6921_/A _5584_/B _5617_/B1 hold392/X vssd1 vssd1 vccd1 vccd1 _5592_/X sky130_fd_sc_hd__a22o_1
X_4612_ _8146_/Q _7545_/Q _7417_/Q _7577_/Q _4741_/S0 _4737_/S1 vssd1 vssd1 vccd1
+ vccd1 _4612_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8380_ _8382_/CLK _8380_/D _7274_/Y vssd1 vssd1 vccd1 vccd1 _8380_/Q sky130_fd_sc_hd__dfrtp_1
Xclkbuf_4_4_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_4_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_4543_ _4541_/X _4542_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4543_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7331_ _8504_/CLK _7331_/D vssd1 vssd1 vccd1 vccd1 _7331_/Q sky130_fd_sc_hd__dfxtp_1
Xhold425 _8300_/Q vssd1 vssd1 vccd1 vccd1 hold425/X sky130_fd_sc_hd__dlygate4sd3_1
X_7262_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7262_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5306__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold414 _5311_/X vssd1 vssd1 vccd1 vccd1 _7542_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _6712_/X vssd1 vssd1 vccd1 vccd1 _8267_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 _5353_/X vssd1 vssd1 vccd1 vccd1 _7580_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold469 _8199_/Q vssd1 vssd1 vccd1 vccd1 hold469/X sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _6552_/A _7913_/Q vssd1 vssd1 vccd1 vccd1 _8045_/D sky130_fd_sc_hd__and2_1
XFILLER_0_111_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5857__A1 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold447 _7420_/Q vssd1 vssd1 vccd1 vccd1 hold447/X sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6008_/A _6362_/B _6130_/A _5876_/X _6251_/A vssd1 vssd1 vccd1 vccd1 _6213_/X
+ sky130_fd_sc_hd__o32a_1
Xhold458 _5601_/X vssd1 vssd1 vccd1 vccd1 _7785_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6855__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6144_ _6064_/X _6143_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _6144_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5609__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6076_/B sky130_fd_sc_hd__nor2_1
Xhold1103 _8155_/Q vssd1 vssd1 vccd1 vccd1 _6583_/B2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 _6924_/X vssd1 vssd1 vccd1 vccd1 _8427_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _4421_/A _4425_/B _5148_/B1 _5025_/X vssd1 vssd1 vccd1 vccd1 _5026_/X sky130_fd_sc_hd__o211a_1
Xhold1136 _6854_/X vssd1 vssd1 vccd1 vccd1 _8393_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7032__A _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1158 _6882_/X vssd1 vssd1 vccd1 vccd1 _8407_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1147 _8395_/Q vssd1 vssd1 vccd1 vccd1 _6858_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 _8440_/Q vssd1 vssd1 vccd1 vccd1 _6950_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 _8349_/Q vssd1 vssd1 vccd1 vccd1 _6824_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout454_A _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6871__A _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4094__C _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_92_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _8090_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6977_ _7356_/Q _6977_/B _7354_/Q _7071_/A vssd1 vssd1 vccd1 vccd1 _6977_/X sky130_fd_sc_hd__and4b_1
X_5928_ _5952_/A _5812_/X _5836_/B vssd1 vssd1 vccd1 vccd1 _5928_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6585__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4691__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5859_ _5779_/X _5782_/X _5859_/S vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6888__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7529_ _7529_/CLK _7529_/D vssd1 vssd1 vccd1 vccd1 _7529_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold981 _8150_/Q vssd1 vssd1 vccd1 vccd1 hold981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold970 _6727_/X vssd1 vssd1 vccd1 vccd1 _8282_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 _6585_/X vssd1 vssd1 vccd1 vccd1 _8157_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5076__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6273__A1 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6812__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1670 _4059_/X vssd1 vssd1 vccd1 vccd1 _6433_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1681 _8509_/Q vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6781__A _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_83_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _8382_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1692 _7672_/Q vssd1 vssd1 vccd1 vccd1 _3967_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_129_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4505__S _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6576__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4682__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4240__S _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7117__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5839__A1 _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5934__S1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4190_ _4190_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4190_/X sky130_fd_sc_hd__xor2_1
XANTENNA__4476__A _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7880_ _8428_/CLK _7880_/D vssd1 vssd1 vccd1 vccd1 _7880_/Q sky130_fd_sc_hd__dfxtp_1
X_6900_ _7023_/A _6900_/A2 _6906_/A3 _6899_/X vssd1 vssd1 vccd1 vccd1 _6900_/X sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_74_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _8501_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6831_ _6963_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6831_/X sky130_fd_sc_hd__and2_1
XANTENNA__6567__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3974_ _6163_/A _5870_/A vssd1 vssd1 vccd1 vccd1 _3974_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6762_ _6947_/A _6773_/A2 _6773_/B1 hold881/X vssd1 vssd1 vccd1 vccd1 _6762_/X sky130_fd_sc_hd__a22o_1
X_8501_ _8501_/CLK _8501_/D vssd1 vssd1 vccd1 vccd1 _8501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5713_ _6318_/A _6334_/A _5716_/S vssd1 vssd1 vccd1 vccd1 _5713_/X sky130_fd_sc_hd__mux2_1
X_6693_ _6953_/A _6701_/A2 _6701_/B1 hold631/X vssd1 vssd1 vccd1 vccd1 _6693_/X sky130_fd_sc_hd__a22o_1
X_8432_ _8466_/CLK _8432_/D vssd1 vssd1 vccd1 vccd1 _8432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5644_ _6953_/A _5652_/A2 _5652_/B1 hold763/X vssd1 vssd1 vccd1 vccd1 _5644_/X sky130_fd_sc_hd__a22o_1
X_8363_ _8363_/CLK _8363_/D _7257_/Y vssd1 vssd1 vccd1 vccd1 _8363_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7314_ _8364_/CLK _7314_/D vssd1 vssd1 vccd1 vccd1 _7314_/Q sky130_fd_sc_hd__dfxtp_1
Xhold211 _5663_/X vssd1 vssd1 vccd1 vccd1 _7843_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold200 _7621_/Q vssd1 vssd1 vccd1 vccd1 _5679_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7027__A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5575_ _6551_/A _5575_/B vssd1 vssd1 vccd1 vccd1 _7764_/D sky130_fd_sc_hd__and2_1
X_8294_ _8456_/CLK _8294_/D vssd1 vssd1 vccd1 vccd1 _8294_/Q sky130_fd_sc_hd__dfxtp_1
Xhold244 _7323_/Q vssd1 vssd1 vccd1 vccd1 _5420_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4526_ _4525_/X _4522_/X _7365_/Q vssd1 vssd1 vccd1 vccd1 _7500_/D sky130_fd_sc_hd__mux2_1
Xhold222 _7377_/Q vssd1 vssd1 vccd1 vccd1 _5444_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _5010_/X vssd1 vssd1 vccd1 vccd1 _7317_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6178__S1 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold255 _5231_/X vssd1 vssd1 vccd1 vccd1 _7439_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _5625_/X vssd1 vssd1 vccd1 vccd1 _7805_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _8383_/Q vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _7018_/A _7930_/Q vssd1 vssd1 vccd1 vccd1 _8062_/D sky130_fd_sc_hd__and2_1
Xhold299 _6743_/X vssd1 vssd1 vccd1 vccd1 _8294_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold288 _7338_/Q vssd1 vssd1 vccd1 vccd1 _5435_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6127_ _6128_/A _6128_/B vssd1 vssd1 vccd1 vccd1 _6130_/A sky130_fd_sc_hd__nor2_4
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4388_ _5050_/A1 _4387_/Y _5465_/C vssd1 vssd1 vccd1 vccd1 _8381_/D sky130_fd_sc_hd__mux2_1
XANTENNA__6255__B2 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5058__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6058_/A _6058_/B vssd1 vssd1 vccd1 vccd1 _6058_/Y sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_65_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _8365_/CLK sky130_fd_sc_hd__clkbuf_16
X_5009_ _7317_/Q _7030_/C vssd1 vssd1 vccd1 vccd1 _5009_/X sky130_fd_sc_hd__or2_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1686_A _7356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4018__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5230__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4664__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5945__A _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4060__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7134__12 _8448_/CLK vssd1 vssd1 vccd1 vccd1 _7511_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_44_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6730__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4995__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5680__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_56_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _8507_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output121_A _7286_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3963__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6016__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5221__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5852__S0 _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3783__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3690_ _7661_/Q _7660_/Q _7663_/Q _7662_/Q vssd1 vssd1 vccd1 vccd1 _3690_/Y sky130_fd_sc_hd__nor4_1
XFILLER_0_82_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6721__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5360_ _6955_/A _5367_/A2 _5367_/B1 hold515/X vssd1 vssd1 vccd1 vccd1 _5360_/X sky130_fd_sc_hd__a22o_1
X_7222__100 _8328_/CLK vssd1 vssd1 vccd1 vccd1 _8232_/CLK sky130_fd_sc_hd__inv_2
X_5291_ _6963_/A _5294_/A2 _5294_/B1 hold745/X vssd1 vssd1 vccd1 vccd1 _5291_/X sky130_fd_sc_hd__a22o_1
X_4311_ _5573_/B _4389_/A _5465_/B vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__mux2_1
X_7030_ _7031_/A _7030_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _7030_/X sky130_fd_sc_hd__and3_1
XANTENNA__5288__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4242_ _8504_/Q _4243_/B vssd1 vssd1 vccd1 vccd1 _4242_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3822__B _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4591__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4173_ _8514_/Q _4173_/B vssd1 vssd1 vccd1 vccd1 _4173_/Y sky130_fd_sc_hd__nand2_1
X_7932_ _8483_/CLK _7932_/D vssd1 vssd1 vccd1 vccd1 _7932_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_47_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8519_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7863_ _8030_/CLK _7863_/D vssd1 vssd1 vccd1 vccd1 _7863_/Q sky130_fd_sc_hd__dfxtp_1
X_7794_ _8460_/CLK _7794_/D vssd1 vssd1 vccd1 vccd1 _7794_/Q sky130_fd_sc_hd__dfxtp_1
X_6814_ _7028_/A _6814_/A2 _6838_/A3 _6813_/X vssd1 vssd1 vccd1 vccd1 _6814_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_133_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6745_ _6847_/A _6741_/B _6774_/B1 hold483/X vssd1 vssd1 vccd1 vccd1 _6745_/X sky130_fd_sc_hd__a22o_1
X_3957_ _4750_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__and2_1
XFILLER_0_45_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5212__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4646__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5484__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6676_ _6853_/A _6669_/B _6702_/B1 hold757/X vssd1 vssd1 vccd1 vccd1 _6676_/X sky130_fd_sc_hd__a22o_1
X_3888_ _4765_/B _3676_/A _4082_/B1 _3886_/X _3887_/X vssd1 vssd1 vccd1 vccd1 _6226_/A
+ sky130_fd_sc_hd__o221a_4
X_8415_ _8483_/CLK _8415_/D vssd1 vssd1 vccd1 vccd1 _8415_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout417_A _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6712__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5627_ _6853_/A _5620_/B _5653_/B1 hold825/X vssd1 vssd1 vccd1 vccd1 _5627_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5558_ _6498_/A _5558_/B vssd1 vssd1 vccd1 vccd1 _7747_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8346_ _8346_/CLK _8346_/D vssd1 vssd1 vccd1 vccd1 _8346_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4509_ _5134_/A1 _4509_/A1 _7082_/B vssd1 vssd1 vccd1 vccd1 _7289_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8277_ _8471_/CLK _8277_/D vssd1 vssd1 vccd1 vccd1 _8277_/Q sky130_fd_sc_hd__dfxtp_1
X_5489_ _7510_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7678_/D sky130_fd_sc_hd__and3_1
XANTENNA__5279__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3986__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _8326_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4885__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5203__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5675__A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3923__A _7282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4573__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4754__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6953__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8426_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4860_ _8338_/Q _7814_/Q _7480_/Q _7448_/Q _4896_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4860_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_75_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3811_ _3811_/A _3811_/B vssd1 vssd1 vccd1 vccd1 _3848_/A sky130_fd_sc_hd__and2_1
XANTENNA__4628__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5585__A _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4791_ _8135_/Q _7534_/Q _7406_/Q _7566_/Q _4895_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4791_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6180__S _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5745__A3 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_17 _6343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6530_ _7024_/A _6530_/B vssd1 vssd1 vccd1 vccd1 _8012_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3756__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3742_ _4771_/B _4071_/A2 _4071_/B1 _3740_/X _3741_/X vssd1 vssd1 vccd1 vccd1 _6334_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_125_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ _5296_/A _7664_/Q _7666_/Q _5581_/A _3672_/Y vssd1 vssd1 vccd1 vccd1 _3675_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_103_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6461_ _6520_/A _6461_/B vssd1 vssd1 vccd1 vccd1 _6461_/X sky130_fd_sc_hd__and2_1
X_8200_ _8326_/CLK _8200_/D vssd1 vssd1 vccd1 vccd1 _8200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5412_ _5412_/A _7082_/A _5442_/C vssd1 vssd1 vccd1 vccd1 _5412_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6392_ _6334_/A _6352_/A _6370_/A _6388_/A _5772_/S _5804_/A vssd1 vssd1 vccd1 vccd1
+ _6392_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4800__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _6921_/A _5335_/B _5368_/B1 hold623/X vssd1 vssd1 vccd1 vccd1 _5343_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput124 _7289_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[7] sky130_fd_sc_hd__buf_12
X_8131_ _8131_/CLK _8131_/D vssd1 vssd1 vccd1 vccd1 _8131_/Q sky130_fd_sc_hd__dfxtp_2
Xoutput113 _7308_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[26] sky130_fd_sc_hd__buf_12
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput102 _7297_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[15] sky130_fd_sc_hd__buf_12
Xoutput135 _8052_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[17] sky130_fd_sc_hd__buf_12
Xoutput146 _8062_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[27] sky130_fd_sc_hd__buf_12
Xoutput157 _8043_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[8] sky130_fd_sc_hd__buf_12
X_5274_ _6929_/A _5262_/B _5295_/B1 hold597/X vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__a22o_1
X_8062_ _8062_/CLK _8062_/D vssd1 vssd1 vccd1 vccd1 _8062_/Q sky130_fd_sc_hd__dfxtp_1
X_4225_ _4225_/A _4225_/B vssd1 vssd1 vccd1 vccd1 _4225_/X sky130_fd_sc_hd__xor2_1
X_7013_ _7028_/A _7013_/B vssd1 vssd1 vccd1 vccd1 _7013_/X sky130_fd_sc_hd__and2_1
XFILLER_0_128_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4156_ _8516_/Q _4156_/B vssd1 vssd1 vccd1 vccd1 _4158_/C sky130_fd_sc_hd__xor2_1
XANTENNA__6863__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6630__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4087_ _6075_/A _6072_/A vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__or2_1
XANTENNA__7040__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5479__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7915_ _8465_/CLK _7915_/D vssd1 vssd1 vccd1 vccd1 _7915_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4867__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7846_ _8369_/CLK hold86/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4619__S1 _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5197__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7777_ _8478_/CLK _7777_/D vssd1 vssd1 vccd1 vccd1 _7777_/Q sky130_fd_sc_hd__dfxtp_1
X_4989_ _8196_/Q _8228_/Q _8292_/Q _7800_/Q _4990_/S0 _4990_/S1 vssd1 vssd1 vccd1
+ vccd1 _4989_/X sky130_fd_sc_hd__mux4_1
X_6728_ _6951_/A _6705_/B _6738_/B1 _6728_/B2 vssd1 vssd1 vccd1 vccd1 _6728_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4603__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6146__B1 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6659_ _6965_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6659_/X sky130_fd_sc_hd__and2_1
XFILLER_0_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1649_A _7344_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6697__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8329_ _8458_/CLK _8329_/D vssd1 vssd1 vccd1 vccd1 _8329_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4555__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout340 _3767_/X vssd1 vssd1 vccd1 vccd1 _6877_/A sky130_fd_sc_hd__buf_4
Xfanout384 _7050_/A vssd1 vssd1 vccd1 vccd1 _4737_/S1 sky130_fd_sc_hd__buf_4
Xfanout373 _5473_/A vssd1 vssd1 vccd1 vccd1 _4742_/S sky130_fd_sc_hd__buf_8
Xfanout351 _5726_/X vssd1 vssd1 vccd1 vccd1 _6414_/A2 sky130_fd_sc_hd__buf_4
Xfanout362 _3678_/X vssd1 vssd1 vccd1 vccd1 _4069_/S sky130_fd_sc_hd__clkbuf_16
Xfanout395 _7072_/B2 vssd1 vssd1 vccd1 vccd1 _4611_/S0 sky130_fd_sc_hd__buf_4
XANTENNA__3683__A1 _3682_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6013__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput26 i_instr_ID[5] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_2
Xinput15 i_instr_ID[24] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__buf_1
Xinput37 i_read_data_M[15] vssd1 vssd1 vccd1 vccd1 _6536_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput48 i_read_data_M[25] vssd1 vssd1 vccd1 vccd1 _6546_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6688__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput59 i_read_data_M[6] vssd1 vssd1 vccd1 vccd1 _6527_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4794__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4749__A _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5360__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6860__A1 _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4010_ _7979_/Q _4079_/A2 _4079_/B1 _8011_/Q _4009_/X vssd1 vssd1 vccd1 vccd1 _4010_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4484__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4849__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5299__B _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _5921_/A _5870_/A _5946_/A _5892_/A _5859_/S _5782_/S vssd1 vssd1 vccd1 vccd1
+ _5961_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6612__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7700_ _8388_/CLK _7700_/D vssd1 vssd1 vccd1 vccd1 _7700_/Q sky130_fd_sc_hd__dfxtp_1
X_4912_ _8185_/Q _8217_/Q _8281_/Q _7789_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4912_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_118_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5892_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5893_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7631_ _8362_/CLK _7631_/D vssd1 vssd1 vccd1 vccd1 _7631_/Q sky130_fd_sc_hd__dfxtp_1
X_4843_ _8465_/Q _8397_/Q _8429_/Q _8303_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4843_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3681__A_N _7282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4774_ _7026_/A _4774_/B vssd1 vssd1 vccd1 vccd1 _8131_/D sky130_fd_sc_hd__and2_1
XFILLER_0_55_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7562_ _8448_/CLK _7562_/D vssd1 vssd1 vccd1 vccd1 _7562_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3729__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7493_ _8481_/CLK _7493_/D vssd1 vssd1 vccd1 vccd1 _7493_/Q sky130_fd_sc_hd__dfxtp_1
X_3725_ _3725_/A _3725_/B vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__and2_1
XFILLER_0_16_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6513_ _6550_/A hold59/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__and2_1
XFILLER_0_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6679__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _8448_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_4_3_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6444_ _7022_/A _6444_/B vssd1 vssd1 vccd1 vccd1 _7926_/D sky130_fd_sc_hd__and2_1
XFILLER_0_130_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3656_ _7939_/Q vssd1 vssd1 vccd1 vccd1 _5581_/A sky130_fd_sc_hd__inv_2
XFILLER_0_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5351__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6375_ _6303_/X _6374_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6375_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8114_ _8114_/CLK _8114_/D vssd1 vssd1 vccd1 vccd1 _8114_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5481__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5326_ _6959_/A _5332_/A2 _5332_/B1 hold777/X vssd1 vssd1 vccd1 vccd1 _5326_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4537__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8045_ _8045_/CLK _8045_/D vssd1 vssd1 vccd1 vccd1 _8045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5257_ _6967_/A _5258_/A2 _5258_/B1 _5257_/B2 vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__a22o_1
X_4208_ _4208_/A _4209_/B vssd1 vssd1 vccd1 vccd1 _4208_/Y sky130_fd_sc_hd__nor2_1
X_5188_ _6741_/A _5188_/B vssd1 vssd1 vccd1 vccd1 _5188_/Y sky130_fd_sc_hd__nor2_1
X_4139_ _6334_/A _6331_/A vssd1 vssd1 vccd1 vccd1 _4139_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__5002__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7829_ _8160_/CLK _7829_/D vssd1 vssd1 vccd1 vccd1 _7829_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6114__A _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4333__S _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5590__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5953__A _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5342__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4776__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4528__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5645__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout192 _5772_/S vssd1 vssd1 vccd1 vccd1 _5782_/S sky130_fd_sc_hd__clkbuf_8
Xfanout181 _6251_/A vssd1 vssd1 vccd1 vccd1 _6163_/A sky130_fd_sc_hd__clkbuf_8
Xfanout170 _7030_/B vssd1 vssd1 vccd1 vccd1 _5540_/B sky130_fd_sc_hd__buf_2
XANTENNA__4508__S _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4751__B _4751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3648__A _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5030__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6959__A _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_752 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold618 _6774_/X vssd1 vssd1 vccd1 vccd1 _8325_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4490_ _5172_/A1 _4385_/B _5463_/C vssd1 vssd1 vccd1 vccd1 _7308_/D sky130_fd_sc_hd__mux2_1
Xhold607 _7451_/Q vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4479__A _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold629 _7483_/Q vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
X_6160_ _6140_/A _6157_/A _6096_/A _6115_/A _5782_/S _5859_/S vssd1 vssd1 vccd1 vccd1
+ _6160_/X sky130_fd_sc_hd__mux4_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5111_ _7078_/A _5523_/C vssd1 vssd1 vccd1 vccd1 _5111_/X sky130_fd_sc_hd__or2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ _4089_/B _6063_/A _6741_/A vssd1 vssd1 vccd1 vccd1 _6091_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5636__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5802__S _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6294__C1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1307 _6648_/X vssd1 vssd1 vccd1 vccd1 _8188_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1318 _8196_/Q vssd1 vssd1 vccd1 vccd1 _6664_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1329 _6658_/X vssd1 vssd1 vccd1 vccd1 _8193_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5042_ _5042_/A1 _4407_/B _5166_/B1 _5041_/X vssd1 vssd1 vccd1 vccd1 _7333_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_33_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5103__A _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6061__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6993_ _7065_/A _7067_/A _5547_/B _6992_/X vssd1 vssd1 vccd1 vccd1 _6993_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5944_ _5946_/A _5946_/B vssd1 vssd1 vccd1 vccd1 _5947_/A sky130_fd_sc_hd__and2_1
XFILLER_0_48_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5875_ _6126_/A _5952_/A _6362_/B vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4826_ _8140_/Q _7539_/Q _7411_/Q _7571_/Q _7063_/A _4976_/S1 vssd1 vssd1 vccd1 vccd1
+ _4826_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7614_ _8019_/CLK _7614_/D vssd1 vssd1 vccd1 vccd1 _7614_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7545_ _8339_/CLK _7545_/D vssd1 vssd1 vccd1 vccd1 _7545_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4757_ _7006_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _8114_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3708_ _4083_/B _3939_/B vssd1 vssd1 vccd1 vccd1 _3708_/Y sky130_fd_sc_hd__nor2_1
X_7476_ _8136_/CLK _7476_/D vssd1 vssd1 vccd1 vccd1 _7476_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4688_ _8350_/Q _7826_/Q _7492_/Q _7460_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4688_/X sky130_fd_sc_hd__mux4_1
X_6427_ _7008_/A _6427_/B vssd1 vssd1 vccd1 vccd1 _7909_/D sky130_fd_sc_hd__and2_1
XANTENNA__5492__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5324__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6358_ _6284_/X _6357_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6358_/X sky130_fd_sc_hd__mux2_1
X_5309_ _6925_/A _5332_/A2 _5332_/B1 hold421/X vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3886__A1 _3885_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5088__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5627__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5712__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6289_ _6279_/A _6281_/A _6288_/X vssd1 vssd1 vccd1 vccd1 _6292_/B sky130_fd_sc_hd__o21a_1
XANTENNA__6824__A1 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8028_ _8028_/CLK _8028_/D vssd1 vssd1 vccd1 vccd1 _8028_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4930__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6588__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4063__B2 _4057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4063__A1 _4756_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5012__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6760__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4998__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4997__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5683__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5315__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7068__A1 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3877__B2 _3875_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3877__A1 _4767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6579__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6961__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3990_ hold55/X _3676_/A _4082_/B1 _6853_/A _3989_/X vssd1 vssd1 vccd1 vccd1 _5892_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5251__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4762__A _7005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5660_ _6520_/A hold35/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__and2_1
XANTENNA__5069__S _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4611_ _8339_/Q _7815_/Q _7481_/Q _7449_/Q _4611_/S0 _4737_/S1 vssd1 vssd1 vccd1
+ vccd1 _4611_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_72_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6751__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5591_ _6853_/A _5584_/B _5617_/B1 hold503/X vssd1 vssd1 vccd1 vccd1 _5591_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_53_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4542_ _8136_/Q _7535_/Q _7407_/Q _7567_/Q _4611_/S0 _4640_/S1 vssd1 vssd1 vccd1
+ vccd1 _4542_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4701__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7330_ _8071_/CLK _7330_/D vssd1 vssd1 vccd1 vccd1 _7330_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold426 _6749_/X vssd1 vssd1 vccd1 vccd1 _8300_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7261_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7261_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5306__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 _7573_/Q vssd1 vssd1 vccd1 vccd1 hold415/X sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _7015_/A _7914_/Q vssd1 vssd1 vccd1 vccd1 _8046_/D sky130_fd_sc_hd__and2_1
Xhold404 _8141_/Q vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5857__A2 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold459 _8212_/Q vssd1 vssd1 vccd1 vccd1 hold459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _5206_/X vssd1 vssd1 vccd1 vccd1 _7420_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6391_/A _6212_/B vssd1 vssd1 vccd1 vccd1 _6212_/Y sky130_fd_sc_hd__nor2_1
Xhold437 _7822_/Q vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6143_ _6140_/A _6096_/A _6115_/A _6075_/A _5859_/S _5744_/S vssd1 vssd1 vccd1 vccd1
+ _6143_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_0_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6074_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6806__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1115 _8402_/Q vssd1 vssd1 vccd1 vccd1 _6872_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1104 _6583_/X vssd1 vssd1 vccd1 vccd1 _8155_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5609__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _5422_/A _5453_/C vssd1 vssd1 vccd1 vccd1 _5025_/X sky130_fd_sc_hd__or2_1
Xhold1137 _8340_/Q vssd1 vssd1 vccd1 vccd1 _6806_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7032__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1148 _6858_/X vssd1 vssd1 vccd1 vccd1 _8395_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _6950_/X vssd1 vssd1 vccd1 vccd1 _8440_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 _8161_/Q vssd1 vssd1 vccd1 vccd1 _6589_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4912__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6871__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout447_A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6976_ _6976_/A _6976_/B vssd1 vssd1 vccd1 vccd1 _6976_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5242__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5487__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6990__A0 _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5927_ _6008_/A _5926_/Y _5925_/X _6008_/B vssd1 vssd1 vccd1 vccd1 _5927_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5858_ _5856_/X _5857_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5858_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5789_ _5820_/A _5765_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5789_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5707__S _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4809_ _4808_/X _4807_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4809_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4979__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7528_ _7528_/CLK _7528_/D vssd1 vssd1 vccd1 vccd1 _7528_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1464_A _7305_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7459_ _8346_/CLK _7459_/D vssd1 vssd1 vccd1 vccd1 _7459_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1729_A _7358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold982 _6578_/X vssd1 vssd1 vccd1 vccd1 _8150_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold960 _5344_/X vssd1 vssd1 vccd1 vccd1 _7571_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold971 _8225_/Q vssd1 vssd1 vccd1 vccd1 hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold993 _8471_/Q vssd1 vssd1 vccd1 vccd1 _7013_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1660 _7690_/Q vssd1 vssd1 vccd1 vccd1 _3855_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4903__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1671 _7649_/Q vssd1 vssd1 vccd1 vccd1 _4285_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1682 _4212_/X vssd1 vssd1 vccd1 vccd1 _5559_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6781__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1693 _3967_/X vssd1 vssd1 vccd1 vccd1 _6425_/B sky130_fd_sc_hd__buf_1
XFILLER_0_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5678__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5233__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3795__B1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6733__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4757__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6830_ _7025_/A _6830_/A2 _6838_/A3 _6829_/X vssd1 vssd1 vccd1 vccd1 _6830_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5775__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6761_ _6945_/A _6773_/A2 _6773_/B1 hold853/X vssd1 vssd1 vccd1 vccd1 _6761_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3973_ _6251_/A _5870_/A vssd1 vssd1 vccd1 vccd1 _3973_/X sky130_fd_sc_hd__or2_1
X_8500_ _8500_/CLK hold91/X vssd1 vssd1 vccd1 vccd1 _8500_/Q sky130_fd_sc_hd__dfxtp_1
X_5712_ _6298_/A _6281_/A _5772_/S vssd1 vssd1 vccd1 vccd1 _5712_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6692_ _6951_/A _6669_/B _6702_/B1 hold685/X vssd1 vssd1 vccd1 vccd1 _6692_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_17_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6724__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5643_ _6951_/A _5620_/B _5653_/B1 hold497/X vssd1 vssd1 vccd1 vccd1 _5643_/X sky130_fd_sc_hd__a22o_1
X_8431_ _8431_/CLK _8431_/D vssd1 vssd1 vccd1 vccd1 _8431_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4431__S _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8362_ _8362_/CLK _8362_/D _7256_/Y vssd1 vssd1 vccd1 vccd1 _8362_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6212__A _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5574_ _7273_/A _5574_/B vssd1 vssd1 vccd1 vccd1 _7763_/D sky130_fd_sc_hd__nor2_1
X_4525_ _4524_/X _4523_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _4525_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7313_ _8360_/CLK _7313_/D _7123_/Y vssd1 vssd1 vccd1 vccd1 _7313_/Q sky130_fd_sc_hd__dfrtp_4
Xhold201 _5679_/X vssd1 vssd1 vccd1 vccd1 _7859_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 _8362_/Q vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
X_8293_ _8451_/CLK _8293_/D vssd1 vssd1 vccd1 vccd1 _8293_/Q sky130_fd_sc_hd__dfxtp_1
Xhold223 _5444_/X vssd1 vssd1 vccd1 vccd1 _7633_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _7316_/Q vssd1 vssd1 vccd1 vccd1 _5413_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold245 _5420_/X vssd1 vssd1 vccd1 vccd1 _7609_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _7735_/Q vssd1 vssd1 vccd1 vccd1 _5657_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold278 _7319_/Q vssd1 vssd1 vccd1 vccd1 _5416_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 _5054_/X vssd1 vssd1 vccd1 vccd1 _7339_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _7028_/A _7931_/Q vssd1 vssd1 vccd1 vccd1 _8063_/D sky130_fd_sc_hd__and2_1
XFILLER_0_1_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4387_ _4387_/A _4387_/B vssd1 vssd1 vccd1 vccd1 _4387_/Y sky130_fd_sc_hd__xnor2_1
Xhold289 _5435_/X vssd1 vssd1 vccd1 vccd1 _7624_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6126_ _6126_/A _6412_/S vssd1 vssd1 vccd1 vccd1 _6128_/B sky130_fd_sc_hd__nor2_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout397_A _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6255__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ _6057_/A _6057_/B vssd1 vssd1 vccd1 vccd1 _6058_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5008_ _4445_/A _5182_/A2 _5182_/B1 _5007_/X vssd1 vssd1 vccd1 vccd1 _7316_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4606__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_clk_A clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3765__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6959_ _6959_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6959_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_87_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6715__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_clk_A clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold790 _5365_/X vssd1 vssd1 vccd1 vccd1 _7592_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_3_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_3_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output114_A _7309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1490 _6457_/X vssd1 vssd1 vccd1 vccd1 _7939_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5206__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5757__A1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5852__S1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6182__A1 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6967__A _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5290_ _6961_/A _5294_/A2 _5294_/B1 hold563/X vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__a22o_1
X_4310_ _4310_/A _4310_/B vssd1 vssd1 vccd1 vccd1 _4310_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_23_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4241_ _4422_/A _4422_/B _4241_/C vssd1 vssd1 vccd1 vccd1 _4419_/A sky130_fd_sc_hd__and3_4
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4591__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4172_ _8514_/Q _4173_/B vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__or2_1
XANTENNA__6788__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7931_ _8476_/CLK _7931_/D vssd1 vssd1 vccd1 vccd1 _7931_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5111__A _7078_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6207__A _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7862_ _8033_/CLK hold80/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7793_ _8346_/CLK _7793_/D vssd1 vssd1 vccd1 vccd1 _7793_/Q sky130_fd_sc_hd__dfxtp_1
X_6813_ _6945_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6813_/X sky130_fd_sc_hd__and2_1
XFILLER_0_135_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6744_ _3939_/C _6742_/B _6742_/Y hold242/X vssd1 vssd1 vccd1 vccd1 _6744_/X sky130_fd_sc_hd__o22a_1
X_3956_ _4750_/B _3676_/A _4082_/B1 _6921_/A _3955_/X vssd1 vssd1 vccd1 vccd1 _5921_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_46_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6960__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6675_ _6917_/A _6701_/A2 _6701_/B1 hold691/X vssd1 vssd1 vccd1 vccd1 _6675_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_115_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5484__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3887_ _3887_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _3887_/X sky130_fd_sc_hd__or2_1
XANTENNA__7038__A _7077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8414_ _8483_/CLK _8414_/D vssd1 vssd1 vccd1 vccd1 _8414_/Q sky130_fd_sc_hd__dfxtp_1
X_5626_ _6917_/A _5652_/A2 _5652_/B1 hold589/X vssd1 vssd1 vccd1 vccd1 _5626_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout312_A _5260_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5557_ _6498_/A _5557_/B vssd1 vssd1 vccd1 vccd1 _7746_/D sky130_fd_sc_hd__and2_1
XANTENNA__6877__A _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8345_ _8448_/CLK _8345_/D vssd1 vssd1 vccd1 vccd1 _8345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3931__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5488_ _7509_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7677_/D sky130_fd_sc_hd__and3_1
X_4508_ _5136_/A1 _4508_/A1 _5449_/C vssd1 vssd1 vccd1 vccd1 _7290_/D sky130_fd_sc_hd__mux2_1
X_8276_ _8402_/CLK _8276_/D vssd1 vssd1 vccd1 vccd1 _8276_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4439_ _4435_/B _5442_/C _4438_/Y _4437_/X vssd1 vssd1 vccd1 vccd1 _8363_/D sky130_fd_sc_hd__a31o_1
X_7089_ _7052_/A _6975_/C _7069_/B _6554_/B _5073_/A vssd1 vssd1 vccd1 vccd1 _7089_/X
+ sky130_fd_sc_hd__o32a_1
X_6109_ _5734_/A _6098_/Y _6108_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6109_/Y sky130_fd_sc_hd__o22ai_1
XANTENNA__5720__S _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5987__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6164__A1 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7245__123 _8086_/CLK vssd1 vssd1 vccd1 vccd1 _8255_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__3923__B _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4573__S1 _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6219__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4790_ _8328_/Q _7804_/Q _7470_/Q _7438_/Q _4895_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4790_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3810_ _6388_/A _6386_/A vssd1 vssd1 vccd1 vccd1 _3811_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4770__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6942__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 _7309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3741_ _3741_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3672_ _7940_/Q _7667_/Q vssd1 vssd1 vccd1 vccd1 _3672_/Y sky130_fd_sc_hd__xnor2_1
X_6460_ _6494_/A _6460_/B vssd1 vssd1 vccd1 vccd1 _6460_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5411_ _5411_/A _7082_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5411_/X sky130_fd_sc_hd__and3_1
XFILLER_0_88_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6391_ _6391_/A _6391_/B vssd1 vssd1 vccd1 vccd1 _6391_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5902__A1 _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput114 _7309_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[27] sky130_fd_sc_hd__buf_12
XFILLER_0_113_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5342_ _6853_/A _5335_/B _5368_/B1 hold919/X vssd1 vssd1 vccd1 vccd1 _5342_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_88_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput125 _7290_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[8] sky130_fd_sc_hd__buf_12
XFILLER_0_70_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput103 _7298_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[16] sky130_fd_sc_hd__buf_12
X_8130_ _8130_/CLK _8130_/D vssd1 vssd1 vccd1 vccd1 _8130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput136 _8053_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[18] sky130_fd_sc_hd__buf_12
Xoutput158 _8044_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[9] sky130_fd_sc_hd__buf_12
X_8061_ _8061_/CLK _8061_/D vssd1 vssd1 vccd1 vccd1 _8061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput147 _8063_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[28] sky130_fd_sc_hd__buf_12
X_5273_ _6927_/A _5262_/B _5295_/B1 hold965/X vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__a22o_1
X_7012_ _7019_/A _7012_/B vssd1 vssd1 vccd1 vccd1 _7012_/X sky130_fd_sc_hd__and2_1
X_4224_ _4215_/Y _4219_/B _4224_/B1 vssd1 vssd1 vccd1 vccd1 _4225_/B sky130_fd_sc_hd__o21a_1
XANTENNA__5130__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4155_ _4155_/A1 _4154_/X _4155_/B1 vssd1 vssd1 vccd1 vccd1 _4155_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4086_ _6072_/A vssd1 vssd1 vccd1 vccd1 _4086_/Y sky130_fd_sc_hd__inv_2
XANTENNA__6091__B1 _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7040__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5479__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7914_ _8425_/CLK _7914_/D vssd1 vssd1 vccd1 vccd1 _7914_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout262_A _5262_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7845_ _8365_/CLK _7845_/D vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5197__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7776_ _8426_/CLK _7776_/D vssd1 vssd1 vccd1 vccd1 _7776_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5495__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4988_ _4986_/X _4987_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3939_ _4083_/B _3939_/B _3939_/C vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__and3b_1
X_7229__107 _8343_/CLK vssd1 vssd1 vccd1 vccd1 _8239_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_73_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6727_ _6949_/A _6737_/A2 _6737_/B1 hold969/X vssd1 vssd1 vccd1 vccd1 _6727_/X sky130_fd_sc_hd__a22o_1
X_6658_ _7024_/A _6658_/A2 _6605_/B _6657_/X vssd1 vssd1 vccd1 vccd1 _6658_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6697__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5609_ _6955_/A _5616_/A2 _5616_/B1 hold539/X vssd1 vssd1 vccd1 vccd1 _5609_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8328_ _8328_/CLK _8328_/D vssd1 vssd1 vccd1 vccd1 _8328_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3904__B1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5715__S _5716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6589_ _6965_/A _6559_/B _6591_/B1 _6589_/B2 vssd1 vssd1 vccd1 vccd1 _6589_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8259_ _8259_/CLK _8259_/D vssd1 vssd1 vccd1 vccd1 _8259_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4555__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout330 _6915_/A vssd1 vssd1 vccd1 vccd1 _6849_/A sky130_fd_sc_hd__clkbuf_8
Xfanout341 _3754_/X vssd1 vssd1 vccd1 vccd1 _6941_/A sky130_fd_sc_hd__buf_4
Xfanout374 _5473_/A vssd1 vssd1 vccd1 vccd1 _4641_/S sky130_fd_sc_hd__buf_4
Xfanout363 _3678_/X vssd1 vssd1 vccd1 vccd1 _4080_/S sky130_fd_sc_hd__buf_6
Xfanout352 _5726_/X vssd1 vssd1 vccd1 vccd1 _6105_/A2 sky130_fd_sc_hd__buf_4
Xfanout385 _7050_/A vssd1 vssd1 vccd1 vccd1 _5472_/A sky130_fd_sc_hd__clkbuf_8
Xfanout396 hold1641/X vssd1 vssd1 vccd1 vccd1 _7072_/B2 sky130_fd_sc_hd__buf_8
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5686__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3918__B _4161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6924__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput16 i_instr_ID[25] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 i_instr_ID[6] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput49 i_read_data_M[26] vssd1 vssd1 vccd1 vccd1 _6547_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__6688__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput38 i_read_data_M[16] vssd1 vssd1 vccd1 vccd1 _6537_/B sky130_fd_sc_hd__buf_1
XANTENNA__3934__A _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4794__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5360__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5648__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6456__S _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4765__A _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5960_ _6105_/A2 _5949_/A _5958_/X _6251_/A vssd1 vssd1 vccd1 vccd1 _5960_/X sky130_fd_sc_hd__a22o_1
X_5891_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4909_/X _4910_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7630_ _8363_/CLK _7630_/D vssd1 vssd1 vccd1 vccd1 _7630_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4704__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4842_ _8175_/Q _8207_/Q _8271_/Q _7779_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4842_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_23_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _6539_/A _4773_/B vssd1 vssd1 vccd1 vccd1 _8130_/D sky130_fd_sc_hd__and2_1
X_7561_ _8427_/CLK _7561_/D vssd1 vssd1 vccd1 vccd1 _7561_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7185__63 _7977_/CLK vssd1 vssd1 vccd1 vccd1 _8065_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3724_ _6318_/A _6315_/A vssd1 vssd1 vccd1 vccd1 _3725_/B sky130_fd_sc_hd__or2_1
X_6512_ _6545_/A hold53/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__and2_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7492_ _8160_/CLK _7492_/D vssd1 vssd1 vccd1 vccd1 _7492_/Q sky130_fd_sc_hd__dfxtp_1
X_6443_ _6999_/A _6443_/B vssd1 vssd1 vccd1 vccd1 _7925_/D sky130_fd_sc_hd__and2_1
XFILLER_0_130_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3655_ _7938_/Q vssd1 vssd1 vccd1 vccd1 _5222_/B sky130_fd_sc_hd__inv_2
XFILLER_0_113_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6679__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5351__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6374_ _6318_/A _6334_/A _6352_/A _6370_/A _5782_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6374_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8113_ _8113_/CLK _8113_/D vssd1 vssd1 vccd1 vccd1 _8113_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5325_ _6891_/A _5299_/B _5331_/B1 hold713/X vssd1 vssd1 vccd1 vccd1 _5325_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4537__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8044_ _8044_/CLK _8044_/D vssd1 vssd1 vccd1 vccd1 _8044_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5639__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5256_ _6965_/A _5258_/A2 _5258_/B1 hold701/X vssd1 vssd1 vccd1 vccd1 _5256_/X sky130_fd_sc_hd__a22o_1
X_4207_ _4432_/A _4432_/B vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__nand2b_1
X_5187_ _6908_/C _6558_/A vssd1 vssd1 vccd1 vccd1 _5189_/B sky130_fd_sc_hd__or2_1
XANTENNA__6064__A0 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4138_ _4138_/A _4138_/B vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4394__B _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4069_ _8082_/Q _4068_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _4069_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6906__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7828_ _8353_/CLK _7828_/D vssd1 vssd1 vccd1 vccd1 _7828_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7759_ _8504_/CLK _7759_/D vssd1 vssd1 vccd1 vccd1 _7759_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1661_A _3855_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1759_A _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5590__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4776__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5342__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6130__A _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4528__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout160 _5370_/Y vssd1 vssd1 vccd1 vccd1 _7090_/A sky130_fd_sc_hd__buf_4
Xfanout182 _3970_/X vssd1 vssd1 vccd1 vccd1 _6251_/A sky130_fd_sc_hd__buf_4
Xfanout171 _7030_/B vssd1 vssd1 vccd1 vccd1 _5465_/B sky130_fd_sc_hd__buf_4
XFILLER_0_135_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout193 _3928_/X vssd1 vssd1 vccd1 vccd1 _5772_/S sky130_fd_sc_hd__buf_6
XFILLER_0_89_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3849__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6305__A _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_121_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6959__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold608 _5243_/X vssd1 vssd1 vccd1 vccd1 _7451_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold619 _8304_/Q vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4136__A3 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6975__A _7356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5884__A3 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6090_ _5734_/A _6078_/X _6089_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _6090_/X sky130_fd_sc_hd__a2bb2o_1
X_5110_ input16/X _5069_/S _5182_/B1 _5109_/X vssd1 vssd1 vccd1 vccd1 _7367_/D sky130_fd_sc_hd__o211a_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _5430_/A _5456_/C vssd1 vssd1 vccd1 vccd1 _5041_/X sky130_fd_sc_hd__or2_1
XFILLER_0_109_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1319 _6664_/X vssd1 vssd1 vccd1 vccd1 _8196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1308 _8443_/Q vssd1 vssd1 vccd1 vccd1 _6956_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5103__B _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6992_ _8529_/Z _5388_/X _6976_/B vssd1 vssd1 vccd1 vccd1 _6992_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_87_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5943_ _5943_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _5946_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5874_ _6393_/A _5874_/B vssd1 vssd1 vccd1 vccd1 _6362_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4825_ _8333_/Q _7809_/Q _7475_/Q _7443_/Q _4983_/S0 _4976_/S1 vssd1 vssd1 vccd1
+ vccd1 _4825_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7613_ _8019_/CLK _7613_/D vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7544_ _8338_/CLK _7544_/D vssd1 vssd1 vccd1 vccd1 _7544_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4756_ _7006_/A _4756_/B vssd1 vssd1 vccd1 vccd1 _8113_/D sky130_fd_sc_hd__and2_1
XANTENNA__6869__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_A _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3707_ _4769_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__and2_1
X_7475_ _8478_/CLK _7475_/D vssd1 vssd1 vccd1 vccd1 _7475_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7046__A _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4687_ _4686_/X _4683_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7523_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5492__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6426_ _7015_/A _6426_/B vssd1 vssd1 vccd1 vccd1 _7908_/D sky130_fd_sc_hd__and2_1
XANTENNA__5324__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4389__B _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6885__A _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6357_ _6298_/A _6318_/A _6334_/A _6352_/A _5782_/S _5804_/A vssd1 vssd1 vccd1 vccd1
+ _6357_/X sky130_fd_sc_hd__mux4_1
X_5308_ _6923_/A _5299_/B _5331_/B1 _5308_/B2 vssd1 vssd1 vccd1 vccd1 _5308_/X sky130_fd_sc_hd__a22o_1
X_6288_ _3736_/Y _6414_/A2 _6398_/B1 _6279_/A _6414_/B1 vssd1 vssd1 vccd1 vccd1 _6288_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4609__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1820 _7883_/Q vssd1 vssd1 vccd1 vccd1 hold1820/X sky130_fd_sc_hd__dlygate4sd3_1
X_5239_ _6931_/A _5258_/A2 _5258_/B1 hold649/X vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__a22o_1
X_8027_ _8090_/CLK _8027_/D vssd1 vssd1 vccd1 vccd1 _8027_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4930__S1 _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6588__A1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4063__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_415 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6779__B _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6760__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4997__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5315__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6795__A _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3877__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6276__B1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__buf_1
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6579__A1 _6945_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5251__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4685__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6035__A _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4254__S _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4610_ _4609_/X _4606_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7512_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5874__A _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6751__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7155__33 _7903_/CLK vssd1 vssd1 vccd1 vccd1 _8035_/CLK sky130_fd_sc_hd__inv_2
X_5590_ _6917_/A _5616_/A2 _5616_/B1 hold727/X vssd1 vssd1 vccd1 vccd1 _5590_/X sky130_fd_sc_hd__a22o_1
X_4541_ _8329_/Q _7805_/Q _7471_/Q _7439_/Q _4611_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4541_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_80_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold427 _8272_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5306__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold416 _5346_/X vssd1 vssd1 vccd1 vccd1 _7573_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4472_ _7007_/A _7915_/Q vssd1 vssd1 vccd1 vccd1 _8047_/D sky130_fd_sc_hd__and2_1
X_7260_ _7264_/A vssd1 vssd1 vccd1 vccd1 _7260_/Y sky130_fd_sc_hd__inv_2
Xhold405 _6569_/X vssd1 vssd1 vccd1 vccd1 _8141_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5857__A3 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6211_ _6211_/A _6211_/B vssd1 vssd1 vccd1 vccd1 _6212_/B sky130_fd_sc_hd__xnor2_1
Xhold438 _5642_/X vssd1 vssd1 vccd1 vccd1 _7822_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _7460_/Q vssd1 vssd1 vccd1 vccd1 hold449/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6142_ _6142_/A _6142_/B vssd1 vssd1 vccd1 vccd1 _6142_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6267__B1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ _6075_/A _6075_/B vssd1 vssd1 vccd1 vccd1 _6076_/A sky130_fd_sc_hd__and2_1
XANTENNA__3841__B _3841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1105 _7792_/Q vssd1 vssd1 vccd1 vccd1 _5608_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5024_/A1 _4425_/B _5148_/B1 _5023_/X vssd1 vssd1 vccd1 vccd1 _7324_/D sky130_fd_sc_hd__o211a_1
Xhold1138 _6806_/X vssd1 vssd1 vccd1 vccd1 _8340_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 _6872_/X vssd1 vssd1 vccd1 vccd1 _8402_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1149 _8446_/Q vssd1 vssd1 vccd1 vccd1 _6962_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1127 _8411_/Q vssd1 vssd1 vccd1 vccd1 _6890_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4912__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A hold1510/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _7356_/Q _7348_/Q _6975_/C vssd1 vssd1 vccd1 vccd1 _6976_/B sky130_fd_sc_hd__and3_1
XANTENNA__5242__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5487__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5926_ _5952_/A _5926_/B vssd1 vssd1 vccd1 vccd1 _5926_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout342_A _3740_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5857_ _5946_/A _5974_/A _5993_/A _6016_/A _5744_/S _5859_/S vssd1 vssd1 vccd1 vccd1
+ _5857_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_63_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5788_ _6911_/A _5788_/B vssd1 vssd1 vccd1 vccd1 _7869_/D sky130_fd_sc_hd__nor2_1
X_4808_ _8460_/Q _8392_/Q _8424_/Q _8298_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4808_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4979__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4739_ _4737_/X _4738_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__mux2_1
X_7527_ _7527_/CLK _7527_/D vssd1 vssd1 vccd1 vccd1 _7527_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7458_ _8484_/CLK _7458_/D vssd1 vssd1 vccd1 vccd1 _7458_/Q sky130_fd_sc_hd__dfxtp_1
X_6409_ _6388_/A _6352_/A _6126_/A _6370_/A _5859_/S _5782_/S vssd1 vssd1 vccd1 vccd1
+ _6409_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold961 _7819_/Q vssd1 vssd1 vccd1 vccd1 hold961/X sky130_fd_sc_hd__dlygate4sd3_1
X_7389_ _8504_/CLK _7389_/D vssd1 vssd1 vccd1 vccd1 _7389_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4600__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold972 _6698_/X vssd1 vssd1 vccd1 vccd1 _8225_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold950 _5327_/X vssd1 vssd1 vccd1 vccd1 _7558_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 _8487_/Q vssd1 vssd1 vccd1 vccd1 _7029_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 _7013_/X vssd1 vssd1 vccd1 vccd1 _8471_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8527__475 vssd1 vssd1 vccd1 vccd1 _8527_/A _8527__475/LO sky130_fd_sc_hd__conb_1
Xhold1661 _3855_/X vssd1 vssd1 vccd1 vccd1 _6443_/B sky130_fd_sc_hd__buf_1
Xhold1650 _7055_/B vssd1 vssd1 vccd1 vccd1 _7046_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__4903__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1694 _7674_/Q vssd1 vssd1 vccd1 vccd1 _3958_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1672 _4285_/Y vssd1 vssd1 vccd1 vccd1 _4286_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1683 _7686_/Q vssd1 vssd1 vccd1 vccd1 _3783_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5233__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4667__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4074__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3795__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4802__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6733__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4757__B _4757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output69_A _8115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5869__A _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4773__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6760_ _6877_/A _6741_/B _6774_/B1 hold643/X vssd1 vssd1 vccd1 vccd1 _6760_/X sky130_fd_sc_hd__a22o_1
X_5711_ _5707_/X _5710_/X _5952_/A vssd1 vssd1 vccd1 vccd1 _5711_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6972__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3972_ _4748_/B _3676_/A _4082_/B1 _3965_/X _3971_/X vssd1 vssd1 vccd1 vccd1 _5870_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_122_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5808__S _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6691_ _6949_/A _6701_/A2 _6701_/B1 hold475/X vssd1 vssd1 vccd1 vccd1 _6691_/X sky130_fd_sc_hd__a22o_1
X_8430_ _8462_/CLK _8430_/D vssd1 vssd1 vccd1 vccd1 _8430_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6724__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5642_ _6949_/A _5652_/A2 _5652_/B1 hold437/X vssd1 vssd1 vccd1 vccd1 _5642_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_127_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7128__6 _8461_/CLK vssd1 vssd1 vccd1 vccd1 _7505_/CLK sky130_fd_sc_hd__inv_2
X_8361_ _8361_/CLK _8361_/D _7255_/Y vssd1 vssd1 vccd1 vccd1 _8361_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5573_ _6551_/A _5573_/B vssd1 vssd1 vccd1 vccd1 _7762_/D sky130_fd_sc_hd__and2_1
XFILLER_0_26_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4524_ _8456_/Q _8388_/Q _8420_/Q _8294_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4524_/X sky130_fd_sc_hd__mux4_1
X_7312_ _8030_/CLK _7312_/D _7122_/Y vssd1 vssd1 vccd1 vccd1 _7312_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold202 _7616_/Q vssd1 vssd1 vccd1 vccd1 _5674_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _7802_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _5012_/X vssd1 vssd1 vccd1 vccd1 _7318_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _5413_/X vssd1 vssd1 vccd1 vccd1 _7602_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8292_ _8450_/CLK _8292_/D vssd1 vssd1 vccd1 vccd1 _8292_/Q sky130_fd_sc_hd__dfxtp_1
Xhold257 _5657_/X vssd1 vssd1 vccd1 vccd1 _7837_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 _7565_/Q vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _7375_/Q vssd1 vssd1 vccd1 vccd1 _5442_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4455_ _7024_/A _7932_/Q vssd1 vssd1 vccd1 vccd1 _8064_/D sky130_fd_sc_hd__and2_1
Xhold279 _5416_/X vssd1 vssd1 vccd1 vccd1 _7605_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5160__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4386_ _5052_/A1 _4385_/X _5456_/C vssd1 vssd1 vccd1 vccd1 _8382_/D sky130_fd_sc_hd__mux2_1
X_6125_ _6414_/A2 _6119_/A _6123_/X _5739_/Y _6124_/X vssd1 vssd1 vccd1 vccd1 _6125_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3710__A1 _3709_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout292_A _6667_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6056_/A _6056_/B vssd1 vssd1 vccd1 vccd1 _6057_/B sky130_fd_sc_hd__or2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _5413_/A _7030_/C vssd1 vssd1 vccd1 vccd1 _5007_/X sky130_fd_sc_hd__or2_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5498__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4018__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5215__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4649__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6958_ _7022_/A _6958_/A2 _6970_/A3 _6957_/X vssd1 vssd1 vccd1 vccd1 _6958_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_91_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5909_ _5745_/X _5783_/X _6144_/S vssd1 vssd1 vccd1 vccd1 _5909_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_64_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6889_ _6955_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6889_/X sky130_fd_sc_hd__and2_1
XFILLER_0_133_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6715__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4821__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold780 _5602_/X vssd1 vssd1 vccd1 vccd1 _7786_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 _7490_/Q vssd1 vssd1 vccd1 vccd1 hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4069__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4888__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1480 _7043_/Y vssd1 vssd1 vccd1 vccd1 _8494_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1491 _7310_/Q vssd1 vssd1 vccd1 vccd1 _5176_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5206__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output107_A _7302_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6954__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4532__S _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4812__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6032__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap355_A _6406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6967__B _6969_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4768__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5142__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4240_ _5563_/B hold637/X _5453_/B vssd1 vssd1 vccd1 vccd1 _4241_/C sky130_fd_sc_hd__mux2_1
X_4171_ _4164_/Y _4171_/B vssd1 vssd1 vccd1 vccd1 _4171_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_117_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4707__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7930_ _8010_/CLK _7930_/D vssd1 vssd1 vccd1 vccd1 _7930_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7861_ _8385_/CLK _7861_/D vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5111__B _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6812_ _7007_/A _6812_/A2 _6779_/B _6811_/X vssd1 vssd1 vccd1 vccd1 _6812_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7792_ _8442_/CLK _7792_/D vssd1 vssd1 vccd1 vccd1 _7792_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6743_ _6777_/A _6742_/B _6742_/Y hold298/X vssd1 vssd1 vccd1 vccd1 _6743_/X sky130_fd_sc_hd__o22a_1
X_3955_ _7706_/Q _4081_/B vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6674_ _6849_/A _6669_/B _6702_/B1 hold529/X vssd1 vssd1 vccd1 vccd1 _6674_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4420__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5625_ _6849_/A _5621_/B _5621_/Y hold276/X vssd1 vssd1 vccd1 vccd1 _5625_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_115_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3886_ _8088_/Q _3885_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8413_ _8413_/CLK _8413_/D vssd1 vssd1 vccd1 vccd1 _8413_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7038__B _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6877__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5556_ _6494_/A _5556_/B vssd1 vssd1 vccd1 vccd1 _7745_/D sky130_fd_sc_hd__and2_1
XFILLER_0_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout305_A _5582_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8344_ _8346_/CLK _8344_/D vssd1 vssd1 vccd1 vccd1 _8344_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3931__B2 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4507_ _5138_/A1 _4432_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _7291_/D sky130_fd_sc_hd__mux2_1
X_5487_ _7508_/Q _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7676_/D sky130_fd_sc_hd__and3_1
X_8275_ _8473_/CLK _8275_/D vssd1 vssd1 vccd1 vccd1 _8275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4438_ _4440_/A _4193_/B _4193_/C vssd1 vssd1 vccd1 vccd1 _4438_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6330__C1 _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4369_ _6419_/B _4370_/B _6418_/B vssd1 vssd1 vccd1 vccd1 _4369_/Y sky130_fd_sc_hd__nor3b_1
XANTENNA__6893__A _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7088_ _7088_/A _7088_/B _7088_/C vssd1 vssd1 vccd1 vccd1 _8518_/D sky130_fd_sc_hd__and3_1
X_6108_ _5952_/A _5926_/B _6309_/B _6107_/Y _6128_/A vssd1 vssd1 vccd1 vccd1 _6108_/X
+ sky130_fd_sc_hd__o32a_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4617__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6039_ _6016_/A _5974_/A _6035_/A _5993_/A _5859_/S _5782_/S vssd1 vssd1 vccd1 vccd1
+ _6039_/X sky130_fd_sc_hd__mux4_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6936__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__B _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3757__A _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_115_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8010_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4411__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5972__A _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6787__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5124__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3686__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4770__B _4770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_19 _7289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3740_ _8094_/Q _3739_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4402__A2 _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8355_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3671_ _7937_/Q _3659_/Y _3661_/Y _7939_/Q _3670_/Y vssd1 vssd1 vccd1 vccd1 _3675_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5410_ _6553_/B _7069_/B _6973_/C _7079_/B vssd1 vssd1 vccd1 vccd1 _7599_/D sky130_fd_sc_hd__o31a_1
X_6390_ _6390_/A _6390_/B vssd1 vssd1 vccd1 vccd1 _6391_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5363__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3913__A1 _3912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_71_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput104 _7299_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[17] sky130_fd_sc_hd__buf_12
XFILLER_0_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput115 _7310_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[28] sky130_fd_sc_hd__buf_12
XFILLER_0_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5341_ _6917_/A _5367_/A2 _5367_/B1 _5341_/B2 vssd1 vssd1 vccd1 vccd1 _5341_/X sky130_fd_sc_hd__a22o_1
Xoutput126 _7291_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[9] sky130_fd_sc_hd__buf_12
XFILLER_0_121_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput137 _8054_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[19] sky130_fd_sc_hd__buf_12
XFILLER_0_50_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput148 _8064_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[29] sky130_fd_sc_hd__buf_12
X_8060_ _8060_/CLK _8060_/D vssd1 vssd1 vccd1 vccd1 _8060_/Q sky130_fd_sc_hd__dfxtp_1
X_5272_ _6925_/A _5262_/B _5295_/B1 hold781/X vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__a22o_1
X_7011_ _7029_/A _7011_/B vssd1 vssd1 vccd1 vccd1 _7011_/X sky130_fd_sc_hd__and2_1
XFILLER_0_11_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4223_ _4221_/Y _4223_/B vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4154_ _4143_/X _4144_/Y _4153_/Y _4152_/A _4152_/Y vssd1 vssd1 vccd1 vccd1 _4154_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_86_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4085_ _4085_/A0 _4084_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _6072_/A sky130_fd_sc_hd__mux2_2
X_7913_ _8011_/CLK _7913_/D vssd1 vssd1 vccd1 vccd1 _7913_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6630__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7844_ _8365_/CLK _7844_/D vssd1 vssd1 vccd1 vccd1 _7844_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6918__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A _5584_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7775_ _8425_/CLK _7775_/D vssd1 vssd1 vccd1 vccd1 _7775_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_24_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5495__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6726_ _6947_/A _6737_/A2 _6737_/B1 _6726_/B2 vssd1 vssd1 vccd1 vccd1 _6726_/X sky130_fd_sc_hd__a22o_1
X_4987_ _8163_/Q _7562_/Q _7434_/Q _7594_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4987_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_19_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3938_ _3939_/C vssd1 vssd1 vccd1 vccd1 _6845_/A sky130_fd_sc_hd__inv_2
XANTENNA_fanout422_A _7357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6657_ _6963_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6657_/X sky130_fd_sc_hd__and2_1
XFILLER_0_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3869_ _4764_/B _4071_/A2 _4071_/B1 _3862_/X _3868_/X vssd1 vssd1 vccd1 vccd1 _6209_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5354__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4900__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8530__471 vssd1 vssd1 vccd1 vccd1 _8530__471/HI _8530_/A sky130_fd_sc_hd__conb_1
XANTENNA__4157__A1 _8517_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_2_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_2_0_clk/X sky130_fd_sc_hd__clkbuf_8
X_5608_ _6953_/A _5616_/A2 _5616_/B1 _5608_/B2 vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__a22o_1
X_6588_ _6963_/A _6559_/B _6591_/B1 hold455/X vssd1 vssd1 vccd1 vccd1 _6588_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_39_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8327_ _8421_/CLK _8327_/D vssd1 vssd1 vccd1 vccd1 _8327_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3904__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5539_ _8258_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7728_/D sky130_fd_sc_hd__and3_1
XFILLER_0_42_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5106__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8258_ _8258_/CLK _8258_/D vssd1 vssd1 vccd1 vccd1 _8258_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout320 _4048_/X vssd1 vssd1 vccd1 vccd1 _6937_/A sky130_fd_sc_hd__buf_4
Xfanout331 _3886_/X vssd1 vssd1 vccd1 vccd1 _6951_/A sky130_fd_sc_hd__buf_4
X_8189_ _8479_/CLK _8189_/D vssd1 vssd1 vccd1 vccd1 _8189_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout375 hold1637/X vssd1 vssd1 vccd1 vccd1 _5473_/A sky130_fd_sc_hd__buf_6
Xfanout353 _5723_/X vssd1 vssd1 vccd1 vccd1 _6405_/B sky130_fd_sc_hd__buf_8
Xfanout364 _3657_/Y vssd1 vssd1 vccd1 vccd1 _4074_/S sky130_fd_sc_hd__buf_8
Xfanout342 _3740_/X vssd1 vssd1 vccd1 vccd1 _6963_/A sky130_fd_sc_hd__buf_4
Xfanout386 hold1633/X vssd1 vssd1 vccd1 vccd1 _7050_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__4347__S _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout397 _7057_/A vssd1 vssd1 vccd1 vccd1 _4999_/S sky130_fd_sc_hd__buf_8
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4093__B1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5593__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 i_instr_ID[26] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_1
Xinput28 i_instr_ID[7] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__buf_2
XFILLER_0_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5345__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput39 i_read_data_M[17] vssd1 vssd1 vccd1 vccd1 _6538_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA__4810__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5648__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6860__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3950__A _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6612__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5890_ _5892_/A _5892_/B vssd1 vssd1 vccd1 vccd1 _5893_/A sky130_fd_sc_hd__and2_1
X_4910_ _8152_/Q _7551_/Q _7423_/Q _7583_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4910_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_114_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _4839_/X _4840_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4841_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_87_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4772_ _6520_/A _4772_/B vssd1 vssd1 vccd1 vccd1 _8129_/D sky130_fd_sc_hd__and2_1
X_7560_ _8419_/CLK _7560_/D vssd1 vssd1 vccd1 vccd1 _7560_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3723_ _3723_/A _6315_/A vssd1 vssd1 vccd1 vccd1 _3725_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7491_ _8346_/CLK _7491_/D vssd1 vssd1 vccd1 vccd1 _7491_/Q sky130_fd_sc_hd__dfxtp_1
X_6511_ _6550_/A hold21/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__and2_1
X_3654_ _7937_/Q vssd1 vssd1 vccd1 vccd1 _5296_/A sky130_fd_sc_hd__inv_2
XFILLER_0_113_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6501__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6442_ _7028_/A _6442_/B vssd1 vssd1 vccd1 vccd1 _7924_/D sky130_fd_sc_hd__and2_1
XFILLER_0_130_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5887__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3844__B _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8112_ _8112_/CLK _8112_/D vssd1 vssd1 vccd1 vccd1 _8112_/Q sky130_fd_sc_hd__dfxtp_2
X_6373_ _6380_/B _6373_/B vssd1 vssd1 vccd1 vccd1 _6373_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5117__A _7075_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5639__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5324_ _6955_/A _5299_/B _5331_/B1 hold901/X vssd1 vssd1 vccd1 vccd1 _5324_/X sky130_fd_sc_hd__a22o_1
X_8043_ _8043_/CLK _8043_/D vssd1 vssd1 vccd1 vccd1 _8043_/Q sky130_fd_sc_hd__dfxtp_1
X_5255_ _6963_/A _5258_/A2 _5258_/B1 hold453/X vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__a22o_1
X_4206_ _5558_/B _5018_/A1 _5453_/B vssd1 vssd1 vccd1 vccd1 _4432_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5186_ _6908_/C _6558_/A vssd1 vssd1 vccd1 vccd1 _5186_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__6064__A1 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4137_ _3750_/B _4136_/X _4135_/Y vssd1 vssd1 vccd1 vccd1 _4138_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout372_A hold1637/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4068_ _7986_/Q _4068_/A2 _4068_/B1 _8018_/Q _4067_/X vssd1 vssd1 vccd1 vccd1 _4068_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_78_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7827_ _8451_/CLK _7827_/D vssd1 vssd1 vccd1 vccd1 _7827_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_7758_ _8020_/CLK _7758_/D vssd1 vssd1 vccd1 vccd1 _7758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6709_ _6847_/A _6706_/B _6706_/Y hold226/X vssd1 vssd1 vccd1 vccd1 _6709_/X sky130_fd_sc_hd__o22a_1
X_7689_ _8481_/CLK _7689_/D vssd1 vssd1 vccd1 vccd1 _7689_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5327__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4630__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3770__A _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 _6307_/A vssd1 vssd1 vccd1 vccd1 _6412_/S sky130_fd_sc_hd__clkbuf_8
Xfanout172 _7030_/B vssd1 vssd1 vccd1 vccd1 _5470_/B sky130_fd_sc_hd__buf_4
Xfanout161 _5182_/B1 vssd1 vssd1 vccd1 vccd1 _5166_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout194 _5950_/S vssd1 vssd1 vccd1 vccd1 _5952_/A sky130_fd_sc_hd__buf_4
XFILLER_0_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5030__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5318__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4540__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold609 _7427_/Q vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output99_A _7294_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5040_/A1 _5067_/S _5172_/B1 _5039_/X vssd1 vssd1 vccd1 vccd1 _7332_/D sky130_fd_sc_hd__o211a_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1309 _6956_/X vssd1 vssd1 vccd1 vccd1 _8443_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6046__A1 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6991__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6046__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6991_ _7090_/A _6991_/B vssd1 vssd1 vccd1 vccd1 _8454_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_125_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5942_ _3962_/B _6011_/A2 _5933_/Y _5941_/X _6911_/A vssd1 vssd1 vccd1 vccd1 _5942_/Y
+ sky130_fd_sc_hd__a221oi_2
XANTENNA__4715__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5873_ _5710_/X _5714_/X _5950_/S vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4824_ _4823_/X _4820_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8236_/D sky130_fd_sc_hd__mux2_1
X_7612_ _8034_/CLK _7612_/D vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4755_ _7026_/A _4755_/B vssd1 vssd1 vccd1 vccd1 _8112_/D sky130_fd_sc_hd__and2_1
X_7543_ _8467_/CLK _7543_/D vssd1 vssd1 vccd1 vccd1 _7543_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3706_ _4083_/B _3941_/B vssd1 vssd1 vccd1 vccd1 _3706_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5309__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7474_ _8426_/CLK _7474_/D vssd1 vssd1 vccd1 vccd1 _7474_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout218_A _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4686_ _4685_/X _4684_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__mux2_1
X_6425_ _6999_/A _6425_/B vssd1 vssd1 vccd1 vccd1 _7907_/D sky130_fd_sc_hd__and2_1
XANTENNA__6885__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6356_ _6354_/Y _6355_/X _6391_/A vssd1 vssd1 vccd1 vccd1 _6356_/X sky130_fd_sc_hd__o21ba_1
X_5307_ _6921_/A _5332_/A2 _5332_/B1 hold865/X vssd1 vssd1 vccd1 vccd1 _5307_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5088__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6287_ _5740_/Y _5984_/Y _6286_/X _6251_/A vssd1 vssd1 vccd1 vccd1 _6287_/X sky130_fd_sc_hd__o2bb2a_1
X_8026_ _8090_/CLK _8026_/D vssd1 vssd1 vccd1 vccd1 _8026_/Q sky130_fd_sc_hd__dfxtp_1
X_5238_ _6929_/A _5226_/B _5259_/B1 hold517/X vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__a22o_1
Xhold1810 _7893_/Q vssd1 vssd1 vccd1 vccd1 hold1810/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6824__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1821 _7630_/Q vssd1 vssd1 vccd1 vccd1 hold1821/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_95_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _8485_/CLK sky130_fd_sc_hd__clkbuf_16
X_5169_ _5464_/A _5465_/C vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__or2_1
XANTENNA__6588__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5012__A2 _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_427 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6760__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6795__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_86_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _7903_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4039__B1 _4035_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6579__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6316__A _6318_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5251__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4685__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6200__B2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6751__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4540_ _4539_/X _4536_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7502_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_10_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _8484_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold406 _8306_/Q vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _8204_/Q vssd1 vssd1 vccd1 vccd1 hold417/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4471_ _7028_/A _7916_/Q vssd1 vssd1 vccd1 vccd1 _8048_/D sky130_fd_sc_hd__and2_1
Xhold439 _8274_/Q vssd1 vssd1 vccd1 vccd1 hold439/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 _6717_/X vssd1 vssd1 vccd1 vccd1 _8272_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5890__A _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6210_ _6210_/A _6210_/B vssd1 vssd1 vccd1 vccd1 _6211_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7170__48 _8010_/CLK vssd1 vssd1 vccd1 vccd1 _8050_/CLK sky130_fd_sc_hd__inv_2
X_6141_ _6141_/A _6141_/B vssd1 vssd1 vccd1 vccd1 _6142_/B sky130_fd_sc_hd__nand2_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ _6072_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6075_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__6806__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1106 _5608_/X vssd1 vssd1 vccd1 vccd1 _7792_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1139 _8426_/Q vssd1 vssd1 vccd1 vccd1 _6922_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1117 _8166_/Q vssd1 vssd1 vccd1 vccd1 _6604_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _5421_/A _5451_/C vssd1 vssd1 vccd1 vccd1 _5023_/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_77_clk clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 _8387_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1128 _6890_/X vssd1 vssd1 vccd1 vccd1 _8411_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6974_ _6974_/A _6981_/B vssd1 vssd1 vccd1 vccd1 _6990_/S sky130_fd_sc_hd__or2_1
XANTENNA__5242__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout168_A hold1510/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6226__A _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5925_ _6270_/A _5925_/B vssd1 vssd1 vccd1 vccd1 _5925_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5856_ _5846_/A _5870_/A _5892_/A _5921_/A _5744_/S _5859_/S vssd1 vssd1 vccd1 vccd1
+ _5856_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout335_A _3826_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4807_ _8170_/Q _8202_/Q _8266_/Q _7774_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4807_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_133_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5787_ _5762_/Y _5775_/X _5786_/X _6011_/A2 _3951_/Y vssd1 vssd1 vccd1 vccd1 _5787_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__7057__A _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4738_ _8164_/Q _7563_/Q _7435_/Q _7595_/Q _4741_/S0 _7050_/A vssd1 vssd1 vccd1 vccd1
+ _4738_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7526_ _7526_/CLK _7526_/D vssd1 vssd1 vccd1 vccd1 _7526_/Q sky130_fd_sc_hd__dfxtp_1
X_4669_ _4667_/X _4668_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4669_/X sky130_fd_sc_hd__mux2_1
X_7457_ _8402_/CLK _7457_/D vssd1 vssd1 vccd1 vccd1 _7457_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6408_ _6402_/Y _6404_/X _6406_/Y _6407_/X _5734_/A vssd1 vssd1 vccd1 vccd1 _6408_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_4_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold940 _6767_/X vssd1 vssd1 vccd1 vccd1 _8318_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold951 _8468_/Q vssd1 vssd1 vccd1 vccd1 _7010_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold962 _5639_/X vssd1 vssd1 vccd1 vccd1 _7819_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4600__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold973 _8289_/Q vssd1 vssd1 vccd1 vccd1 hold973/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7388_ _8195_/CLK _7388_/D vssd1 vssd1 vccd1 vccd1 _7388_/Q sky130_fd_sc_hd__dfxtp_1
Xhold995 _7549_/Q vssd1 vssd1 vccd1 vccd1 hold995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 _7029_/X vssd1 vssd1 vccd1 vccd1 _8487_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ _6337_/Y _6338_/X _6391_/A vssd1 vssd1 vccd1 vccd1 _6339_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_hold1617_A _3981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8009_ _8477_/CLK _8009_/D vssd1 vssd1 vccd1 vccd1 _8009_/Q sky130_fd_sc_hd__dfxtp_2
Xhold1651 _7678_/Q vssd1 vssd1 vccd1 vccd1 _4004_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1640 _4183_/Y vssd1 vssd1 vccd1 vccd1 _5555_/B sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_68_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _8361_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1662 _7679_/Q vssd1 vssd1 vccd1 vccd1 _4028_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1695 _3958_/X vssd1 vssd1 vccd1 vccd1 _6427_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1684 _3783_/X vssd1 vssd1 vccd1 vccd1 _6439_/B sky130_fd_sc_hd__buf_1
Xhold1673 _4286_/Y vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5233__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4667__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3795__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6733__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_59_clk clkbuf_4_15_0_clk/X vssd1 vssd1 vccd1 vccd1 _8011_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4773__B _4773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3971_ _3971_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _3971_/X sky130_fd_sc_hd__or2_1
X_5710_ _5708_/X _5709_/X _5838_/A vssd1 vssd1 vccd1 vccd1 _5710_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7215__93 _8382_/CLK vssd1 vssd1 vccd1 vccd1 _8128_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_15_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6690_ _6947_/A _6701_/A2 _6701_/B1 hold587/X vssd1 vssd1 vccd1 vccd1 _6690_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6724__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5641_ _6947_/A _5652_/A2 _5652_/B1 hold889/X vssd1 vssd1 vccd1 vccd1 _5641_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5932__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8360_ _8360_/CLK _8360_/D _7254_/Y vssd1 vssd1 vccd1 vccd1 _8360_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5572_ _7273_/A _5572_/B vssd1 vssd1 vccd1 vccd1 _7761_/D sky130_fd_sc_hd__nor2_1
X_4523_ _8166_/Q _8198_/Q _8262_/Q _7770_/Q _7362_/Q _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4523_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5109__B _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7311_ _8385_/CLK _7311_/D _7121_/Y vssd1 vssd1 vccd1 vccd1 _7311_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8291_ _8350_/CLK _8291_/D vssd1 vssd1 vccd1 vccd1 _8291_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold225 _5622_/X vssd1 vssd1 vccd1 vccd1 _7802_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _7376_/Q vssd1 vssd1 vccd1 vccd1 _5443_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _5674_/X vssd1 vssd1 vccd1 vccd1 _7854_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _5338_/X vssd1 vssd1 vccd1 vccd1 _7565_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold258 _7566_/Q vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _6498_/A _7933_/Q vssd1 vssd1 vccd1 vccd1 _8065_/D sky130_fd_sc_hd__and2_1
Xhold269 _5442_/X vssd1 vssd1 vccd1 vccd1 _7631_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3852__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold236 _7857_/Q vssd1 vssd1 vccd1 vccd1 _6478_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4594__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4385_ _4385_/A _4385_/B vssd1 vssd1 vccd1 vccd1 _4385_/X sky130_fd_sc_hd__xor2_1
X_6124_ _4077_/A _6414_/B1 _6398_/B1 _6112_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6124_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6056_/A _6056_/B vssd1 vssd1 vccd1 vccd1 _6055_/Y sky130_fd_sc_hd__nor2_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _4448_/A _4448_/B _5140_/B1 _5005_/X vssd1 vssd1 vccd1 vccd1 _7315_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6660__A1 _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout285_A _6775_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout452_A _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6099__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5498__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5215__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4649__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6957_ _6957_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6957_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5908_ _5777_/X _5780_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5908_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6888_ _7026_/A _6888_/A2 _6906_/A3 _6887_/X vssd1 vssd1 vccd1 vccd1 _6888_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6715__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6403__B _6406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5839_ _6393_/A _5952_/B _5836_/A vssd1 vssd1 vccd1 vccd1 _5840_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4821__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7509_ _7509_/CLK _7509_/D vssd1 vssd1 vccd1 vccd1 _7509_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8489_ _8500_/CLK _8489_/D vssd1 vssd1 vccd1 vccd1 _8489_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold781 _7476_/Q vssd1 vssd1 vccd1 vccd1 hold781/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3762__B _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold770 _5366_/X vssd1 vssd1 vccd1 vccd1 _7593_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _5286_/X vssd1 vssd1 vccd1 vccd1 _7490_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4888__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1470 _7300_/Q vssd1 vssd1 vccd1 vccd1 _5156_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4085__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold1492 _7309_/Q vssd1 vssd1 vccd1 vccd1 _5174_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 _7299_/Q vssd1 vssd1 vccd1 vccd1 _5154_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5206__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4813__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6167__B1 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4812__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output81_A _8126_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7140__18 _8339_/CLK vssd1 vssd1 vccd1 vccd1 _7517_/CLK sky130_fd_sc_hd__inv_2
X_4170_ _5553_/B _4445_/A _7030_/B vssd1 vssd1 vccd1 vccd1 _4171_/B sky130_fd_sc_hd__mux2_1
XANTENNA__6890__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6642__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7130__8 _8173_/CLK vssd1 vssd1 vccd1 vccd1 _7507_/CLK sky130_fd_sc_hd__inv_2
X_7860_ _8032_/CLK _7860_/D vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6811_ _6877_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6811_/X sky130_fd_sc_hd__and2_1
X_7791_ _8283_/CLK _7791_/D vssd1 vssd1 vccd1 vccd1 _7791_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6742_ _6999_/A _6742_/B vssd1 vssd1 vccd1 vccd1 _6742_/Y sky130_fd_sc_hd__nand2_1
X_3954_ _8073_/Q _3953_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _3954_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6673_ _6847_/A _6670_/B _6670_/Y hold252/X vssd1 vssd1 vccd1 vccd1 _6673_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6223__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3885_ _7992_/Q _4079_/A2 _4079_/B1 _8024_/Q _3884_/X vssd1 vssd1 vccd1 vccd1 _3885_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5624_ _6847_/A _5620_/B _5653_/B1 hold695/X vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__a22o_1
X_8412_ _8480_/CLK _8412_/D vssd1 vssd1 vccd1 vccd1 _8412_/Q sky130_fd_sc_hd__dfxtp_1
X_8343_ _8343_/CLK _8343_/D vssd1 vssd1 vccd1 vccd1 _8343_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5555_ _6494_/A _5555_/B vssd1 vssd1 vccd1 vccd1 _7744_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8274_ _8466_/CLK _8274_/D vssd1 vssd1 vccd1 vccd1 _8274_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3931__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4506_ _5140_/A1 _4430_/B _5449_/C vssd1 vssd1 vccd1 vccd1 _7292_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5486_ _7507_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7675_/D sky130_fd_sc_hd__and3_1
X_4437_ _4437_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4437_/X sky130_fd_sc_hd__and2_1
XANTENNA__7054__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4368_ _4361_/X _4362_/Y _4367_/X vssd1 vssd1 vccd1 vccd1 _4370_/B sky130_fd_sc_hd__o21a_1
XANTENNA__6893__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6107_ _6008_/A _5928_/Y _5955_/Y vssd1 vssd1 vccd1 vccd1 _6107_/Y sky130_fd_sc_hd__a21oi_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7087_ _5544_/A _6975_/C _7080_/X _7050_/A vssd1 vssd1 vccd1 vccd1 _7088_/C sky130_fd_sc_hd__a22o_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _8496_/Q _4299_/B vssd1 vssd1 vccd1 vccd1 _4299_/Y sky130_fd_sc_hd__nand2_1
X_6038_ _6038_/A _6038_/B vssd1 vssd1 vccd1 vccd1 _6038_/X sky130_fd_sc_hd__xor2_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold1684_A _3783_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7989_ _8071_/CLK _7989_/D vssd1 vssd1 vccd1 vccd1 _7989_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3757__B _3757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4558__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6872__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3686__B2 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6624__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4730__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4543__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5060__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3670_ _7938_/Q _7665_/Q vssd1 vssd1 vccd1 vccd1 _3670_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4797__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5363__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput105 _7300_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[18] sky130_fd_sc_hd__buf_12
X_5340_ _6849_/A _5336_/B _5336_/Y hold290/X vssd1 vssd1 vccd1 vccd1 _5340_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_112_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput116 _7311_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[29] sky130_fd_sc_hd__buf_12
XFILLER_0_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5271_ _6923_/A _5294_/A2 _5294_/B1 _5271_/B2 vssd1 vssd1 vccd1 vccd1 _5271_/X sky130_fd_sc_hd__a22o_1
Xoutput138 _8036_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[1] sky130_fd_sc_hd__buf_12
Xoutput127 _8035_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[0] sky130_fd_sc_hd__buf_12
Xoutput149 _8037_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[2] sky130_fd_sc_hd__buf_12
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4549__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7010_ _7010_/A _7010_/B vssd1 vssd1 vccd1 vccd1 _7010_/X sky130_fd_sc_hd__and2_1
X_4222_ _8507_/Q _4222_/B vssd1 vssd1 vccd1 vccd1 _4222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_128_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4153_ _4153_/A _5690_/A vssd1 vssd1 vccd1 vccd1 _4153_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4718__S _4735_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5403__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4084_ _4084_/A1 _4084_/A2 _6935_/A _4084_/B2 _4083_/X vssd1 vssd1 vccd1 vccd1 _4084_/X
+ sky130_fd_sc_hd__a221o_2
X_7912_ _8426_/CLK _7912_/D vssd1 vssd1 vccd1 vccd1 _7912_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6091__A2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7843_ _8363_/CLK _7843_/D vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__6379__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3858__A _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4986_ _8356_/Q _7832_/Q _7498_/Q _7466_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4986_/X sky130_fd_sc_hd__mux4_1
X_7774_ _8350_/CLK _7774_/D vssd1 vssd1 vccd1 vccd1 _7774_/Q sky130_fd_sc_hd__dfxtp_1
X_3937_ _8068_/Q _3677_/Y _4079_/B1 _8004_/Q _3936_/X vssd1 vssd1 vccd1 vccd1 _3939_/C
+ sky130_fd_sc_hd__a221o_4
XANTENNA_fanout248_A _6705_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6725_ _6945_/A _6737_/A2 _6737_/B1 hold625/X vssd1 vssd1 vccd1 vccd1 _6725_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_A _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6656_ _7024_/A _6656_/A2 _6666_/A3 _6655_/X vssd1 vssd1 vccd1 vccd1 _6656_/X sky130_fd_sc_hd__a31o_1
X_3868_ _3868_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3868_/X sky130_fd_sc_hd__or2_1
XANTENNA__5354__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5607_ _6951_/A _5584_/B _5617_/B1 hold683/X vssd1 vssd1 vccd1 vccd1 _5607_/X sky130_fd_sc_hd__a22o_1
X_3799_ _3799_/A _3799_/B vssd1 vssd1 vccd1 vccd1 _3800_/D sky130_fd_sc_hd__and2_1
X_6587_ _6961_/A _6559_/B _6591_/B1 hold921/X vssd1 vssd1 vccd1 vccd1 _6587_/X sky130_fd_sc_hd__a22o_1
X_8326_ _8326_/CLK _8326_/D vssd1 vssd1 vccd1 vccd1 _8326_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7065__A _7065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3904__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5538_ _8257_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7727_/D sky130_fd_sc_hd__and3_1
XANTENNA__6303__A0 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8257_ _8257_/CLK _8257_/D vssd1 vssd1 vccd1 vccd1 _8257_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6854__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5469_ _5469_/A _5470_/B _7030_/C vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__and3_1
Xfanout310 _5297_/Y vssd1 vssd1 vccd1 vccd1 _5332_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_111_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout321 _4035_/X vssd1 vssd1 vccd1 vccd1 _6927_/A sky130_fd_sc_hd__buf_4
Xfanout332 _3875_/X vssd1 vssd1 vccd1 vccd1 _6955_/A sky130_fd_sc_hd__buf_4
X_8188_ _8442_/CLK _8188_/D vssd1 vssd1 vccd1 vccd1 _8188_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout365 _3657_/Y vssd1 vssd1 vccd1 vccd1 _4085_/S sky130_fd_sc_hd__buf_4
Xfanout354 _5723_/X vssd1 vssd1 vccd1 vccd1 _6094_/B sky130_fd_sc_hd__clkbuf_8
Xfanout343 _6957_/A vssd1 vssd1 vccd1 vccd1 _6891_/A sky130_fd_sc_hd__buf_4
XANTENNA__6606__A1 _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 _7057_/A vssd1 vssd1 vccd1 vccd1 _4929_/S sky130_fd_sc_hd__buf_8
XFILLER_0_94_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6067__C1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout387 _4720_/S0 vssd1 vssd1 vccd1 vccd1 _4706_/S0 sky130_fd_sc_hd__buf_8
Xfanout376 _4741_/S1 vssd1 vssd1 vccd1 vccd1 _4733_/S1 sky130_fd_sc_hd__clkbuf_8
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4093__A1 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4712__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5290__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3840__A1 _6452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5593__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5042__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 i_instr_ID[27] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput29 i_instr_ID[8] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4779__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5345__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5648__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4951__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5281__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4084__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4703__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4840_ _8142_/Q _7541_/Q _7413_/Q _7573_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4840_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6054__A _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3678__A _7282_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6510_ _7005_/A _6510_/B vssd1 vssd1 vccd1 vccd1 _6510_/X sky130_fd_sc_hd__and2_1
X_4771_ _6551_/A _4771_/B vssd1 vssd1 vccd1 vccd1 _8128_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3722_ _3722_/A0 _6447_/B _4074_/S vssd1 vssd1 vccd1 vccd1 _6315_/A sky130_fd_sc_hd__mux2_2
X_7490_ _8484_/CLK _7490_/D vssd1 vssd1 vccd1 vccd1 _7490_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3653_ _7835_/Q vssd1 vssd1 vccd1 vccd1 _3653_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6441_ _7267_/A _6441_/B vssd1 vssd1 vccd1 vccd1 _7923_/D sky130_fd_sc_hd__nor2_2
X_6372_ _6355_/A _6355_/B _6353_/A vssd1 vssd1 vccd1 vccd1 _6373_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_24_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8111_ _8111_/CLK _8111_/D vssd1 vssd1 vccd1 vccd1 _8111_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__7089__A1 _7052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5323_ _6953_/A _5299_/B _5331_/B1 hold693/X vssd1 vssd1 vccd1 vccd1 _5323_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5117__B _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5639__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8042_ _8042_/CLK _8042_/D vssd1 vssd1 vccd1 vccd1 _8042_/Q sky130_fd_sc_hd__dfxtp_1
X_5254_ _6961_/A _5258_/A2 _5258_/B1 hold549/X vssd1 vssd1 vccd1 vccd1 _5254_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6836__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5185_ _7939_/Q _7940_/Q vssd1 vssd1 vccd1 vccd1 _6558_/A sky130_fd_sc_hd__nand2_4
X_4205_ _4205_/A _4205_/B vssd1 vssd1 vccd1 vccd1 _4205_/X sky130_fd_sc_hd__xor2_1
XANTENNA_fanout198_A _6393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4136_ _3750_/A _3733_/Y _6281_/A _3711_/Y _6298_/A vssd1 vssd1 vccd1 vccd1 _4136_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6064__A2 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5272__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _3657_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7235__113 _8467_/CLK vssd1 vssd1 vccd1 vccd1 _8245_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4067_ _4067_/A_N _7954_/Q vssd1 vssd1 vccd1 vccd1 _4067_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7826_ _8350_/CLK _7826_/D vssd1 vssd1 vccd1 vccd1 _7826_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5024__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6899__A _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4969_ _8483_/Q _8415_/Q _8447_/Q _8321_/Q _4983_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4969_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6772__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7757_ _8373_/CLK _7757_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
X_6708_ _3939_/C _6706_/B _6706_/Y hold262/X vssd1 vssd1 vccd1 vccd1 _6708_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7176__54 _8471_/CLK vssd1 vssd1 vccd1 vccd1 _8056_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__4911__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7688_ _8442_/CLK _7688_/D vssd1 vssd1 vccd1 vccd1 _7688_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5327__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6639_ _6945_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6639_/X sky130_fd_sc_hd__and2_1
XFILLER_0_34_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8309_ _8471_/CLK _8309_/D vssd1 vssd1 vccd1 vccd1 _8309_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6288__C1 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4358__S _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6139__A _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout173 hold1510/X vssd1 vssd1 vccd1 vccd1 _7030_/B sky130_fd_sc_hd__clkbuf_4
Xfanout162 _5182_/B1 vssd1 vssd1 vccd1 vccd1 _5172_/B1 sky130_fd_sc_hd__buf_4
XANTENNA__4933__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 _5879_/S vssd1 vssd1 vccd1 vccd1 _5950_/S sky130_fd_sc_hd__clkbuf_4
Xfanout184 _6307_/A vssd1 vssd1 vccd1 vccd1 _6198_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_70_clk_A clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__B2 _8031_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6763__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_85_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5318__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3961__A _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6818__A1 _6434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4268__S _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4924__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3900__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6990_ _7074_/A _6989_/Y _6990_/S vssd1 vssd1 vccd1 vccd1 _6991_/B sky130_fd_sc_hd__mux2_1
Xclkbuf_4_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_1_0_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_38_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _5734_/A _5923_/Y _5940_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _5941_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5254__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5872_ _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5872_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5006__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4823_ _4822_/X _4821_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__mux2_1
X_7611_ _8034_/CLK _7611_/D vssd1 vssd1 vccd1 vccd1 _7611_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6754__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4754_ _7006_/A _4754_/B vssd1 vssd1 vccd1 vccd1 _8111_/D sky130_fd_sc_hd__and2_1
X_7542_ _8143_/CLK _7542_/D vssd1 vssd1 vccd1 vccd1 _7542_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3705_ _3705_/A _3705_/B _3705_/C _3705_/D vssd1 vssd1 vccd1 vccd1 _3941_/B sky130_fd_sc_hd__or4_1
XANTENNA__5309__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7473_ _8425_/CLK _7473_/D vssd1 vssd1 vccd1 vccd1 _7473_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4685_ _8479_/Q _8411_/Q _8443_/Q _8317_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4685_/X sky130_fd_sc_hd__mux4_1
X_6424_ _6741_/A _6424_/B vssd1 vssd1 vccd1 vccd1 _7906_/D sky130_fd_sc_hd__nor2_1
X_6355_ _6355_/A _6355_/B _6355_/C vssd1 vssd1 vccd1 vccd1 _6355_/X sky130_fd_sc_hd__and3_1
X_5306_ _6853_/A _5332_/A2 _5332_/B1 hold783/X vssd1 vssd1 vccd1 vccd1 _5306_/X sky130_fd_sc_hd__a22o_1
X_6286_ _6144_/X _6285_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6286_/X sky130_fd_sc_hd__mux2_1
X_5237_ _6927_/A _5226_/B _5259_/B1 hold545/X vssd1 vssd1 vccd1 vccd1 _5237_/X sky130_fd_sc_hd__a22o_1
X_8025_ _8090_/CLK _8025_/D vssd1 vssd1 vccd1 vccd1 _8025_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1811 _7894_/Q vssd1 vssd1 vccd1 vccd1 hold1811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1800 _8373_/Q vssd1 vssd1 vccd1 vccd1 hold1800/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1822 _7353_/Q vssd1 vssd1 vccd1 vccd1 hold1822/X sky130_fd_sc_hd__dlygate4sd3_1
X_5168_ _5168_/A1 _5067_/S _5172_/B1 _5167_/X vssd1 vssd1 vccd1 vccd1 _7396_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4048__A1 _4047_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4119_ _6388_/A _6386_/A vssd1 vssd1 vccd1 vccd1 _4119_/Y sky130_fd_sc_hd__nand2b_1
X_5099_ _7052_/A _5099_/B vssd1 vssd1 vccd1 vccd1 _5099_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5245__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6406__B _6406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6745__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7809_ _8478_/CLK _7809_/D vssd1 vssd1 vccd1 vccd1 _7809_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4641__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5720__A1 _5719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7253__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4906__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4816__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5236__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4039__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6984__A0 _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5882__S1 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6736__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6332__A _6334_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold407 _6755_/X vssd1 vssd1 vccd1 vccd1 _8306_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _6677_/X vssd1 vssd1 vccd1 vccd1 _8204_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4470_ _7018_/A _7917_/Q vssd1 vssd1 vccd1 vccd1 _8049_/D sky130_fd_sc_hd__and2_1
XFILLER_0_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold429 _7457_/Q vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6140_ _6140_/A _6140_/B vssd1 vssd1 vccd1 vccd1 _6141_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ _4066_/B _6063_/A _6063_/Y _6070_/X _6741_/A vssd1 vssd1 vccd1 vccd1 _6071_/Y
+ sky130_fd_sc_hd__a221oi_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1129 _8422_/Q vssd1 vssd1 vccd1 vccd1 _6914_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 _6604_/X vssd1 vssd1 vccd1 vccd1 _8166_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5022_ _5022_/A1 _5144_/A2 _5146_/B1 _5021_/X vssd1 vssd1 vccd1 vccd1 _7323_/D sky130_fd_sc_hd__o211a_1
Xhold1107 _7449_/Q vssd1 vssd1 vccd1 vccd1 _5241_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6507__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6973_ _7090_/A _6973_/B _6973_/C vssd1 vssd1 vccd1 vccd1 _8452_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_88_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5924_ _5803_/B _5808_/X _6393_/A vssd1 vssd1 vccd1 vccd1 _5925_/B sky130_fd_sc_hd__mux2_1
X_5855_ _6105_/A2 _5850_/A _5853_/X _5739_/Y vssd1 vssd1 vccd1 vccd1 _5855_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6727__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout230_A _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4806_ _4804_/X _4805_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_106_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5786_ _6163_/A _5786_/B _5785_/X vssd1 vssd1 vccd1 vccd1 _5786_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7057__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7146__24 _8486_/CLK vssd1 vssd1 vccd1 vccd1 _7523_/CLK sky130_fd_sc_hd__inv_2
X_4737_ _8357_/Q _7833_/Q _7499_/Q _7467_/Q _4741_/S0 _4737_/S1 vssd1 vssd1 vccd1
+ vccd1 _4737_/X sky130_fd_sc_hd__mux4_1
X_7525_ _7525_/CLK _7525_/D vssd1 vssd1 vccd1 vccd1 _7525_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4668_ _8154_/Q _7553_/Q _7425_/Q _7585_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4668_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7456_ _8440_/CLK _7456_/D vssd1 vssd1 vccd1 vccd1 _7456_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6407_ _6390_/A _6387_/X _6403_/Y _6405_/Y _6389_/B vssd1 vssd1 vccd1 vccd1 _6407_/X
+ sky130_fd_sc_hd__o221a_1
Xhold930 _5593_/X vssd1 vssd1 vccd1 vccd1 _7777_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 _7010_/X vssd1 vssd1 vccd1 vccd1 _8468_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _8139_/Q vssd1 vssd1 vccd1 vccd1 hold941/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7073__A _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold963 _8163_/Q vssd1 vssd1 vccd1 vccd1 hold963/X sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _4597_/X _4598_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4599_/X sky130_fd_sc_hd__mux2_1
X_7387_ _8485_/CLK _7387_/D vssd1 vssd1 vccd1 vccd1 _7387_/Q sky130_fd_sc_hd__dfxtp_1
Xhold996 _5318_/X vssd1 vssd1 vccd1 vccd1 _7549_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 _7560_/Q vssd1 vssd1 vccd1 vccd1 hold985/X sky130_fd_sc_hd__dlygate4sd3_1
X_6338_ _6338_/A _6338_/B vssd1 vssd1 vccd1 vccd1 _6338_/X sky130_fd_sc_hd__or2_1
XFILLER_0_8_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold974 _6734_/X vssd1 vssd1 vccd1 vccd1 _8289_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1512_A _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6269_ _6195_/X _6268_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6270_/B sky130_fd_sc_hd__mux2_1
X_8008_ _8008_/CLK _8008_/D vssd1 vssd1 vccd1 vccd1 _8008_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1652 _4004_/X vssd1 vssd1 vccd1 vccd1 _6431_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1641 _7362_/Q vssd1 vssd1 vccd1 vccd1 hold1641/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold1630 _8501_/Q vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__buf_1
Xhold1663 _4028_/X vssd1 vssd1 vccd1 vccd1 _6432_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5218__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1696 _8498_/Q vssd1 vssd1 vccd1 vccd1 _3891_/A0 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1674 _4288_/X vssd1 vssd1 vccd1 vccd1 _5570_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1685 _8504_/Q vssd1 vssd1 vccd1 vccd1 _4074_/A0 sky130_fd_sc_hd__buf_1
XFILLER_0_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6718__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3776__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5991__A _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5941__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5941__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4546__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5209__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _4074_/S _3967_/X _3968_/X vssd1 vssd1 vccd1 vccd1 _3970_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6972__A3 _6908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _6945_/A _5652_/A2 _5652_/B1 hold400/X vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_26_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5571_ _7027_/A _5571_/B vssd1 vssd1 vccd1 vccd1 _7760_/D sky130_fd_sc_hd__and2_1
X_4522_ _4520_/X _4521_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _4522_/X sky130_fd_sc_hd__mux2_1
X_8290_ _8319_/CLK _8290_/D vssd1 vssd1 vccd1 vccd1 _8290_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7310_ _8385_/CLK _7310_/D _7120_/Y vssd1 vssd1 vccd1 vccd1 _7310_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold226 _8264_/Q vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 _5443_/X vssd1 vssd1 vccd1 vccd1 _7632_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _7022_/A _7934_/Q vssd1 vssd1 vccd1 vccd1 _8066_/D sky130_fd_sc_hd__and2_1
Xhold204 _7332_/Q vssd1 vssd1 vccd1 vccd1 _5429_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold259 _5339_/X vssd1 vssd1 vccd1 vccd1 _7566_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _7380_/Q vssd1 vssd1 vccd1 vccd1 _5447_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5696__A0 _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold237 _6478_/X vssd1 vssd1 vccd1 vccd1 _7960_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4594__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4384_ _4334_/Y _5468_/C _4383_/X _4382_/X vssd1 vssd1 vccd1 vccd1 _8383_/D sky130_fd_sc_hd__a31o_1
XANTENNA__5160__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6123_ _5962_/X _6122_/X _6411_/S vssd1 vssd1 vccd1 vccd1 _6123_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6056_/A _6056_/B vssd1 vssd1 vccd1 vccd1 _6057_/A sky130_fd_sc_hd__nand2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5412_/A _5442_/C vssd1 vssd1 vccd1 vccd1 _5005_/X sky130_fd_sc_hd__or2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout278_A _6971_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout180_A _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6099__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout445_A _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6956_ _7018_/A _6956_/A2 _6970_/A3 _6955_/X vssd1 vssd1 vccd1 vccd1 _6956_/X sky130_fd_sc_hd__a31o_1
X_5907_ _6144_/S _5797_/S _5773_/C _5906_/Y vssd1 vssd1 vccd1 vccd1 _5907_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_119_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4191__S _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6887_ _6953_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6887_/X sky130_fd_sc_hd__and2_1
XFILLER_0_106_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5838_ _5838_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _5952_/B sky130_fd_sc_hd__or2_1
XFILLER_0_48_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5769_ _5769_/A _5769_/B vssd1 vssd1 vccd1 vccd1 _5769_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7508_ _7508_/CLK _7508_/D vssd1 vssd1 vccd1 vccd1 _7508_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_121_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8488_ _8500_/CLK _8488_/D vssd1 vssd1 vccd1 vccd1 _8488_/Q sky130_fd_sc_hd__dfxtp_1
X_7439_ _8458_/CLK _7439_/D vssd1 vssd1 vccd1 vccd1 _7439_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold782 _5272_/X vssd1 vssd1 vccd1 vccd1 _7476_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 _5215_/X vssd1 vssd1 vccd1 vccd1 _7429_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 _8290_/Q vssd1 vssd1 vccd1 vccd1 hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold793 _8284_/Q vssd1 vssd1 vccd1 vccd1 hold793/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1460 _8363_/Q vssd1 vssd1 vccd1 vccd1 _4437_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold1482 _7733_/Q vssd1 vssd1 vccd1 vccd1 _5655_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 _7313_/Q vssd1 vssd1 vccd1 vccd1 _5182_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1471 _7898_/Q vssd1 vssd1 vccd1 vccd1 _4774_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_67_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5611__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6954__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6167__A1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5226__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5142__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4576__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output74_A _8120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6810_ _7017_/A _6810_/A2 _6838_/A3 _6809_/X vssd1 vssd1 vccd1 vccd1 _6810_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7790_ _8440_/CLK _7790_/D vssd1 vssd1 vccd1 vccd1 _7790_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5602__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6741_ _6741_/A _6741_/B vssd1 vssd1 vccd1 vccd1 _6741_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3953_ _7977_/Q _4079_/A2 _4079_/B1 _8009_/Q _3952_/X vssd1 vssd1 vccd1 vccd1 _3953_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6672_ _3939_/C _6669_/B _6702_/B1 hold469/X vssd1 vssd1 vccd1 vccd1 _6672_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _7283_/Q _7960_/Q vssd1 vssd1 vccd1 vccd1 _3884_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_18_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5623_ _3939_/C _5620_/B _5653_/B1 hold443/X vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8411_ _8479_/CLK _8411_/D vssd1 vssd1 vccd1 vccd1 _8411_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6520__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8342_ _8445_/CLK _8342_/D vssd1 vssd1 vccd1 vccd1 _8342_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5554_ _6494_/A _5554_/B vssd1 vssd1 vccd1 vccd1 _7743_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4505_ _5142_/A1 _4505_/A1 _7088_/B vssd1 vssd1 vccd1 vccd1 _7293_/D sky130_fd_sc_hd__mux2_1
X_5485_ _7506_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7674_/D sky130_fd_sc_hd__and3_1
X_8273_ _8431_/CLK _8273_/D vssd1 vssd1 vccd1 vccd1 _8273_/Q sky130_fd_sc_hd__dfxtp_1
X_4436_ _4432_/A _5449_/C _4435_/Y _4434_/X vssd1 vssd1 vccd1 vccd1 _8364_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_41_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4367_ _4367_/A _4367_/B _4367_/C _4367_/D vssd1 vssd1 vccd1 vccd1 _4367_/X sky130_fd_sc_hd__or4_1
XANTENNA_fanout395_A _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6106_ _6094_/A _5732_/X _6063_/A _6104_/X _6105_/X vssd1 vssd1 vccd1 vccd1 _6106_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7086_ _7088_/A _7088_/B _7086_/C vssd1 vssd1 vccd1 vccd1 _8517_/D sky130_fd_sc_hd__and3_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _8496_/Q _4299_/B vssd1 vssd1 vccd1 vccd1 _4298_/Y sky130_fd_sc_hd__nor2_1
X_6037_ _6018_/A _6017_/A _6015_/Y vssd1 vssd1 vccd1 vccd1 _6038_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_96_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4914__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6936__A3 _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7988_ _8020_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 _7988_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6939_ _6939_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6939_/X sky130_fd_sc_hd__and2_1
XANTENNA__6149__B2 _5719_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6430__A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4558__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5124__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold590 _5626_/X vssd1 vssd1 vccd1 vccd1 _7806_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7261__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3686__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4824__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1290 _8191_/Q vssd1 vssd1 vccd1 vccd1 _6654_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4730__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7200__78 _8079_/CLK vssd1 vssd1 vccd1 vccd1 _8113_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_82_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4797__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5363__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput106 _7301_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[19] sky130_fd_sc_hd__buf_12
XFILLER_0_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput128 _8045_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[10] sky130_fd_sc_hd__buf_12
X_5270_ _6921_/A _5262_/B _5295_/B1 hold787/X vssd1 vssd1 vccd1 vccd1 _5270_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6312__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput139 _8055_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[20] sky130_fd_sc_hd__buf_12
Xoutput117 _7284_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[2] sky130_fd_sc_hd__buf_12
XFILLER_0_121_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4221_ _4221_/A _4222_/B vssd1 vssd1 vccd1 vccd1 _4221_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5746__S0 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4549__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ _4152_/A _5733_/C vssd1 vssd1 vccd1 vccd1 _4152_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_37_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4083_ _4757_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _4083_/X sky130_fd_sc_hd__and2_1
X_7911_ _8283_/CLK _7911_/D vssd1 vssd1 vccd1 vccd1 _7911_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4019__B _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7842_ _7977_/CLK _7842_/D vssd1 vssd1 vccd1 vccd1 _7842_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6918__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6515__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7773_ _8338_/CLK _7773_/D vssd1 vssd1 vccd1 vccd1 _7773_/Q sky130_fd_sc_hd__dfxtp_1
X_4985_ _4984_/X _4981_/X _7057_/A vssd1 vssd1 vccd1 vccd1 _8259_/D sky130_fd_sc_hd__mux2_1
X_3936_ _7282_/Q _7283_/Q _7972_/Q vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6724_ _6877_/A _6705_/B _6738_/B1 _6724_/B2 vssd1 vssd1 vccd1 vccd1 _6724_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_129_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3867_ _3968_/A _6441_/B _3865_/Y vssd1 vssd1 vccd1 vccd1 _3871_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6655_ _6961_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6655_/X sky130_fd_sc_hd__and2_1
XFILLER_0_27_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5354__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6586_ _6959_/A _6592_/A2 _6592_/B1 hold386/X vssd1 vssd1 vccd1 vccd1 _6586_/X sky130_fd_sc_hd__a22o_1
X_3798_ _6191_/A _6188_/A vssd1 vssd1 vccd1 vccd1 _3799_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout408_A _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5606_ _6949_/A _5616_/A2 _5616_/B1 hold465/X vssd1 vssd1 vccd1 vccd1 _5606_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_131_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7065__B _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8325_ _8487_/CLK _8325_/D vssd1 vssd1 vccd1 vccd1 _8325_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5537_ _8256_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7726_/D sky130_fd_sc_hd__and3_1
XFILLER_0_131_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5106__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6303__A1 _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8256_ _8256_/CLK _8256_/D vssd1 vssd1 vccd1 vccd1 _8256_/Q sky130_fd_sc_hd__dfxtp_1
X_5468_ _5468_/A _5470_/B _5468_/C vssd1 vssd1 vccd1 vccd1 _5468_/X sky130_fd_sc_hd__and3_1
X_4419_ _4419_/A _4425_/B vssd1 vssd1 vccd1 vccd1 _4419_/Y sky130_fd_sc_hd__nor2_1
X_5399_ _5399_/A vssd1 vssd1 vccd1 vccd1 _5399_/Y sky130_fd_sc_hd__inv_2
X_8187_ _8283_/CLK _8187_/D vssd1 vssd1 vccd1 vccd1 _8187_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout300 _5731_/Y vssd1 vssd1 vccd1 vccd1 _6398_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout322 _4024_/X vssd1 vssd1 vccd1 vccd1 _6931_/A sky130_fd_sc_hd__buf_4
Xfanout311 _5260_/Y vssd1 vssd1 vccd1 vccd1 _5294_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout366 hold1725/X vssd1 vssd1 vccd1 vccd1 _3968_/A sky130_fd_sc_hd__buf_8
Xfanout344 _3717_/X vssd1 vssd1 vccd1 vccd1 _6961_/A sky130_fd_sc_hd__buf_4
Xfanout333 _3862_/X vssd1 vssd1 vccd1 vccd1 _6949_/A sky130_fd_sc_hd__buf_4
X_7069_ _7069_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7069_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout388 _4720_/S0 vssd1 vssd1 vccd1 vccd1 _4734_/S0 sky130_fd_sc_hd__buf_4
Xfanout399 hold1659/X vssd1 vssd1 vccd1 vccd1 _7057_/A sky130_fd_sc_hd__clkbuf_8
Xfanout377 _4741_/S1 vssd1 vssd1 vccd1 vccd1 _4734_/S1 sky130_fd_sc_hd__clkbuf_4
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4712__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5290__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6425__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4644__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3768__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6790__A1 _7008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5593__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7256__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput19 i_instr_ID[28] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_1
XFILLER_0_18_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4779__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5345__A2 _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4951__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5281__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4084__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4703__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4554__S _7365_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3678__B _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6230__B1 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _6524_/A _4770_/B vssd1 vssd1 vccd1 vccd1 _8127_/D sky130_fd_sc_hd__and2_1
XFILLER_0_7_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3721_ _3721_/A1 _4073_/A2 _6961_/A _4073_/B2 _3720_/X vssd1 vssd1 vccd1 vccd1 _6447_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_130_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3652_ _7660_/Q vssd1 vssd1 vccd1 vccd1 _3652_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_113_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6440_ _7017_/A _6440_/B vssd1 vssd1 vccd1 vccd1 _7922_/D sky130_fd_sc_hd__and2_1
XFILLER_0_3_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6371_ _6371_/A _6371_/B vssd1 vssd1 vccd1 vccd1 _6380_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8110_ _8110_/CLK _8110_/D vssd1 vssd1 vccd1 vccd1 _8110_/Q sky130_fd_sc_hd__dfxtp_1
X_5322_ _6951_/A _5332_/A2 _5332_/B1 hold471/X vssd1 vssd1 vccd1 vccd1 _5322_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_121_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8041_ _8041_/CLK _8041_/D vssd1 vssd1 vccd1 vccd1 _8041_/Q sky130_fd_sc_hd__dfxtp_1
X_5253_ _6959_/A _5226_/B _5259_/B1 hold376/X vssd1 vssd1 vccd1 vccd1 _5253_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6392__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4729__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5184_ _7937_/Q _5222_/B _5183_/X vssd1 vssd1 vccd1 vccd1 _6908_/C sky130_fd_sc_hd__or3b_4
X_4204_ _4194_/Y _4198_/B _4196_/B vssd1 vssd1 vccd1 vccd1 _4205_/B sky130_fd_sc_hd__o21a_1
XANTENNA__6049__B1 _6048_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4135_ _6318_/A _6315_/A vssd1 vssd1 vccd1 vccd1 _4135_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5272__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4066_ _4066_/A _4066_/B vssd1 vssd1 vccd1 vccd1 _4090_/B sky130_fd_sc_hd__and2_1
XANTENNA__6064__A3 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A _5299_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7825_ _8486_/CLK _7825_/D vssd1 vssd1 vccd1 vccd1 _7825_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6221__B1 _6347_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6899__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7756_ _8071_/CLK _7756_/D vssd1 vssd1 vccd1 vccd1 _7756_/Q sky130_fd_sc_hd__dfxtp_1
X_4968_ _8193_/Q _8225_/Q _8289_/Q _7797_/Q _4983_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4968_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6772__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6707_ _6777_/A _6705_/B _6738_/B1 hold767/X vssd1 vssd1 vccd1 vccd1 _6707_/X sky130_fd_sc_hd__a22o_1
X_4899_ _8473_/Q _8405_/Q _8437_/Q _8311_/Q _4997_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4899_/X sky130_fd_sc_hd__mux4_1
X_3919_ _4014_/A _3917_/Y _3918_/Y vssd1 vssd1 vccd1 vccd1 _3919_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_74_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7687_ _8319_/CLK _7687_/D vssd1 vssd1 vccd1 vccd1 _7687_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3808__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__7076__A _7076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6638_ _7015_/A _6638_/A2 _6605_/B _6637_/X vssd1 vssd1 vccd1 vccd1 _6638_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5327__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_7191__69 _8328_/CLK vssd1 vssd1 vccd1 vccd1 _8104_/CLK sky130_fd_sc_hd__inv_2
X_6569_ _6925_/A _6592_/A2 _6592_/B1 hold404/X vssd1 vssd1 vccd1 vccd1 _6569_/X sky130_fd_sc_hd__a22o_1
X_8308_ _8477_/CLK _8308_/D vssd1 vssd1 vccd1 vccd1 _8308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_131_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6288__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8239_ _8239_/CLK _8239_/D vssd1 vssd1 vccd1 vccd1 _8239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout174 hold1510/X vssd1 vssd1 vccd1 vccd1 _5542_/B sky130_fd_sc_hd__buf_4
Xfanout163 _5002_/X vssd1 vssd1 vccd1 vccd1 _5182_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__4933__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _5879_/S vssd1 vssd1 vccd1 vccd1 _5963_/S sky130_fd_sc_hd__buf_4
Xfanout185 _5797_/S vssd1 vssd1 vccd1 vccd1 _5859_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__6155__A _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6763__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5318__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4621__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6374__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4924__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5254__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5940_ _5694_/Y _5939_/X _5936_/Y _6083_/A vssd1 vssd1 vccd1 vccd1 _5940_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4688__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7610_ _8368_/CLK _7610_/D vssd1 vssd1 vccd1 vccd1 _7610_/Q sky130_fd_sc_hd__dfxtp_1
X_5871_ _5871_/A _5871_/B vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4822_ _8462_/Q _8394_/Q _8426_/Q _8300_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4822_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6754__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7541_ _8343_/CLK _7541_/D vssd1 vssd1 vccd1 vccd1 _7541_/Q sky130_fd_sc_hd__dfxtp_1
X_4753_ _7006_/A _4753_/B vssd1 vssd1 vccd1 vccd1 _8110_/D sky130_fd_sc_hd__and2_1
XFILLER_0_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4860__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3704_ _3705_/A _3705_/B _3705_/C _3705_/D vssd1 vssd1 vccd1 vccd1 _3939_/B sky130_fd_sc_hd__nor4_1
XANTENNA__5309__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7472_ _8350_/CLK _7472_/D vssd1 vssd1 vccd1 vccd1 _7472_/Q sky130_fd_sc_hd__dfxtp_1
X_4684_ _8189_/Q _8221_/Q _8285_/Q _7793_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4684_/X sky130_fd_sc_hd__mux4_1
X_6423_ _7267_/A _6423_/B vssd1 vssd1 vccd1 vccd1 _7905_/D sky130_fd_sc_hd__nor2_1
XANTENNA__4612__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5190__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6354_ _6355_/B _6355_/C _6355_/A vssd1 vssd1 vccd1 vccd1 _6354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6285_ _6215_/X _6284_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6285_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3871__B _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5305_ _6917_/A _5299_/B _5331_/B1 hold725/X vssd1 vssd1 vccd1 vccd1 _5305_/X sky130_fd_sc_hd__a22o_1
X_8024_ _8457_/CLK _8024_/D vssd1 vssd1 vccd1 vccd1 _8024_/Q sky130_fd_sc_hd__dfxtp_2
X_5236_ _6925_/A _5226_/B _5259_/B1 hold873/X vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6690__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1801 _7892_/Q vssd1 vssd1 vccd1 vccd1 hold1801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1812 _7897_/Q vssd1 vssd1 vccd1 vccd1 hold1812/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1823 _7872_/Q vssd1 vssd1 vccd1 vccd1 hold1823/X sky130_fd_sc_hd__dlygate4sd3_1
X_5167_ _5463_/A _5463_/C vssd1 vssd1 vccd1 vccd1 _5167_/X sky130_fd_sc_hd__or2_1
XANTENNA__5245__A1 _6877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5098_ input10/X _4448_/B _5140_/B1 _5097_/X vssd1 vssd1 vccd1 vccd1 _7361_/D sky130_fd_sc_hd__o211a_1
X_4118_ _4118_/A _5955_/A vssd1 vssd1 vccd1 vccd1 _4118_/Y sky130_fd_sc_hd__nand2_1
X_4049_ _4049_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _4049_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6993__A1 _7065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1492_A _7309_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6745__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7808_ _8426_/CLK _7808_/D vssd1 vssd1 vccd1 vccd1 _7808_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4922__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7739_ _8519_/CLK _7739_/D vssd1 vssd1 vccd1 vccd1 _7739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6681__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4906__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5236__A1 _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4039__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5501__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6613__A _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6736__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4842__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold408 _7315_/Q vssd1 vssd1 vccd1 vccd1 _5412_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3970__A1 _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold419 _7452_/Q vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5172__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3722__A1 _6447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ _5734_/A _6058_/Y _6069_/Y _6163_/A vssd1 vssd1 vccd1 vccd1 _6070_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5899__A _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6672__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5021_ _5420_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5021_/X sky130_fd_sc_hd__or2_1
Xhold1108 _5241_/X vssd1 vssd1 vccd1 vccd1 _7449_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1119 _8441_/Q vssd1 vssd1 vccd1 vccd1 _6952_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5411__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6972_ _7029_/A _6972_/A2 _6908_/X _6971_/X vssd1 vssd1 vccd1 vccd1 _6972_/X sky130_fd_sc_hd__a31o_1
X_5923_ _5923_/A _5923_/B vssd1 vssd1 vccd1 vccd1 _5923_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4027__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6523__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5854_ _3910_/B _6398_/A2 _6413_/B1 _6302_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _5854_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4742__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6727__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4805_ _8137_/Q _7536_/Q _7408_/Q _7568_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4805_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4833__S0 _7357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4043__A _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5785_ _5778_/X _5784_/X _6302_/A vssd1 vssd1 vccd1 vccd1 _5785_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6242__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7524_ _7524_/CLK _7524_/D vssd1 vssd1 vccd1 vccd1 _7524_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout223_A _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4736_ _4735_/X _4732_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7530_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4667_ _8347_/Q _7823_/Q _7489_/Q _7457_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4667_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7455_ _8445_/CLK _7455_/D vssd1 vssd1 vccd1 vccd1 _7455_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7161__39 _8466_/CLK vssd1 vssd1 vccd1 vccd1 _8041_/CLK sky130_fd_sc_hd__inv_2
X_7386_ _8368_/CLK _7386_/D vssd1 vssd1 vccd1 vccd1 _7386_/Q sky130_fd_sc_hd__dfxtp_1
Xhold931 _7417_/Q vssd1 vssd1 vccd1 vccd1 hold931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold920 _5342_/X vssd1 vssd1 vccd1 vccd1 _7569_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6406_ _6406_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6406_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold942 _6567_/X vssd1 vssd1 vccd1 vccd1 _8139_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 _7874_/Q vssd1 vssd1 vccd1 vccd1 _4750_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7073__B _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6337_ _6338_/A _6338_/B vssd1 vssd1 vccd1 vccd1 _6337_/Y sky130_fd_sc_hd__nand2_1
X_4598_ _8144_/Q _7543_/Q _7415_/Q _7575_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4598_/X sky130_fd_sc_hd__mux4_1
Xhold964 _6591_/X vssd1 vssd1 vccd1 vccd1 _8163_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 _5329_/X vssd1 vssd1 vccd1 vccd1 _7560_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 _7423_/Q vssd1 vssd1 vccd1 vccd1 hold997/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 _7455_/Q vssd1 vssd1 vccd1 vccd1 hold975/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6268_ _6244_/A _6209_/A _6262_/A _6226_/A _5859_/S _5782_/S vssd1 vssd1 vccd1 vccd1
+ _6268_/X sky130_fd_sc_hd__mux4_1
X_6199_ _3799_/A _6414_/B1 _6398_/B1 _6188_/A _6417_/A2 vssd1 vssd1 vccd1 vccd1 _6199_/X
+ sky130_fd_sc_hd__a221o_1
X_5219_ _6967_/A _5188_/B _5220_/B1 _5219_/B2 vssd1 vssd1 vccd1 vccd1 _5219_/X sky130_fd_sc_hd__a22o_1
X_8007_ _8032_/CLK _8007_/D vssd1 vssd1 vccd1 vccd1 _8007_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1631 _7677_/Q vssd1 vssd1 vccd1 vccd1 _4039_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1642 _8506_/Q vssd1 vssd1 vccd1 vccd1 _4085_/A0 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1653 _7346_/Q vssd1 vssd1 vccd1 vccd1 _5391_/A sky130_fd_sc_hd__clkbuf_4
Xhold1620 _4324_/X vssd1 vssd1 vccd1 vccd1 _4325_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_84_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1686 _7356_/Q vssd1 vssd1 vccd1 vccd1 _6986_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1664 _7699_/Q vssd1 vssd1 vccd1 vccd1 _3839_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5218__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1675 _7698_/Q vssd1 vssd1 vccd1 vccd1 _3807_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1697 _7683_/Q vssd1 vssd1 vccd1 vccd1 _4073_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6966__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6433__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_99_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4652__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6718__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7264__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_0_0_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5154__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4827__S _7059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5209__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6709__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4815__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5932__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ _7005_/A _5570_/B vssd1 vssd1 vccd1 vccd1 _7759_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4521_ _8133_/Q _7532_/Q _7404_/Q _7564_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4521_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_81_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4452_ _7935_/Q _7018_/A vssd1 vssd1 vccd1 vccd1 _8099_/D sky130_fd_sc_hd__and2_1
Xhold216 _7335_/Q vssd1 vssd1 vccd1 vccd1 _5432_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 _5429_/X vssd1 vssd1 vccd1 vccd1 _7618_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _6709_/X vssd1 vssd1 vccd1 vccd1 _8264_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _7534_/Q vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 _5447_/X vssd1 vssd1 vccd1 vccd1 _7636_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5696__A1 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4383_ _4383_/A _4383_/B vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__or2_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6122_ _6039_/X _6121_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6122_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ _6053_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6056_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__6518__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _7258_/A _5004_/B hold1512/X vssd1 vssd1 vccd1 vccd1 _7314_/D sky130_fd_sc_hd__or3b_1
XANTENNA__4120__B2 _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__B _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6660__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4038__A _4753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A hold1510/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6948__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__7070__B1 _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6955_ _6955_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6955_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout340_A _3767_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5906_ _6144_/S _5906_/B vssd1 vssd1 vccd1 vccd1 _5906_/Y sky130_fd_sc_hd__nand2_1
X_7206__84 _8463_/CLK vssd1 vssd1 vccd1 vccd1 _8119_/CLK sky130_fd_sc_hd__inv_2
X_6886_ _7019_/A _6886_/A2 _6845_/B _6885_/X vssd1 vssd1 vccd1 vccd1 _6886_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout438_A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5837_ _5832_/X _5836_/Y _6270_/A vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5768_ _3934_/B _5971_/B _5772_/S vssd1 vssd1 vccd1 vccd1 _5769_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_16_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8487_ _8487_/CLK _8487_/D vssd1 vssd1 vccd1 vccd1 _8487_/Q sky130_fd_sc_hd__dfxtp_1
X_4719_ _8194_/Q _8226_/Q _8290_/Q _7798_/Q _4720_/S0 _4741_/S1 vssd1 vssd1 vccd1
+ vccd1 _4719_/X sky130_fd_sc_hd__mux4_1
X_7507_ _7507_/CLK _7507_/D vssd1 vssd1 vccd1 vccd1 _7507_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7438_ _8339_/CLK _7438_/D vssd1 vssd1 vccd1 vccd1 _7438_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7084__A _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5136__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5699_ _6016_/A _5974_/A _6035_/A _5993_/A _5860_/S _5789_/S vssd1 vssd1 vccd1 vccd1
+ _5699_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_71_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7369_ _8028_/CLK _7369_/D vssd1 vssd1 vccd1 vccd1 _7369_/Q sky130_fd_sc_hd__dfxtp_1
Xhold772 _6735_/X vssd1 vssd1 vccd1 vccd1 _8290_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold761 _7797_/Q vssd1 vssd1 vccd1 vccd1 hold761/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold750 _5357_/X vssd1 vssd1 vccd1 vccd1 _7584_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 _7537_/Q vssd1 vssd1 vccd1 vccd1 hold783/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold794 _6729_/X vssd1 vssd1 vccd1 vccd1 _8284_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1450 _4219_/X vssd1 vssd1 vccd1 vccd1 _5560_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _7882_/Q vssd1 vssd1 vccd1 vccd1 _4758_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1483 _7296_/Q vssd1 vssd1 vccd1 vccd1 _5148_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1494 hold1816/X vssd1 vssd1 vccd1 vccd1 _4765_/B sky130_fd_sc_hd__buf_1
Xhold1472 hold1812/X vssd1 vssd1 vccd1 vccd1 _4773_/B sky130_fd_sc_hd__buf_2
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7259__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6163__A _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5611__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5226__B _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6890__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4557__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4102__A1 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6642__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3861__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6740_ _7939_/Q _7940_/Q _6740_/C vssd1 vssd1 vccd1 vccd1 _6742_/B sky130_fd_sc_hd__or3_1
XANTENNA__5602__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_109_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8483_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4405__A2 _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3952_ _3923_/B _7945_/Q vssd1 vssd1 vccd1 vccd1 _3952_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6671_ _6777_/A _6670_/B _6670_/Y hold274/X vssd1 vssd1 vccd1 vccd1 _6671_/X sky130_fd_sc_hd__o22a_1
X_3883_ _3883_/A _3883_/B vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__and2_1
X_5622_ _6777_/A _5621_/B _5621_/Y hold224/X vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5905__A2 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8410_ _8427_/CLK _8410_/D vssd1 vssd1 vccd1 vccd1 _8410_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5366__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5553_ _6520_/A _5553_/B vssd1 vssd1 vccd1 vccd1 _7742_/D sky130_fd_sc_hd__and2_1
XFILLER_0_54_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8341_ _8450_/CLK _8341_/D vssd1 vssd1 vccd1 vccd1 _8341_/Q sky130_fd_sc_hd__dfxtp_1
X_4504_ _5144_/A1 _4504_/A1 _5451_/C vssd1 vssd1 vccd1 vccd1 _7294_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5118__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8272_ _8462_/CLK _8272_/D vssd1 vssd1 vccd1 vccd1 _8272_/Q sky130_fd_sc_hd__dfxtp_1
X_5484_ _7505_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7673_/D sky130_fd_sc_hd__and3_1
XFILLER_0_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4435_ _4200_/B _4435_/B vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__nand2b_1
X_4366_ _5477_/A _7734_/Q vssd1 vssd1 vccd1 vccd1 _4367_/D sky130_fd_sc_hd__xor2_1
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6105_ _4090_/A _6105_/A2 _6103_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6105_/X sky130_fd_sc_hd__a22o_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout290_A _6703_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7085_ _5545_/A _6975_/C _7080_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _7086_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _4398_/A _4395_/B vssd1 vssd1 vccd1 vccd1 _4392_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout388_A _4720_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6036_ _6036_/A _6036_/B vssd1 vssd1 vccd1 vccd1 _6038_/A sky130_fd_sc_hd__nor2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7043__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7987_ _8019_/CLK hold58/X vssd1 vssd1 vccd1 vccd1 _7987_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6938_ _7019_/A _6938_/A2 _6943_/B _6937_/X vssd1 vssd1 vccd1 vccd1 _6938_/X sky130_fd_sc_hd__a31o_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6869_ _6935_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6869_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6149__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5357__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3907__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold580 _7000_/X vssd1 vssd1 vccd1 vccd1 _8458_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6872__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold591 _8269_/Q vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6624__A3 _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1280 _8178_/Q vssd1 vssd1 vccd1 vccd1 _6628_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1291 _6654_/X vssd1 vssd1 vccd1 vccd1 _8191_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6605__B _6605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output105_A _7300_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5596__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5060__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7197__75 _8519_/CLK vssd1 vssd1 vccd1 vccd1 _8110_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_95_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6621__A _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5348__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput107 _7302_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[20] sky130_fd_sc_hd__buf_12
Xoutput129 _8046_/Q vssd1 vssd1 vccd1 vccd1 o_write_data_M[11] sky130_fd_sc_hd__buf_12
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput118 _7312_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[30] sky130_fd_sc_hd__buf_12
XFILLER_0_121_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4220_ _4219_/X _5022_/A1 _5453_/B vssd1 vssd1 vccd1 vccd1 _4227_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3980__A _4751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4151_ _5690_/A _5727_/C _4149_/X vssd1 vssd1 vccd1 vccd1 _5733_/C sky130_fd_sc_hd__o21a_1
X_4082_ _4757_/B _3676_/A _4082_/B1 _6935_/A _4081_/X vssd1 vssd1 vccd1 vccd1 _6075_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7910_ _8090_/CLK _7910_/D vssd1 vssd1 vccd1 vccd1 _7910_/Q sky130_fd_sc_hd__dfxtp_1
X_7841_ _8360_/CLK _7841_/D vssd1 vssd1 vccd1 vccd1 _7841_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6379__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7772_ _8326_/CLK _7772_/D vssd1 vssd1 vccd1 vccd1 _7772_/Q sky130_fd_sc_hd__dfxtp_1
X_4984_ _4983_/X _4982_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4984_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3935_ _3935_/A _3935_/B vssd1 vssd1 vccd1 vccd1 _3935_/X sky130_fd_sc_hd__and2_1
X_6723_ _6941_/A _6705_/B _6738_/B1 hold583/X vssd1 vssd1 vccd1 vccd1 _6723_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6531__A _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6654_ _7017_/A _6654_/A2 _6666_/A3 _6653_/X vssd1 vssd1 vccd1 vccd1 _6654_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_6_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5605_ _6947_/A _5616_/A2 _5616_/B1 hold739/X vssd1 vssd1 vccd1 vccd1 _5605_/X sky130_fd_sc_hd__a22o_1
X_3866_ _3968_/A _6441_/B _3865_/Y vssd1 vssd1 vccd1 vccd1 _6206_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3797_ _6191_/A _6188_/A vssd1 vssd1 vccd1 vccd1 _3799_/A sky130_fd_sc_hd__or2_1
XFILLER_0_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6585_ _6891_/A _6559_/B _6591_/B1 hold991/X vssd1 vssd1 vccd1 vccd1 _6585_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_131_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5536_ _8255_/Q _5538_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7725_/D sky130_fd_sc_hd__and3_1
XANTENNA_fanout303_A _5618_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8324_ _8450_/CLK _8324_/D vssd1 vssd1 vccd1 vccd1 _8324_/Q sky130_fd_sc_hd__dfxtp_1
X_8255_ _8255_/CLK _8255_/D vssd1 vssd1 vccd1 vccd1 _8255_/Q sky130_fd_sc_hd__dfxtp_1
X_5467_ hold67/X _5470_/B _5468_/C vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__and3_1
XFILLER_0_41_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4418_ _4425_/A _4422_/B _4241_/C vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6303__A2 _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6854__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout312 _5260_/Y vssd1 vssd1 vccd1 vccd1 _5262_/B sky130_fd_sc_hd__buf_6
Xfanout323 _4011_/X vssd1 vssd1 vccd1 vccd1 _6925_/A sky130_fd_sc_hd__buf_4
X_5398_ _7065_/A _6977_/B _7071_/A vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__o21a_1
Xfanout301 _5734_/A vssd1 vssd1 vccd1 vccd1 _6391_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8186_ _8346_/CLK _8186_/D vssd1 vssd1 vccd1 vccd1 _8186_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout356 _6909_/A vssd1 vssd1 vccd1 vccd1 _6777_/A sky130_fd_sc_hd__clkbuf_8
Xfanout345 _3966_/B vssd1 vssd1 vccd1 vccd1 _4072_/B sky130_fd_sc_hd__buf_8
X_4349_ _8489_/Q _7658_/Q vssd1 vssd1 vccd1 vccd1 _4350_/B sky130_fd_sc_hd__nand2_1
Xfanout334 _3851_/X vssd1 vssd1 vccd1 vccd1 _6953_/A sky130_fd_sc_hd__buf_4
Xfanout367 hold1725/X vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__buf_4
X_7068_ _7071_/B _7068_/A2 _7090_/A vssd1 vssd1 vccd1 vccd1 _7068_/Y sky130_fd_sc_hd__a21oi_1
Xfanout378 _4741_/S1 vssd1 vssd1 vccd1 vccd1 _4731_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout389 _4720_/S0 vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__buf_8
XANTENNA__4925__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6019_ _6008_/A _5814_/B _5955_/Y vssd1 vssd1 vccd1 vccd1 _6019_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6706__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3825__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5290__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6425__B _6425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4101__A_N _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6441__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4002__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7272__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5504__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5281__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3816__B1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6230__A1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3720_ _4770_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3720_/X sky130_fd_sc_hd__and2_1
XFILLER_0_130_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _8428_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6351__A _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3651_ _3651_/A vssd1 vssd1 vccd1 vccd1 _5073_/A sky130_fd_sc_hd__inv_2
XFILLER_0_130_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6370_ _6370_/A _6370_/B vssd1 vssd1 vccd1 vccd1 _6371_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7089__A3 _7069_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5321_ _6949_/A _5299_/B _5331_/B1 _5321_/B2 vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__a22o_1
X_8040_ _8040_/CLK _8040_/D vssd1 vssd1 vccd1 vccd1 _8040_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6392__S1 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6836__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5252_ _6891_/A _5258_/A2 _5258_/B1 hold449/X vssd1 vssd1 vccd1 vccd1 _5252_/X sky130_fd_sc_hd__a22o_1
X_5183_ _7006_/A _7936_/Q vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__and2_1
X_4203_ _4201_/Y _4203_/B vssd1 vssd1 vccd1 vccd1 _4203_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__5414__B _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6049__A1 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6049__B2 _6198_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4134_ _4128_/X _4132_/X _4133_/Y _3897_/A vssd1 vssd1 vccd1 vccd1 _4134_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5272__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4065_ _6053_/A _4065_/B vssd1 vssd1 vccd1 vccd1 _4066_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6526__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4124__A_N _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7824_ _8478_/CLK _7824_/D vssd1 vssd1 vccd1 vccd1 _7824_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout253_A _5620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5024__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7755_ _8379_/CLK _7755_/D vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__6772__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4967_ _4965_/X _4966_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__mux2_1
X_6706_ _6706_/A _6706_/B vssd1 vssd1 vccd1 vccd1 _6706_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_31_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8462_/CLK sky130_fd_sc_hd__clkbuf_16
X_4898_ _8183_/Q _8215_/Q _8279_/Q _7787_/Q _4996_/S0 _4997_/S1 vssd1 vssd1 vccd1
+ vccd1 _4898_/X sky130_fd_sc_hd__mux4_1
X_3918_ _4014_/A _4161_/A vssd1 vssd1 vccd1 vccd1 _3918_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_fanout420_A _7357_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6261__A _6262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7686_ _8355_/CLK _7686_/D vssd1 vssd1 vccd1 vccd1 _7686_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6637_ _6877_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6637_/X sky130_fd_sc_hd__and2_1
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3849_ _4067_/A_N _7961_/Q vssd1 vssd1 vccd1 vccd1 _3849_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_34_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6568_ _6923_/A _6559_/B _6591_/B1 hold729/X vssd1 vssd1 vccd1 vccd1 _6568_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5519_ _8238_/Q _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7708_/D sky130_fd_sc_hd__and3_1
X_8307_ _8469_/CLK _8307_/D vssd1 vssd1 vccd1 vccd1 _8307_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6499_ _6534_/A _6499_/B vssd1 vssd1 vccd1 vccd1 _6499_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8238_ _8238_/CLK _8238_/D vssd1 vssd1 vccd1 vccd1 _8238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8169_ _8468_/CLK _8169_/D vssd1 vssd1 vccd1 vccd1 _8169_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_98_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _8504_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout164 _5148_/B1 vssd1 vssd1 vccd1 vccd1 _5146_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout175 hold1510/X vssd1 vssd1 vccd1 vccd1 _5528_/B sky130_fd_sc_hd__buf_2
Xfanout197 _3920_/Y vssd1 vssd1 vccd1 vccd1 _5879_/S sky130_fd_sc_hd__clkbuf_4
Xfanout186 _5797_/S vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__buf_4
XANTENNA__4655__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6436__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6994__A1_N _7074_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6763__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7267__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7167__45 _8465_/CLK vssd1 vssd1 vccd1 vccd1 _8047_/CLK sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_22_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8477_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4621__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6818__A3 _6838_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6374__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_89_clk clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 _8091_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5254__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4688__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5870_ _5870_/A _5870_/B vssd1 vssd1 vccd1 vccd1 _5871_/B sky130_fd_sc_hd__or2_1
X_4821_ _8172_/Q _8204_/Q _8268_/Q _7776_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4821_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5006__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6203__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6754__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4752_ _6498_/A _4752_/B vssd1 vssd1 vccd1 vccd1 _8109_/D sky130_fd_sc_hd__and2_1
X_7540_ _8270_/CLK _7540_/D vssd1 vssd1 vccd1 vccd1 _7540_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_13_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _8419_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4860__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7471_ _7805_/CLK _7471_/D vssd1 vssd1 vccd1 vccd1 _7471_/Q sky130_fd_sc_hd__dfxtp_1
X_3703_ _3652_/Y _7937_/Q _7936_/Q vssd1 vssd1 vccd1 vccd1 _3705_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4683_ _4681_/X _4682_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4683_/X sky130_fd_sc_hd__mux2_1
X_6422_ _3939_/X _3940_/X _6422_/A3 _5667_/A vssd1 vssd1 vccd1 vccd1 _6422_/X sky130_fd_sc_hd__o31a_2
XANTENNA__4612__S1 _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5190__A1 _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6353_ _6353_/A vssd1 vssd1 vccd1 vccd1 _6355_/C sky130_fd_sc_hd__inv_2
XFILLER_0_12_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5304_ _6849_/A _5300_/B _5300_/Y hold360/X vssd1 vssd1 vccd1 vccd1 _5304_/X sky130_fd_sc_hd__o22a_1
X_6284_ _6281_/A _6244_/A _6262_/A _6226_/A _5859_/S _5744_/S vssd1 vssd1 vccd1 vccd1
+ _6284_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_11_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5235_ _6923_/A _5258_/A2 _5258_/B1 hold989/X vssd1 vssd1 vccd1 vccd1 _5235_/X sky130_fd_sc_hd__a22o_1
X_8023_ _8032_/CLK _8023_/D vssd1 vssd1 vccd1 vccd1 _8023_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1802 _7890_/Q vssd1 vssd1 vccd1 vccd1 hold1802/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6690__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1824 _7361_/Q vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1813 _7884_/Q vssd1 vssd1 vccd1 vccd1 hold1813/X sky130_fd_sc_hd__dlygate4sd3_1
X_5166_ _5166_/A1 _4416_/B _5166_/B1 _5165_/X vssd1 vssd1 vccd1 vccd1 _7395_/D sky130_fd_sc_hd__o211a_1
X_4117_ _4111_/X _4115_/X _4116_/Y _4092_/A vssd1 vssd1 vccd1 vccd1 _4117_/Y sky130_fd_sc_hd__a31oi_2
XFILLER_0_79_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout468_A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5097_ hold89/X _7030_/C vssd1 vssd1 vccd1 vccd1 _5097_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout370_A _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5245__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4048_ _8081_/Q _4047_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4048_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6745__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7807_ _8461_/CLK _7807_/D vssd1 vssd1 vccd1 vccd1 _7807_/Q sky130_fd_sc_hd__dfxtp_1
X_5999_ _6302_/A _5999_/B vssd1 vssd1 vccd1 vccd1 _5999_/Y sky130_fd_sc_hd__nor2_1
X_7738_ _8519_/CLK _7738_/D vssd1 vssd1 vccd1 vccd1 _7738_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1652_A _4004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7669_ _8080_/CLK _7669_/D vssd1 vssd1 vccd1 vccd1 _7669_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5705__A0 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5335__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6681__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5070__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5236__A2 _5226_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5501__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6613__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6736__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4842__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7225__103 _8461_/CLK vssd1 vssd1 vccd1 vccd1 _8235_/CLK sky130_fd_sc_hd__inv_2
Xhold409 _5412_/X vssd1 vssd1 vccd1 vccd1 _7601_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3970__A2 _3967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_output97_A _7292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6672__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5020_ _5020_/A1 _4425_/B _5146_/B1 _5019_/X vssd1 vssd1 vccd1 vccd1 _7322_/D sky130_fd_sc_hd__o211a_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clkbuf_4_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _8450_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold1109 _8417_/Q vssd1 vssd1 vccd1 vccd1 _6902_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5411__C _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6971_ _6971_/A _6971_/B vssd1 vssd1 vccd1 vccd1 _6971_/X sky130_fd_sc_hd__and2_1
XANTENNA__4530__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5922_ _5922_/A _5922_/B vssd1 vssd1 vccd1 vccd1 _5923_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5853_ _6342_/S _6144_/S _5853_/C vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__and3_1
XFILLER_0_61_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6727__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5784_ _5780_/X _5783_/X _5963_/S vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4804_ _8330_/Q _7806_/Q _7472_/Q _7440_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4804_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4833__S1 _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5139__B _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4735_ _4734_/X _4733_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4735_/X sky130_fd_sc_hd__mux2_1
X_7523_ _7523_/CLK _7523_/D vssd1 vssd1 vccd1 vccd1 _7523_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout216_A _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7454_ _8218_/CLK _7454_/D vssd1 vssd1 vccd1 vccd1 _7454_/Q sky130_fd_sc_hd__dfxtp_1
X_4666_ _4665_/X _4662_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7520_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_114_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7385_ _8370_/CLK _7385_/D vssd1 vssd1 vccd1 vccd1 _7385_/Q sky130_fd_sc_hd__dfxtp_1
X_6405_ _6405_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6405_/Y sky130_fd_sc_hd__nor2_1
X_4597_ _8337_/Q _7813_/Q _7479_/Q _7447_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4597_/X sky130_fd_sc_hd__mux4_1
Xhold910 _7020_/X vssd1 vssd1 vccd1 vccd1 _8478_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4597__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold921 _8159_/Q vssd1 vssd1 vccd1 vccd1 hold921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 _8107_/D vssd1 vssd1 vccd1 vccd1 _8073_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold932 _5203_/X vssd1 vssd1 vccd1 vccd1 _7417_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _8154_/Q vssd1 vssd1 vccd1 vccd1 hold943/X sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ _6320_/A _6319_/A _6317_/Y vssd1 vssd1 vccd1 vccd1 _6338_/B sky130_fd_sc_hd__a21o_1
Xhold965 _7477_/Q vssd1 vssd1 vccd1 vccd1 hold965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _5209_/X vssd1 vssd1 vccd1 vccd1 _7423_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 _5247_/X vssd1 vssd1 vccd1 vccd1 _7455_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 _8151_/Q vssd1 vssd1 vccd1 vccd1 hold987/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_782 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6267_ _6265_/Y _6266_/X _6391_/A vssd1 vssd1 vccd1 vccd1 _6267_/Y sky130_fd_sc_hd__a21oi_1
X_6198_ _5853_/X _6197_/X _6198_/S vssd1 vssd1 vccd1 vccd1 _6198_/X sky130_fd_sc_hd__mux2_1
X_5218_ _6965_/A _5188_/B _5220_/B1 hold955/X vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__a22o_1
X_8006_ _8096_/CLK _8006_/D vssd1 vssd1 vccd1 vccd1 _8006_/Q sky130_fd_sc_hd__dfxtp_1
Xhold1610 _4253_/X vssd1 vssd1 vccd1 vccd1 _5565_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1632 _4039_/X vssd1 vssd1 vccd1 vccd1 _6430_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1643 _7736_/Q vssd1 vssd1 vccd1 vccd1 _4155_/A1 sky130_fd_sc_hd__dlygate4sd3_1
X_5149_ _5454_/A _5454_/C vssd1 vssd1 vccd1 vccd1 _5149_/X sky130_fd_sc_hd__or2_1
Xhold1621 _4325_/Y vssd1 vssd1 vccd1 vccd1 _5575_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1687 _7693_/Q vssd1 vssd1 vccd1 vccd1 _3709_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6415__B2 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1676 _3807_/X vssd1 vssd1 vccd1 vccd1 _6451_/B sky130_fd_sc_hd__buf_1
XANTENNA__5218__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1654 _8492_/Q vssd1 vssd1 vccd1 vccd1 _3745_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1665 _7651_/Q vssd1 vssd1 vccd1 vccd1 _4299_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1698 _4073_/X vssd1 vssd1 vccd1 vccd1 _6436_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4521__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6718__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7137__15 _8154_/CLK vssd1 vssd1 vccd1 vccd1 _7514_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_62_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3792__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5065__A _5404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7280__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6654__A1 _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5512__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5209__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5090__B1 _5002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4815__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3983__A _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6590__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4520_ _8326_/Q _7802_/Q _7468_/Q _7436_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4520_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4579__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4451_ _5003_/A0 _4163_/Y _5442_/C vssd1 vssd1 vccd1 vccd1 _8358_/D sky130_fd_sc_hd__mux2_1
Xhold217 _5432_/X vssd1 vssd1 vccd1 vccd1 _7621_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold206 _7617_/Q vssd1 vssd1 vccd1 vccd1 _5675_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _7564_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _5303_/X vssd1 vssd1 vccd1 vccd1 _7534_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5696__A2 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6121_ _6096_/A _6056_/A _6115_/A _6075_/A _5859_/S _5782_/S vssd1 vssd1 vccd1 vccd1
+ _6121_/X sky130_fd_sc_hd__mux4_1
X_4382_ _4382_/A _5069_/S vssd1 vssd1 vccd1 vccd1 _4382_/X sky130_fd_sc_hd__and2_1
XFILLER_0_0_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6034_/Y _6038_/B _6036_/B vssd1 vssd1 vccd1 vccd1 _6058_/A sky130_fd_sc_hd__a21o_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5422__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5003_ _5003_/A0 _5411_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5004_/B sky130_fd_sc_hd__mux2_1
XANTENNA__4120__A2 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4038__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7070__A1 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6534__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout166_A _5002_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6954_ _7026_/A _6954_/A2 _6970_/A3 _6953_/X vssd1 vssd1 vccd1 vccd1 _6954_/X sky130_fd_sc_hd__a31o_1
X_5905_ _5846_/A _5820_/A _5892_/A _5870_/A _5744_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _5906_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6885_ _6951_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6885_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7221__99 _8388_/CLK vssd1 vssd1 vccd1 vccd1 _8231_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_91_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5836_ _5836_/A _5836_/B vssd1 vssd1 vccd1 vccd1 _5836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5767_ _5765_/X _5767_/B vssd1 vssd1 vccd1 vccd1 _5769_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_72_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3893__A _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6581__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7506_ _7506_/CLK _7506_/D vssd1 vssd1 vccd1 vccd1 _7506_/Q sky130_fd_sc_hd__dfxtp_1
X_5698_ _6016_/A _6035_/A _5789_/S vssd1 vssd1 vccd1 vccd1 _5698_/X sky130_fd_sc_hd__mux2_1
X_4718_ _4716_/X _4717_/X _4735_/S vssd1 vssd1 vccd1 vccd1 _4718_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8486_ _8486_/CLK _8486_/D vssd1 vssd1 vccd1 vccd1 _8486_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7437_ _8458_/CLK _7437_/D vssd1 vssd1 vccd1 vccd1 _7437_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7084__B _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4649_ _8184_/Q _8216_/Q _8280_/Q _7788_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4649_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6884__A1 _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7368_ _8462_/CLK _7368_/D vssd1 vssd1 vccd1 vccd1 _7368_/Q sky130_fd_sc_hd__dfxtp_1
Xhold773 _8268_/Q vssd1 vssd1 vccd1 vccd1 hold773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 _7418_/Q vssd1 vssd1 vccd1 vccd1 hold751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 _5605_/X vssd1 vssd1 vccd1 vccd1 _7789_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _5613_/X vssd1 vssd1 vccd1 vccd1 _7797_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4928__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold784 _5306_/X vssd1 vssd1 vccd1 vccd1 _7537_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ _6319_/A _6319_/B vssd1 vssd1 vccd1 vccd1 _6320_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4990__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold795 _8321_/Q vssd1 vssd1 vccd1 vccd1 hold795/X sky130_fd_sc_hd__dlygate4sd3_1
X_7299_ _8373_/CLK _7299_/D _7109_/Y vssd1 vssd1 vccd1 vccd1 _7299_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__6636__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1451 _4227_/B vssd1 vssd1 vccd1 vccd1 _4427_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1440 hold1817/X vssd1 vssd1 vccd1 vccd1 _4764_/B sky130_fd_sc_hd__buf_2
Xhold1495 _8168_/Q vssd1 vssd1 vccd1 vccd1 _6607_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1473 _7301_/Q vssd1 vssd1 vccd1 vccd1 _5158_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 _7298_/Q vssd1 vssd1 vccd1 vccd1 _5152_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1462 _7306_/Q vssd1 vssd1 vccd1 vccd1 _5168_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5072__B1 _5140_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5611__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6572__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7275__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5507__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4838__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6619__A _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4102__A2 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4733__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3951_ _5838_/A _5765_/A vssd1 vssd1 vccd1 vccd1 _3951_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5602__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6670_ _6706_/A _6670_/B vssd1 vssd1 vccd1 vccd1 _6670_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3882_ _3882_/A _6259_/A vssd1 vssd1 vccd1 vccd1 _3883_/B sky130_fd_sc_hd__nand2_1
XANTENNA__6801__B _6839_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5621_ _6706_/A _5621_/B vssd1 vssd1 vccd1 vccd1 _5621_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5366__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5905__A3 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5552_ _6494_/A _5552_/B vssd1 vssd1 vccd1 vccd1 _7741_/D sky130_fd_sc_hd__and2_1
X_8340_ _8481_/CLK _8340_/D vssd1 vssd1 vccd1 vccd1 _8340_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4503_ _5146_/A1 _4422_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _7295_/D sky130_fd_sc_hd__mux2_1
X_8271_ _8425_/CLK _8271_/D vssd1 vssd1 vccd1 vccd1 _8271_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5417__B _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_83_clk_A clkbuf_4_5_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6866__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5483_ _7504_/Q _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _7672_/D sky130_fd_sc_hd__and3_1
X_4434_ _4434_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4434_/X sky130_fd_sc_hd__and2_1
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6529__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4365_ _5476_/A _7733_/Q vssd1 vssd1 vccd1 vccd1 _4367_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_111_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4972__S0 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7084_ _7088_/A _7088_/B _7084_/C vssd1 vssd1 vccd1 vccd1 _7084_/X sky130_fd_sc_hd__and3_1
X_6104_ _6096_/A _6094_/A _6398_/A2 vssd1 vssd1 vccd1 vccd1 _6104_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6618__A1 _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6035_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _6036_/B sky130_fd_sc_hd__nor2_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _5571_/B _4394_/A _5503_/B vssd1 vssd1 vccd1 vccd1 _4395_/B sky130_fd_sc_hd__mux2_1
XANTENNA_fanout283_A _6776_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4724__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout450_A _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5054__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7986_ _8090_/CLK hold38/X vssd1 vssd1 vccd1 vccd1 _7986_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6937_ _6937_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6937_/X sky130_fd_sc_hd__and2_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6868_ _7010_/A _6868_/A2 _6845_/B _6867_/X vssd1 vssd1 vccd1 vccd1 _6868_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_76_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5819_ _5963_/S _5971_/B vssd1 vssd1 vccd1 vccd1 _5820_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_91_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5357__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3907__A2 _3904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7095__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6799_ _6931_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6799_/X sky130_fd_sc_hd__and2_1
XFILLER_0_17_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8469_ _8469_/CLK _8469_/D vssd1 vssd1 vccd1 vccd1 _8469_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6439__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold581 _8270_/Q vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold570 _6699_/X vssd1 vssd1 vccd1 vccd1 _8226_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4658__S _5103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold592 _6714_/X vssd1 vssd1 vccd1 vccd1 _8269_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_109_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5293__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1270 _6818_/X vssd1 vssd1 vccd1 vccd1 _8346_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1281 _6628_/X vssd1 vssd1 vccd1 vccd1 _8178_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6174__A _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3798__A _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1292 _7886_/Q vssd1 vssd1 vccd1 vccd1 _4762_/B sky130_fd_sc_hd__buf_1
XANTENNA__5596__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6621__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5348__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3898__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6848__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput119 _7313_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[31] sky130_fd_sc_hd__buf_12
Xoutput108 _7303_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[21] sky130_fd_sc_hd__buf_12
XANTENNA__4568__S _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4954__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3980__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4150_ _8453_/Q _5732_/C _5688_/A vssd1 vssd1 vccd1 vccd1 _5727_/C sky130_fd_sc_hd__or3b_2
XFILLER_0_128_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput90 _8105_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[4] sky130_fd_sc_hd__buf_12
XFILLER_0_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4081_ _4081_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _4081_/X sky130_fd_sc_hd__or2_1
XANTENNA__5284__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4706__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7840_ _8030_/CLK hold36/X vssd1 vssd1 vccd1 vccd1 _7840_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5036__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5587__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7771_ _8326_/CLK _7771_/D vssd1 vssd1 vccd1 vccd1 _7771_/Q sky130_fd_sc_hd__dfxtp_1
X_4983_ _8485_/Q _8417_/Q _8449_/Q _8323_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4983_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_129_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3934_ _5789_/S _3934_/B vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__or2_1
X_6722_ _6939_/A _6737_/A2 _6737_/B1 hold703/X vssd1 vssd1 vccd1 vccd1 _6722_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5339__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6653_ _6959_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6653_/X sky130_fd_sc_hd__and2_1
XFILLER_0_46_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3865_ _3968_/A _4277_/A vssd1 vssd1 vccd1 vccd1 _3865_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5604_ _6945_/A _5616_/A2 _5616_/B1 hold495/X vssd1 vssd1 vccd1 vccd1 _5604_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_27_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3796_ _3796_/A0 _3795_/X _4074_/S vssd1 vssd1 vccd1 vccd1 _6188_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_42_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6584_ _6955_/A _6559_/B _6591_/B1 hold869/X vssd1 vssd1 vccd1 vccd1 _6584_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5147__B _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4051__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8323_ _8350_/CLK _8323_/D vssd1 vssd1 vccd1 vccd1 _8323_/Q sky130_fd_sc_hd__dfxtp_1
X_5535_ _8254_/Q _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _7724_/D sky130_fd_sc_hd__and3_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5466_ hold63/X _5470_/B _5468_/C vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__and3_1
XFILLER_0_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8254_ _8254_/CLK _8254_/D vssd1 vssd1 vccd1 vccd1 _8254_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6303__A3 _6244_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4417_ _5030_/A1 _4416_/B _4415_/X _4416_/Y vssd1 vssd1 vccd1 vccd1 _8371_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5397_ _7067_/A _7069_/A _6597_/B vssd1 vssd1 vccd1 vccd1 _5397_/Y sky130_fd_sc_hd__o21bai_1
Xfanout302 _6030_/A1 vssd1 vssd1 vccd1 vccd1 _5734_/A sky130_fd_sc_hd__clkbuf_8
X_8185_ _8445_/CLK _8185_/D vssd1 vssd1 vccd1 vccd1 _8185_/Q sky130_fd_sc_hd__dfxtp_1
Xfanout313 _5226_/B vssd1 vssd1 vccd1 vccd1 _5258_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4945__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout324 _4000_/X vssd1 vssd1 vccd1 vccd1 _6929_/A sky130_fd_sc_hd__buf_4
Xfanout346 _3966_/B vssd1 vssd1 vccd1 vccd1 _4083_/B sky130_fd_sc_hd__buf_4
Xfanout357 _3837_/X vssd1 vssd1 vccd1 vccd1 _6971_/A sky130_fd_sc_hd__buf_4
X_4348_ _8489_/Q _7658_/Q vssd1 vssd1 vccd1 vccd1 _4350_/A sky130_fd_sc_hd__or2_1
Xfanout335 _3826_/X vssd1 vssd1 vccd1 vccd1 _6967_/A sky130_fd_sc_hd__buf_4
X_7067_ _7067_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7067_/Y sky130_fd_sc_hd__nand2_1
Xfanout379 _7050_/A vssd1 vssd1 vccd1 vccd1 _4741_/S1 sky130_fd_sc_hd__clkbuf_4
Xfanout368 _7083_/B2 vssd1 vssd1 vccd1 vccd1 _7046_/A sky130_fd_sc_hd__buf_8
X_4279_ _4277_/Y _4279_/B vssd1 vssd1 vccd1 vccd1 _4281_/A sky130_fd_sc_hd__nand2b_1
X_6018_ _6018_/A _6018_/B vssd1 vssd1 vccd1 vccd1 _6018_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5275__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3825__B2 _8032_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7969_ _8030_/CLK _7969_/D vssd1 vssd1 vccd1 vccd1 _7969_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6790__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6441__B _6441_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4002__B2 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5772__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5057__B _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3761__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4388__S _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5504__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4069__A1 _4068_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5266__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3816__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5018__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6766__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4851__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3650_ _7067_/A vssd1 vssd1 vccd1 vccd1 _6977_/B sky130_fd_sc_hd__inv_2
XFILLER_0_130_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5320_ _6947_/A _5299_/B _5331_/B1 hold957/X vssd1 vssd1 vccd1 vccd1 _5320_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5251_ _6955_/A _5258_/A2 _5258_/B1 hold535/X vssd1 vssd1 vccd1 vccd1 _5251_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4927__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4202_ _8510_/Q _4202_/B vssd1 vssd1 vccd1 vccd1 _4202_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5414__C _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5182_ _5182_/A1 _5182_/A2 _5182_/B1 _5181_/X vssd1 vssd1 vccd1 vccd1 _7403_/D sky130_fd_sc_hd__o211a_1
X_4133_ _6262_/A _6259_/A vssd1 vssd1 vccd1 vccd1 _4133_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__6807__A _6939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4064_ _6053_/A _6056_/A vssd1 vssd1 vccd1 vccd1 _4066_/A sky130_fd_sc_hd__or2_1
XANTENNA__5257__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3807__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6757__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7823_ _8413_/CLK _7823_/D vssd1 vssd1 vccd1 vccd1 _7823_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6542__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6221__A2 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7754_ _8485_/CLK _7754_/D vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
X_6705_ _6741_/A _6705_/B vssd1 vssd1 vccd1 vccd1 _6705_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4966_ _8160_/Q _7559_/Q _7431_/Q _7591_/Q _4990_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4966_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7685_ _8464_/CLK _7685_/D vssd1 vssd1 vccd1 vccd1 _7685_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4897_ _4895_/X _4896_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4897_/X sky130_fd_sc_hd__mux2_1
X_3917_ _3917_/A1 _4084_/A2 _6847_/A _4084_/B2 _3916_/X vssd1 vssd1 vccd1 vccd1 _3917_/Y
+ sky130_fd_sc_hd__a221oi_4
XANTENNA__5980__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout413_A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7076__C _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6636_ _7019_/A _6636_/A2 _6666_/A3 _6635_/X vssd1 vssd1 vccd1 vccd1 _6636_/X sky130_fd_sc_hd__a31o_1
X_3848_ _3848_/A _3848_/B _3848_/C _6405_/A vssd1 vssd1 vccd1 vccd1 _3897_/C sky130_fd_sc_hd__or4_1
XFILLER_0_6_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6567_ _6921_/A _6592_/A2 _6592_/B1 hold941/X vssd1 vssd1 vccd1 vccd1 _6567_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3779_ _8085_/Q _3778_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8306_ _8466_/CLK _8306_/D vssd1 vssd1 vccd1 vccd1 _8306_/Q sky130_fd_sc_hd__dfxtp_1
X_5518_ _8237_/Q _5541_/B _7073_/B vssd1 vssd1 vccd1 vccd1 _7707_/D sky130_fd_sc_hd__and3_1
XFILLER_0_42_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3743__B1 _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6498_ _6498_/A hold94/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__and2_1
XANTENNA__6288__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5449_ _5449_/A _5453_/B _5449_/C vssd1 vssd1 vccd1 vccd1 _5449_/X sky130_fd_sc_hd__and3_1
X_8237_ _8237_/CLK _8237_/D vssd1 vssd1 vccd1 vccd1 _8237_/Q sky130_fd_sc_hd__dfxtp_1
X_8168_ _8458_/CLK _8168_/D vssd1 vssd1 vccd1 vccd1 _8168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout165 _5148_/B1 vssd1 vssd1 vccd1 vccd1 _5140_/B1 sky130_fd_sc_hd__clkbuf_8
X_7119_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7119_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4936__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5621__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 _3946_/X vssd1 vssd1 vccd1 vccd1 _5797_/S sky130_fd_sc_hd__buf_4
Xfanout176 _7073_/A vssd1 vssd1 vccd1 vccd1 _7082_/A sky130_fd_sc_hd__buf_4
Xfanout198 _6393_/A vssd1 vssd1 vccd1 vccd1 _6410_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__3840__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8099_ _8099_/CLK _8099_/D vssd1 vssd1 vccd1 vccd1 _8099_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5248__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6748__B1 _6774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4099__A_N _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5068__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4909__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5515__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5239__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820_ _4818_/X _4819_/X _5477_/A vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4581__S _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6362__A _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _6494_/A _4751_/B vssd1 vssd1 vccd1 vccd1 _8108_/D sky130_fd_sc_hd__and2_1
XFILLER_0_56_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3702_ _3700_/Y _3701_/X _3690_/Y vssd1 vssd1 vccd1 vccd1 _3705_/C sky130_fd_sc_hd__a21o_1
X_7470_ _8339_/CLK _7470_/D vssd1 vssd1 vccd1 vccd1 _7470_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4682_ _8156_/Q _7555_/Q _7427_/Q _7587_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4682_/X sky130_fd_sc_hd__mux4_1
X_6421_ _7258_/A _6421_/B vssd1 vssd1 vccd1 vccd1 _7903_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_71_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5190__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6352_ _6352_/A _6352_/B vssd1 vssd1 vccd1 vccd1 _6353_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_3_466 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5303_ _6847_/A _5300_/B _5300_/Y hold238/X vssd1 vssd1 vccd1 vccd1 _5303_/X sky130_fd_sc_hd__o22a_1
X_6283_ _6283_/A _6283_/B vssd1 vssd1 vccd1 vccd1 _6283_/X sky130_fd_sc_hd__xor2_1
XANTENNA__5425__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5234_ _6921_/A _5226_/B _5259_/B1 hold801/X vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__a22o_1
X_8022_ _8440_/CLK _8022_/D vssd1 vssd1 vccd1 vccd1 _8022_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__6690__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5165_ _5462_/A _5454_/C vssd1 vssd1 vccd1 vccd1 _5165_/X sky130_fd_sc_hd__or2_1
Xhold1814 _7369_/Q vssd1 vssd1 vccd1 vccd1 hold1814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1825 _7373_/Q vssd1 vssd1 vccd1 vccd1 hold1825/X sky130_fd_sc_hd__dlygate4sd3_1
X_4116_ _6115_/A _6112_/A vssd1 vssd1 vccd1 vccd1 _4116_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1803 _8376_/Q vssd1 vssd1 vccd1 vccd1 hold1803/X sky130_fd_sc_hd__dlygate4sd3_1
X_5096_ input9/X _5067_/S _5172_/B1 _5095_/X vssd1 vssd1 vccd1 vccd1 _7360_/D sky130_fd_sc_hd__o211a_1
X_4047_ _7985_/Q _4079_/A2 _4079_/B1 _8017_/Q _4046_/X vssd1 vssd1 vccd1 vccd1 _4047_/X
+ sky130_fd_sc_hd__a221o_4
XANTENNA__5650__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7806_ _8350_/CLK _7806_/D vssd1 vssd1 vccd1 vccd1 _7806_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4491__S _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5998_ _5906_/B _6080_/B _6144_/S vssd1 vssd1 vccd1 vccd1 _5999_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_59_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7737_ _8454_/CLK _7737_/D vssd1 vssd1 vccd1 vccd1 _7737_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4949_ _4948_/X _4947_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_129_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7668_ _8080_/CLK _7668_/D vssd1 vssd1 vccd1 vccd1 _7668_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3964__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6619_ _6925_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6619_/X sky130_fd_sc_hd__and2_1
XANTENNA__5705__A1 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7599_ _8507_/CLK _7599_/D vssd1 vssd1 vccd1 vccd1 _7599_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3716__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5335__B _5335_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6681__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4666__S _7046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5641__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7278__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5172__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6121__A1 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6672__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6970_ _6434_/A _6970_/A2 _6970_/A3 _6969_/X vssd1 vssd1 vccd1 vccd1 _6970_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5632__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5921_ _5921_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5922_/B sky130_fd_sc_hd__or2_1
XFILLER_0_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4530__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5852_ _5846_/A _5820_/A _5765_/A _3934_/B _5789_/S _5838_/A vssd1 vssd1 vccd1 vccd1
+ _5853_/C sky130_fd_sc_hd__mux4_2
XFILLER_0_76_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4803_ _4802_/X _4799_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8233_/D sky130_fd_sc_hd__mux2_1
X_5783_ _5781_/X _5782_/X _5860_/S vssd1 vssd1 vccd1 vccd1 _5783_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7522_ _7522_/CLK _7522_/D vssd1 vssd1 vccd1 vccd1 _7522_/Q sky130_fd_sc_hd__dfxtp_1
X_4734_ _8486_/Q _8418_/Q _8450_/Q _8324_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4734_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7453_ _8343_/CLK _7453_/D vssd1 vssd1 vccd1 vccd1 _7453_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5699__A0 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4665_ _4664_/X _4663_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4665_/X sky130_fd_sc_hd__mux2_1
X_7384_ _8368_/CLK _7384_/D vssd1 vssd1 vccd1 vccd1 _7384_/Q sky130_fd_sc_hd__dfxtp_1
X_4596_ _4595_/X _4592_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7510_/D sky130_fd_sc_hd__mux2_1
Xhold900 _5347_/X vssd1 vssd1 vccd1 vccd1 _7574_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5794__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6360__B2 _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6360__A1 _5739_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6404_ _6406_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6404_/X sky130_fd_sc_hd__or2_1
Xhold911 _7813_/Q vssd1 vssd1 vccd1 vccd1 hold911/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4597__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold922 _6587_/X vssd1 vssd1 vccd1 vccd1 _8159_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 _6582_/X vssd1 vssd1 vccd1 vccd1 _8154_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 _7432_/Q vssd1 vssd1 vccd1 vccd1 hold955/X sky130_fd_sc_hd__dlygate4sd3_1
X_6335_ _6335_/A _6335_/B vssd1 vssd1 vccd1 vccd1 _6338_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold933 _8320_/Q vssd1 vssd1 vccd1 vccd1 hold933/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold966 _5273_/X vssd1 vssd1 vccd1 vccd1 _7477_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 _7577_/Q vssd1 vssd1 vccd1 vccd1 hold977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 _6579_/X vssd1 vssd1 vccd1 vccd1 _8151_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8005_ _8028_/CLK _8005_/D vssd1 vssd1 vccd1 vccd1 _8005_/Q sky130_fd_sc_hd__dfxtp_1
Xhold999 _7773_/Q vssd1 vssd1 vccd1 vccd1 hold999/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6266_ _6266_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6266_/X sky130_fd_sc_hd__or2_1
X_6197_ _6040_/X _6196_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6197_/X sky130_fd_sc_hd__mux2_1
Xhold1600 _4169_/Y vssd1 vssd1 vccd1 vccd1 _5553_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4486__S _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5217_ _6963_/A _5188_/B _5220_/B1 hold467/X vssd1 vssd1 vccd1 vccd1 _5217_/X sky130_fd_sc_hd__a22o_1
Xhold1633 _7363_/Q vssd1 vssd1 vccd1 vccd1 hold1633/X sky130_fd_sc_hd__dlygate4sd3_1
X_5148_ _5148_/A1 _4425_/B _5148_/B1 _5147_/X vssd1 vssd1 vccd1 vccd1 _7386_/D sky130_fd_sc_hd__o211a_1
Xhold1611 _7634_/Q vssd1 vssd1 vccd1 vccd1 _4181_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1644 _7657_/Q vssd1 vssd1 vccd1 vccd1 _4343_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1622 _7650_/Q vssd1 vssd1 vccd1 vccd1 _4292_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5079_ _5546_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5079_/X sky130_fd_sc_hd__or2_1
Xhold1655 _7689_/Q vssd1 vssd1 vccd1 vccd1 _3890_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1666 _4299_/Y vssd1 vssd1 vccd1 vccd1 _4300_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1677 _7695_/Q vssd1 vssd1 vccd1 vccd1 _3743_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5623__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1688 _3709_/X vssd1 vssd1 vccd1 vccd1 _6446_/B sky130_fd_sc_hd__buf_1
XANTENNA__6966__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1699 _8497_/Q vssd1 vssd1 vccd1 vccd1 _3856_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4521__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7098__A _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1595_A _3757_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3937__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7248__126 _8354_/CLK vssd1 vssd1 vccd1 vccd1 _8258_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_35_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5065__B _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6103__A1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5512__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6905__A _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6590__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4579__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5776__S0 _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4450_ _4164_/Y _5442_/C _4449_/X _4448_/X vssd1 vssd1 vccd1 vccd1 _8359_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_41_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 _5675_/X vssd1 vssd1 vccd1 vccd1 _7855_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold229 _5337_/X vssd1 vssd1 vccd1 vccd1 _7564_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 _7381_/Q vssd1 vssd1 vccd1 vccd1 _5448_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5696__A3 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4381_ _4377_/A _5468_/C _4380_/X _4379_/X vssd1 vssd1 vccd1 vccd1 _8384_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6120_ _6118_/Y _6119_/X _6391_/A vssd1 vssd1 vccd1 vccd1 _6120_/Y sky130_fd_sc_hd__a21oi_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ _6045_/X _6046_/X _6049_/Y _6050_/Y vssd1 vssd1 vccd1 vccd1 _7879_/D sky130_fd_sc_hd__o31a_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _6551_/A _5465_/B vssd1 vssd1 vccd1 vccd1 _5002_/X sky130_fd_sc_hd__and2_4
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5605__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6948__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6953_ _6953_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6953_/X sky130_fd_sc_hd__and2_1
XFILLER_0_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5904_ _3996_/A _6398_/A2 _6413_/B1 _5889_/A _6011_/A2 vssd1 vssd1 vccd1 vccd1 _5914_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6884_ _7018_/A _6884_/A2 _6906_/A3 _6883_/X vssd1 vssd1 vccd1 vccd1 _6884_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5835_ _6126_/A _5952_/A vssd1 vssd1 vccd1 vccd1 _5836_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5766_ _5765_/B _5765_/C _5765_/A vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5384__A2 _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout326_A _3977_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6550__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6581__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7505_ _7505_/CLK _7505_/D vssd1 vssd1 vccd1 vccd1 _7505_/Q sky130_fd_sc_hd__dfxtp_1
X_5697_ _5695_/X _5696_/X _5879_/S vssd1 vssd1 vccd1 vccd1 _5697_/X sky130_fd_sc_hd__mux2_1
X_4717_ _8161_/Q _7560_/Q _7432_/Q _7592_/Q _4720_/S0 _4731_/S1 vssd1 vssd1 vccd1
+ vccd1 _4717_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_17_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8485_ _8485_/CLK _8485_/D vssd1 vssd1 vccd1 vccd1 _8485_/Q sky130_fd_sc_hd__dfxtp_1
X_7436_ _8458_/CLK _7436_/D vssd1 vssd1 vccd1 vccd1 _7436_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5136__A2 _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4648_ _4646_/X _4647_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4648_/X sky130_fd_sc_hd__mux2_1
Xhold730 _6568_/X vssd1 vssd1 vccd1 vccd1 _8140_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4579_ _8174_/Q _8206_/Q _8270_/Q _7778_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4579_/X sky130_fd_sc_hd__mux4_1
Xhold752 _5204_/X vssd1 vssd1 vccd1 vccd1 _7418_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7367_ _8360_/CLK _7367_/D vssd1 vssd1 vccd1 vccd1 _7367_/Q sky130_fd_sc_hd__dfxtp_1
Xhold763 _7824_/Q vssd1 vssd1 vccd1 vccd1 hold763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 _8479_/Q vssd1 vssd1 vccd1 vccd1 _7021_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 _6713_/X vssd1 vssd1 vccd1 vccd1 _8268_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 _7780_/Q vssd1 vssd1 vccd1 vccd1 hold785/X sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ _6318_/A _6318_/B vssd1 vssd1 vccd1 vccd1 _6319_/B sky130_fd_sc_hd__or2_1
XANTENNA__4990__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold796 _6770_/X vssd1 vssd1 vccd1 vccd1 _8321_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7298_ _8485_/CLK _7298_/D _7108_/Y vssd1 vssd1 vccd1 vccd1 _7298_/Q sky130_fd_sc_hd__dfrtp_4
X_6249_ _6178_/X _6248_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6249_/X sky130_fd_sc_hd__mux2_1
Xhold1441 _7295_/Q vssd1 vssd1 vccd1 vccd1 _5146_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _7284_/Q vssd1 vssd1 vccd1 vccd1 _5124_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1430 hold1798/X vssd1 vssd1 vccd1 vccd1 _4771_/B sky130_fd_sc_hd__buf_2
Xhold1474 _7294_/Q vssd1 vssd1 vccd1 vccd1 _5144_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1485 hold1825/X vssd1 vssd1 vccd1 vccd1 _7031_/A sky130_fd_sc_hd__buf_2
Xhold1463 _8360_/Q vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1496 _6608_/X vssd1 vssd1 vccd1 vccd1 _8168_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5072__A1 input27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6444__B _6444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6021__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6460__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6572__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5507__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5804__A _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6619__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4733__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6635__A _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3861__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3978__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3950_ _5838_/A _5765_/A vssd1 vssd1 vccd1 vccd1 _3950_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3994__A _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3881_ _6262_/A _6259_/A vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__or2_1
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6563__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5620_ _6741_/A _5620_/B vssd1 vssd1 vccd1 vccd1 _5620_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__5997__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6370__A _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5366__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5551_ _6498_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _7740_/D sky130_fd_sc_hd__and2_1
XFILLER_0_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4502_ _5148_/A1 _4241_/C _5451_/C vssd1 vssd1 vccd1 vccd1 _7296_/D sky130_fd_sc_hd__mux2_1
X_8270_ _8270_/CLK _8270_/D vssd1 vssd1 vccd1 vccd1 _8270_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5417__C _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5118__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5482_ _7503_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7671_/D sky130_fd_sc_hd__and3_1
XANTENNA__5749__S0 _5716_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4433_ _5018_/A1 _4432_/Y _5453_/C vssd1 vssd1 vccd1 vccd1 _8365_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4364_ _7057_/A _7735_/Q vssd1 vssd1 vccd1 vccd1 _4367_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_111_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6079__A0 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4972__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7083_ _5546_/A _6975_/C _7080_/X _7083_/B2 vssd1 vssd1 vccd1 vccd1 _7083_/X sky130_fd_sc_hd__a22o_1
X_6103_ _5740_/B _6101_/X _6102_/X _5694_/Y vssd1 vssd1 vccd1 vccd1 _6103_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5433__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4295_ _4295_/A _4295_/B vssd1 vssd1 vccd1 vccd1 _4295_/X sky130_fd_sc_hd__xor2_1
X_6034_ _6035_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _6034_/Y sky130_fd_sc_hd__nand2_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4049__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4724__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout276_A _6908_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7985_ _8370_/CLK _7985_/D vssd1 vssd1 vccd1 vccd1 _7985_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ _7029_/A _6936_/A2 _6943_/B _6935_/X vssd1 vssd1 vccd1 vccd1 _6936_/X sky130_fd_sc_hd__a31o_1
XANTENNA__7079__C _7079_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout443_A _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6867_ _6933_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6867_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6003__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6798_ _7008_/A _6798_/A2 _6779_/B _6797_/X vssd1 vssd1 vccd1 vccd1 _6798_/X sky130_fd_sc_hd__a31o_1
X_5818_ _6144_/S _6094_/B vssd1 vssd1 vccd1 vccd1 _5820_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6280__A _6281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5357__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5749_ _6298_/A _6318_/A _6334_/A _6352_/A _5716_/S _5838_/A vssd1 vssd1 vccd1 vccd1
+ _5750_/B sky130_fd_sc_hd__mux4_1
XANTENNA__6306__A1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4660__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8468_ _8468_/CLK _8468_/D vssd1 vssd1 vccd1 vccd1 _8468_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_114_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8399_ _8475_/CLK _8399_/D vssd1 vssd1 vccd1 vccd1 _8399_/Q sky130_fd_sc_hd__dfxtp_1
X_7419_ _8431_/CLK _7419_/D vssd1 vssd1 vccd1 vccd1 _7419_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4939__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold571 _8224_/Q vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 _5363_/X vssd1 vssd1 vccd1 vccd1 _7590_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6439__B _6439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 _6715_/X vssd1 vssd1 vccd1 vccd1 _8270_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _7548_/Q vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5293__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1260 _6886_/X vssd1 vssd1 vccd1 vccd1 _8409_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 _8430_/Q vssd1 vssd1 vccd1 vccd1 _6930_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1282 _8187_/Q vssd1 vssd1 vccd1 vccd1 _6646_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 _8119_/D vssd1 vssd1 vccd1 vccd1 _8085_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5596__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6190__A _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5348__A2 _5367_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5518__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput109 _7304_/Q vssd1 vssd1 vccd1 vccd1 o_pc_IF[22] sky130_fd_sc_hd__buf_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output72_A _8118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4954__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput91 _8106_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[5] sky130_fd_sc_hd__buf_12
XFILLER_0_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput80 _8125_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[24] sky130_fd_sc_hd__buf_12
XFILLER_0_128_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4080_ _8080_/Q _4079_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _4080_/X sky130_fd_sc_hd__mux2_2
XANTENNA__5284__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4706__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6233__A0 _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6784__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7770_ _8326_/CLK _7770_/D vssd1 vssd1 vccd1 vccd1 _7770_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4982_ _8195_/Q _8227_/Q _8291_/Q _7799_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4982_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_129_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7188__66 _8507_/CLK vssd1 vssd1 vccd1 vccd1 _8101_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3933_ _5789_/S _3934_/B vssd1 vssd1 vccd1 vccd1 _3935_/A sky130_fd_sc_hd__nand2_1
X_6721_ _6937_/A _6705_/B _6738_/B1 hold601/X vssd1 vssd1 vccd1 vccd1 _6721_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6652_ _7022_/A _6652_/A2 _6666_/A3 _6651_/X vssd1 vssd1 vccd1 vccd1 _6652_/X sky130_fd_sc_hd__a31o_1
X_3864_ _4764_/B _4072_/B _3863_/X vssd1 vssd1 vccd1 vccd1 _6441_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5603_ _6877_/A _5584_/B _5617_/B1 hold885/X vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4642__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3795_ _3795_/A1 _4073_/A2 _6947_/A _4073_/B2 _3794_/X vssd1 vssd1 vccd1 vccd1 _3795_/X
+ sky130_fd_sc_hd__a221o_2
X_8322_ _8448_/CLK _8322_/D vssd1 vssd1 vccd1 vccd1 _8322_/Q sky130_fd_sc_hd__dfxtp_1
X_6583_ _6953_/A _6559_/B _6591_/B1 _6583_/B2 vssd1 vssd1 vccd1 vccd1 _6583_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_14_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5534_ _8253_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7723_/D sky130_fd_sc_hd__and3_1
X_5465_ hold65/X _5465_/B _5465_/C vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__and3_1
X_8253_ _8253_/CLK _8253_/D vssd1 vssd1 vccd1 vccd1 _8253_/Q sky130_fd_sc_hd__dfxtp_1
X_8184_ _8346_/CLK _8184_/D vssd1 vssd1 vccd1 vccd1 _8184_/Q sky130_fd_sc_hd__dfxtp_1
X_4416_ _4416_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_111_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout314 _5224_/Y vssd1 vssd1 vccd1 vccd1 _5226_/B sky130_fd_sc_hd__buf_6
X_5396_ _6983_/B _6981_/B vssd1 vssd1 vccd1 vccd1 _6600_/B sky130_fd_sc_hd__and2_1
Xfanout303 _5618_/Y vssd1 vssd1 vccd1 vccd1 _5652_/A2 sky130_fd_sc_hd__buf_6
XANTENNA__6259__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4945__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout347 _3696_/Y vssd1 vssd1 vccd1 vccd1 _3966_/B sky130_fd_sc_hd__buf_4
Xfanout325 _6787_/A vssd1 vssd1 vccd1 vccd1 _6853_/A sky130_fd_sc_hd__buf_4
XANTENNA_fanout393_A _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _3814_/X vssd1 vssd1 vccd1 vccd1 _6965_/A sky130_fd_sc_hd__buf_4
X_4347_ _4346_/X _5058_/A1 _5470_/B vssd1 vssd1 vccd1 vccd1 _4377_/B sky130_fd_sc_hd__mux2_1
X_7066_ _7071_/B _7066_/A2 _7090_/A vssd1 vssd1 vccd1 vccd1 _7066_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout369 _7083_/B2 vssd1 vssd1 vccd1 vccd1 _5474_/A sky130_fd_sc_hd__buf_8
Xfanout358 _4079_/B1 vssd1 vssd1 vccd1 vccd1 _4068_/B1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__5275__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4278_ _8499_/Q _4278_/B vssd1 vssd1 vccd1 vccd1 _4278_/Y sky130_fd_sc_hd__nand2_1
X_6017_ _6017_/A _6017_/B vssd1 vssd1 vccd1 vccd1 _6018_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3825__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7968_ _8096_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 _7968_/Q sky130_fd_sc_hd__dfxtp_1
X_6919_ _6919_/A _6943_/B vssd1 vssd1 vccd1 vccd1 _6919_/X sky130_fd_sc_hd__and2_1
XFILLER_0_77_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7899_ _8454_/CLK _7899_/D vssd1 vssd1 vccd1 vccd1 _7899_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4881__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4002__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4633__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4669__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5073__B _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 _7387_/Q vssd1 vssd1 vccd1 vccd1 _5454_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5266__A1 _6847_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3715__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5520__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3816__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_82_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1090 _6848_/X vssd1 vssd1 vccd1 vccd1 _8390_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6215__A0 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6913__A _6913_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output110_A _7305_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6766__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_97_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_clk_A clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3991__B _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5250_ _6953_/A _5258_/A2 _5258_/B1 hold677/X vssd1 vssd1 vccd1 vccd1 _5250_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_35_clk_A clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4927__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4201_ _8510_/Q _4202_/B vssd1 vssd1 vccd1 vccd1 _4201_/Y sky130_fd_sc_hd__nor2_1
X_5181_ _5470_/A _5470_/C vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4132_ _4132_/A _4132_/B vssd1 vssd1 vccd1 vccd1 _4132_/X sky130_fd_sc_hd__or2_1
XFILLER_0_47_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4756_/B _3676_/A _4082_/B1 _4057_/X _4062_/X vssd1 vssd1 vccd1 vccd1 _6056_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__6807__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5257__A1 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3807__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6757__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6823__A _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7822_ _8218_/CLK _7822_/D vssd1 vssd1 vccd1 vccd1 _7822_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7753_ _8019_/CLK _7753_/D vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4965_ _8353_/Q _7829_/Q _7495_/Q _7463_/Q _4990_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4965_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4863__S0 _4896_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6704_ _6908_/C _6704_/B vssd1 vssd1 vccd1 vccd1 _6706_/B sky130_fd_sc_hd__or2_1
XFILLER_0_117_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3916_ _4746_/B _4083_/B vssd1 vssd1 vccd1 vccd1 _3916_/X sky130_fd_sc_hd__and2_1
XFILLER_0_117_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4896_ _8150_/Q _7549_/Q _7421_/Q _7581_/Q _4896_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4896_/X sky130_fd_sc_hd__mux4_1
XANTENNA_fanout239_A _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5980__A2 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7684_ _8086_/CLK _7684_/D vssd1 vssd1 vccd1 vccd1 _7684_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_108_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4062__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4615__S0 _4741_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6635_ _6941_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6635_/X sky130_fd_sc_hd__and2_1
X_3847_ _6406_/A vssd1 vssd1 vccd1 vccd1 _6405_/A sky130_fd_sc_hd__inv_2
XFILLER_0_132_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6566_ _6853_/A _6592_/A2 _6592_/B1 _6566_/B2 vssd1 vssd1 vccd1 vccd1 _6566_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3778_ _7989_/Q _4068_/A2 _4068_/B1 _8021_/Q _3777_/X vssd1 vssd1 vccd1 vccd1 _3778_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout406_A _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5517_ _8236_/Q _5528_/B _5523_/C vssd1 vssd1 vccd1 vccd1 _7706_/D sky130_fd_sc_hd__and3_1
X_8305_ _8431_/CLK _8305_/D vssd1 vssd1 vccd1 vccd1 _8305_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3743__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8236_ _8236_/CLK _8236_/D vssd1 vssd1 vccd1 vccd1 _8236_/Q sky130_fd_sc_hd__dfxtp_1
X_6497_ _6498_/A _6497_/B vssd1 vssd1 vccd1 vccd1 _6497_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5448_ _5448_/A _5453_/B _5453_/C vssd1 vssd1 vccd1 vccd1 _5448_/X sky130_fd_sc_hd__and3_1
XANTENNA__3738__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6693__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8167_ _8421_/CLK _8167_/D vssd1 vssd1 vccd1 vccd1 _8167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5379_ _6974_/A _6973_/B _5373_/Y vssd1 vssd1 vccd1 vccd1 _5395_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_1_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8098_ _8515_/CLK _8132_/D vssd1 vssd1 vccd1 vccd1 _8098_/Q sky130_fd_sc_hd__dfxtp_1
X_7118_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7118_/Y sky130_fd_sc_hd__inv_2
Xfanout177 _7073_/A vssd1 vssd1 vccd1 vccd1 _7088_/A sky130_fd_sc_hd__buf_4
Xfanout199 _6393_/A vssd1 vssd1 vccd1 vccd1 _6144_/S sky130_fd_sc_hd__buf_4
Xfanout188 _3945_/Y vssd1 vssd1 vccd1 vccd1 _5860_/S sky130_fd_sc_hd__clkbuf_8
Xfanout166 _5002_/X vssd1 vssd1 vccd1 vccd1 _5148_/B1 sky130_fd_sc_hd__buf_6
X_7049_ _7031_/Y _7049_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8497_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__5248__A1 _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6748__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6452__B _6452_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4854__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3982__A1 _3981_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5783__S _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_564 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6920__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6920__B2 _7015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4909__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6684__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6627__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5531__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5239__A1 _6931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4862__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6643__A _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _7007_/A _4750_/B vssd1 vssd1 vccd1 vccd1 _8107_/D sky130_fd_sc_hd__and2_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7158__36 _8472_/CLK vssd1 vssd1 vccd1 vccd1 _8038_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3701_ _7663_/Q _7940_/Q vssd1 vssd1 vccd1 vccd1 _3701_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4681_ _8349_/Q _7825_/Q _7491_/Q _7459_/Q _4734_/S0 _4734_/S1 vssd1 vssd1 vccd1
+ vccd1 _4681_/X sky130_fd_sc_hd__mux4_1
X_6420_ _6534_/A _6420_/B vssd1 vssd1 vccd1 vccd1 _6420_/X sky130_fd_sc_hd__and2_1
XFILLER_0_71_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6351_ _6352_/A _6352_/B vssd1 vssd1 vccd1 vccd1 _6355_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5302_ _3939_/C _5332_/A2 _5332_/B1 hold463/X vssd1 vssd1 vccd1 vccd1 _5302_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6124__C1 _6417_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6282_ _6280_/Y _6282_/B vssd1 vssd1 vccd1 vccd1 _6283_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5233_ _6853_/A _5226_/B _5259_/B1 hold753/X vssd1 vssd1 vccd1 vccd1 _5233_/X sky130_fd_sc_hd__a22o_1
X_8021_ _8096_/CLK _8021_/D vssd1 vssd1 vccd1 vccd1 _8021_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6675__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5164_ _5164_/A1 _4416_/B _5166_/B1 _5163_/X vssd1 vssd1 vccd1 vccd1 _7394_/D sky130_fd_sc_hd__o211a_1
Xhold1804 _7869_/Q vssd1 vssd1 vccd1 vccd1 hold1804/X sky130_fd_sc_hd__dlygate4sd3_1
X_4115_ _4115_/A _4115_/B vssd1 vssd1 vccd1 vccd1 _4115_/X sky130_fd_sc_hd__or2_1
XANTENNA__5441__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1815 _7887_/Q vssd1 vssd1 vccd1 vccd1 hold1815/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6537__B _6537_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5095_ _7057_/A _5463_/C vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__or2_1
X_4046_ _3923_/B _7953_/Q vssd1 vssd1 vccd1 vccd1 _4046_/X sky130_fd_sc_hd__and2b_1
XANTENNA__5650__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7805_ _7805_/CLK _7805_/D vssd1 vssd1 vccd1 vccd1 _7805_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout356_A _6909_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4836__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5997_ _5921_/A _5946_/A _5974_/A _5993_/A _5772_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6080_/B sky130_fd_sc_hd__mux4_1
XFILLER_0_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7736_ _8358_/CLK _7736_/D vssd1 vssd1 vccd1 vccd1 _7736_/Q sky130_fd_sc_hd__dfxtp_1
X_4948_ _8480_/Q _8412_/Q _8444_/Q _8318_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4948_/X sky130_fd_sc_hd__mux4_1
X_7667_ _8388_/CLK _7667_/D vssd1 vssd1 vccd1 vccd1 _7667_/Q sky130_fd_sc_hd__dfxtp_1
X_4879_ _4878_/X _4877_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4879_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3964__B2 _8007_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6618_ _7026_/A _6618_/A2 _6666_/A3 _6617_/X vssd1 vssd1 vccd1 vccd1 _6618_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_7_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5166__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7598_ _8507_/CLK _7598_/D vssd1 vssd1 vccd1 vccd1 _7598_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3716__B2 _8029_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6902__A1 _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7172__50 _8468_/CLK vssd1 vssd1 vccd1 vccd1 _8052_/CLK sky130_fd_sc_hd__inv_2
X_6549_ _7007_/A _6549_/B vssd1 vssd1 vccd1 vccd1 _8031_/D sky130_fd_sc_hd__and2_1
XANTENNA_hold1540_A _7356_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8219_ _8283_/CLK _8219_/D vssd1 vssd1 vccd1 vccd1 _8219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3851__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6447__B _6447_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4248__A _4419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6463__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5641__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5526__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6121__A2 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6409__A0 _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4158__A _4161_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4592__S _4742_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5632__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5920_ _5921_/A _5921_/B vssd1 vssd1 vccd1 vccd1 _5920_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4818__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5851_ _5849_/Y _5850_/X _5734_/A vssd1 vssd1 vccd1 vccd1 _5851_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4802_ _4801_/X _4800_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5782_ _6096_/A _6075_/A _5782_/S vssd1 vssd1 vccd1 vccd1 _5782_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7521_ _7521_/CLK _7521_/D vssd1 vssd1 vccd1 vccd1 _7521_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_56_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4733_ _8196_/Q _8228_/Q _8292_/Q _7800_/Q _4734_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4733_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_16_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5148__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7452_ _8472_/CLK _7452_/D vssd1 vssd1 vccd1 vccd1 _7452_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5699__A1 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6403_ _6406_/A _6406_/B vssd1 vssd1 vccd1 vccd1 _6403_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5436__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4664_ _8476_/Q _8408_/Q _8440_/Q _8314_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4664_/X sky130_fd_sc_hd__mux4_1
X_4595_ _4594_/X _4593_/X _4641_/S vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7383_ _8507_/CLK _7383_/D vssd1 vssd1 vccd1 vccd1 _7383_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold912 _5633_/X vssd1 vssd1 vccd1 vccd1 _7813_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold901 _7555_/Q vssd1 vssd1 vccd1 vccd1 hold901/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _7482_/Q vssd1 vssd1 vccd1 vccd1 hold923/X sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ _6334_/A _6334_/B vssd1 vssd1 vccd1 vccd1 _6335_/B sky130_fd_sc_hd__nor2_1
Xhold945 _7586_/Q vssd1 vssd1 vccd1 vccd1 hold945/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 _6769_/X vssd1 vssd1 vccd1 vccd1 _8320_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 _5350_/X vssd1 vssd1 vccd1 vccd1 _7577_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _7467_/Q vssd1 vssd1 vccd1 vccd1 hold967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 _5218_/X vssd1 vssd1 vccd1 vccd1 _7432_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 _7443_/Q vssd1 vssd1 vccd1 vccd1 hold989/X sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ _6266_/A _6266_/B vssd1 vssd1 vccd1 vccd1 _6265_/Y sky130_fd_sc_hd__nand2_1
X_8004_ _8426_/CLK _8004_/D vssd1 vssd1 vccd1 vccd1 _8004_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5216_ _6961_/A _5188_/B _5220_/B1 hold501/X vssd1 vssd1 vccd1 vccd1 _5216_/X sky130_fd_sc_hd__a22o_1
Xhold1601 _7633_/Q vssd1 vssd1 vccd1 vccd1 _4173_/B sky130_fd_sc_hd__dlygate4sd3_1
X_6196_ _6121_/X _6195_/X _6410_/S vssd1 vssd1 vccd1 vccd1 _6196_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5320__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5147_ _5453_/A _5451_/C vssd1 vssd1 vccd1 vccd1 _5147_/X sky130_fd_sc_hd__or2_1
Xhold1612 _4181_/Y vssd1 vssd1 vccd1 vccd1 _4182_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1634 _7050_/Y vssd1 vssd1 vccd1 vccd1 _7051_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1623 _4292_/Y vssd1 vssd1 vccd1 vccd1 _4293_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5078_ input30/X _5144_/A2 _5146_/B1 _5077_/X vssd1 vssd1 vccd1 vccd1 _7351_/D sky130_fd_sc_hd__o211a_1
Xhold1656 _3890_/X vssd1 vssd1 vccd1 vccd1 _6442_/B sky130_fd_sc_hd__buf_1
Xhold1645 _4344_/B vssd1 vssd1 vccd1 vccd1 _4351_/B1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1667 _4300_/Y vssd1 vssd1 vccd1 vccd1 _4302_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold1678 _7691_/Q vssd1 vssd1 vccd1 vccd1 _3879_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5623__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4426__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4029_ _4029_/A0 _4028_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _6032_/A sky130_fd_sc_hd__mux2_2
Xhold1689 _8512_/Q vssd1 vssd1 vccd1 vccd1 _3982_/A0 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4515__B _5404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1588_A _3904_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3937__B2 _8004_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7719_ _8319_/CLK _7719_/D vssd1 vssd1 vccd1 vccd1 _7719_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5311__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__B _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6654__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7064__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6905__B _6905_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__A1 _6965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4417__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5090__A2 _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4425__B _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6921__A _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4050__B1 _4082_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6132__S _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6590__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold208 _7390_/Q vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 _5448_/X vssd1 vssd1 vccd1 vccd1 _7637_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5776__S1 _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4380_ _4383_/A _4383_/B _4341_/C vssd1 vssd1 vccd1 vccd1 _4380_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6368__A _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6050_ _6050_/A1 _6063_/A _6741_/A vssd1 vssd1 vccd1 vccd1 _6050_/Y sky130_fd_sc_hd__a21oi_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _6534_/A _5001_/B vssd1 vssd1 vccd1 vccd1 _5001_/X sky130_fd_sc_hd__and2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6815__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5605__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4408__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6952_ _7019_/A _6952_/A2 _6943_/B _6951_/X vssd1 vssd1 vccd1 vccd1 _6952_/X sky130_fd_sc_hd__a31o_1
X_5903_ _5881_/C _5902_/Y _5900_/X vssd1 vssd1 vccd1 vccd1 _5903_/X sky130_fd_sc_hd__a21bo_1
X_6883_ _6949_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6883_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5834_ _6410_/S _5834_/B vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__nand2_1
XANTENNA__6831__A _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6030__B2 _6163_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5765_ _5765_/A _5765_/B _5765_/C vssd1 vssd1 vccd1 vccd1 _5765_/X sky130_fd_sc_hd__and3_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6581__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout319_A _4057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5696_ _5921_/A _5870_/A _5946_/A _5892_/A _5804_/A _5789_/S vssd1 vssd1 vccd1 vccd1
+ _5696_/X sky130_fd_sc_hd__mux4_1
XANTENNA_fanout221_A _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4716_ _8354_/Q _7830_/Q _7496_/Q _7464_/Q _4720_/S0 _4741_/S1 vssd1 vssd1 vccd1
+ vccd1 _4716_/X sky130_fd_sc_hd__mux4_1
X_8484_ _8484_/CLK _8484_/D vssd1 vssd1 vccd1 vccd1 _8484_/Q sky130_fd_sc_hd__dfxtp_1
X_7504_ _7504_/CLK _7504_/D vssd1 vssd1 vccd1 vccd1 _7504_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7435_ _8487_/CLK _7435_/D vssd1 vssd1 vccd1 vccd1 _7435_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4070__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4647_ _8151_/Q _7550_/Q _7422_/Q _7582_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4647_/X sky130_fd_sc_hd__mux4_1
Xhold720 _7008_/X vssd1 vssd1 vccd1 vccd1 _8466_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7142__20 _8445_/CLK vssd1 vssd1 vccd1 vccd1 _7519_/CLK sky130_fd_sc_hd__inv_2
X_7366_ _8480_/CLK _7366_/D vssd1 vssd1 vccd1 vccd1 _7366_/Q sky130_fd_sc_hd__dfxtp_1
Xhold731 _8464_/Q vssd1 vssd1 vccd1 vccd1 _7006_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _4576_/X _4577_/X _5473_/A vssd1 vssd1 vccd1 vccd1 _4578_/X sky130_fd_sc_hd__mux2_1
Xhold753 _7441_/Q vssd1 vssd1 vccd1 vccd1 hold753/X sky130_fd_sc_hd__dlygate4sd3_1
X_6317_ _6318_/A _6318_/B vssd1 vssd1 vccd1 vccd1 _6317_/Y sky130_fd_sc_hd__nor2_1
Xhold764 _5644_/X vssd1 vssd1 vccd1 vccd1 _7824_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 _7021_/X vssd1 vssd1 vccd1 vccd1 _8479_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6884__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold786 _5596_/X vssd1 vssd1 vccd1 vccd1 _7780_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 _7438_/Q vssd1 vssd1 vccd1 vccd1 hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 _8286_/Q vssd1 vssd1 vccd1 vccd1 hold797/X sky130_fd_sc_hd__dlygate4sd3_1
X_7297_ _8480_/CLK _7297_/D _7107_/Y vssd1 vssd1 vccd1 vccd1 _7297_/Q sky130_fd_sc_hd__dfrtp_4
X_6248_ _6191_/A _6209_/A _6226_/A _6244_/A _3928_/X _5804_/A vssd1 vssd1 vccd1 vccd1
+ _6248_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6636__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6179_ _6099_/X _6178_/X _6393_/A vssd1 vssd1 vccd1 vccd1 _6179_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1420 _7659_/Q vssd1 vssd1 vccd1 vccd1 _4356_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1503_A _7297_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1431 _8371_/Q vssd1 vssd1 vccd1 vccd1 _5030_/A1 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold1442 _7303_/Q vssd1 vssd1 vccd1 vccd1 _5162_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 _7287_/Q vssd1 vssd1 vccd1 vccd1 _5130_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 _7030_/X vssd1 vssd1 vccd1 vccd1 _8488_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 _7305_/Q vssd1 vssd1 vccd1 vccd1 _5166_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 _7308_/Q vssd1 vssd1 vccd1 vccd1 _5172_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1497 _7732_/Q vssd1 vssd1 vccd1 vccd1 _5654_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5072__A2 _4448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6741__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4960__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6572__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5780__A0 _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6088__A1 _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5523__C _5523_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7037__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6635__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5599__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6651__A _6891_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_70_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _8515_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3880_ _3880_/A0 _6444_/B _4074_/S vssd1 vssd1 vccd1 vccd1 _6259_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4023__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5997__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5550_ _7006_/A _5550_/B vssd1 vssd1 vccd1 vccd1 _5550_/X sky130_fd_sc_hd__and2_1
X_5481_ _7502_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7670_/D sky130_fd_sc_hd__and3_1
XFILLER_0_81_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6377__A1_N _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4501_ _5150_/A1 _4415_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _7297_/D sky130_fd_sc_hd__mux2_1
X_4432_ _4432_/A _4432_/B vssd1 vssd1 vccd1 vccd1 _4432_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5749__S1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6866__A3 _6906_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ _5475_/A _7732_/Q vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__xor2_1
XANTENNA__6079__A1 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7082_ _7082_/A _7082_/B _7082_/C vssd1 vssd1 vccd1 vccd1 _8515_/D sky130_fd_sc_hd__and3_1
X_6102_ _5925_/B _5938_/X _6250_/S vssd1 vssd1 vccd1 vccd1 _6102_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6618__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5433__C _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4294_ _4284_/Y _4288_/B _4285_/Y vssd1 vssd1 vccd1 vccd1 _4295_/B sky130_fd_sc_hd__o21a_1
X_6033_ _6035_/A _6035_/B vssd1 vssd1 vccd1 vccd1 _6036_/A sky130_fd_sc_hd__and2_1
XANTENNA__5826__B2 _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7984_ _8034_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 _7984_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout171_A _7030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6935_ _6935_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6935_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout269_A _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5054__A2 _5069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5876__S _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _8370_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6866_ _7023_/A _6866_/A2 _6906_/A3 _6865_/X vssd1 vssd1 vccd1 vccd1 _6866_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout436_A _7027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6797_ _6929_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6797_/X sky130_fd_sc_hd__and2_1
X_5817_ _5765_/X _5769_/B _5767_/B vssd1 vssd1 vccd1 vccd1 _5823_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_57_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5748_ _6270_/A _5748_/B vssd1 vssd1 vccd1 vccd1 _5748_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4660__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1453_A _7287_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8467_ _8467_/CLK _8467_/D vssd1 vssd1 vccd1 vccd1 _8467_/Q sky130_fd_sc_hd__dfxtp_1
X_5679_ _6545_/A _5679_/B vssd1 vssd1 vccd1 vccd1 _5679_/X sky130_fd_sc_hd__and2_1
XFILLER_0_130_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8398_ _8466_/CLK _8398_/D vssd1 vssd1 vccd1 vccd1 _8398_/Q sky130_fd_sc_hd__dfxtp_1
X_7418_ _8154_/CLK _7418_/D vssd1 vssd1 vccd1 vccd1 _7418_/Q sky130_fd_sc_hd__dfxtp_1
X_7349_ _8519_/CLK _7349_/D vssd1 vssd1 vccd1 vccd1 _7349_/Q sky130_fd_sc_hd__dfxtp_1
Xhold561 _7579_/Q vssd1 vssd1 vccd1 vccd1 hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 _6697_/X vssd1 vssd1 vccd1 vccd1 _8224_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _5254_/X vssd1 vssd1 vccd1 vccd1 _7462_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _5317_/X vssd1 vssd1 vccd1 vccd1 _7548_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _8278_/Q vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3828__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5293__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1250 _6860_/X vssd1 vssd1 vccd1 vccd1 _8396_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1261 _8450_/Q vssd1 vssd1 vccd1 vccd1 _6970_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 _6930_/X vssd1 vssd1 vccd1 vccd1 _8430_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1283 _6646_/X vssd1 vssd1 vccd1 vccd1 _8187_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 _8345_/Q vssd1 vssd1 vccd1 vccd1 _6816_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4690__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_52_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8457_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6471__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5087__A _7065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5518__C _7073_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6848__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5534__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput70 _8116_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[15] sky130_fd_sc_hd__buf_12
Xoutput81 _8126_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[25] sky130_fd_sc_hd__buf_12
XANTENNA__4865__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput92 _8107_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[6] sky130_fd_sc_hd__buf_12
XANTENNA_output65_A _8111_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5550__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5284__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3989__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6233__A1 _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5036__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6784__A2 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4981_ _4979_/X _4980_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_43_clk _7871_/CLK vssd1 vssd1 vccd1 vccd1 _8328_/CLK sky130_fd_sc_hd__clkbuf_16
X_6720_ _6935_/A _6705_/B _6738_/B1 _6720_/B2 vssd1 vssd1 vccd1 vccd1 _6720_/X sky130_fd_sc_hd__a22o_1
X_3932_ _3934_/B vssd1 vssd1 vccd1 vccd1 _4094_/B sky130_fd_sc_hd__inv_2
XFILLER_0_19_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6651_ _6891_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6651_/X sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_9_clk_A clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3863_ _3863_/A1 _4073_/A2 _6949_/A _4073_/B2 vssd1 vssd1 vccd1 vccd1 _3863_/X sky130_fd_sc_hd__a22o_1
X_6582_ _6951_/A _6592_/A2 _6592_/B1 hold943/X vssd1 vssd1 vccd1 vccd1 _6582_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5744__A0 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5602_ _6941_/A _5584_/B _5617_/B1 hold779/X vssd1 vssd1 vccd1 vccd1 _5602_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5428__C _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4642__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3794_ _4763_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__and2_1
XFILLER_0_54_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5533_ _8252_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7722_/D sky130_fd_sc_hd__and3_1
XFILLER_0_5_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8321_ _8483_/CLK _8321_/D vssd1 vssd1 vccd1 vccd1 _8321_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8252_ _8252_/CLK _8252_/D vssd1 vssd1 vccd1 vccd1 _8252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5464_ _5464_/A _5465_/B _5465_/C vssd1 vssd1 vccd1 vccd1 _5464_/X sky130_fd_sc_hd__and3_1
XFILLER_0_111_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8183_ _8473_/CLK _8183_/D vssd1 vssd1 vccd1 vccd1 _8183_/Q sky130_fd_sc_hd__dfxtp_1
X_5395_ _5395_/A _7055_/B _7071_/A _5409_/A vssd1 vssd1 vccd1 vccd1 _6981_/B sky130_fd_sc_hd__or4b_1
XANTENNA__5444__B _7082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4415_ _4419_/A _4415_/B vssd1 vssd1 vccd1 vccd1 _4415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout304 _5618_/Y vssd1 vssd1 vccd1 vccd1 _5620_/B sky130_fd_sc_hd__buf_6
X_4346_ _4346_/A _4346_/B vssd1 vssd1 vccd1 vccd1 _4346_/X sky130_fd_sc_hd__xor2_1
Xfanout315 _5186_/Y vssd1 vssd1 vccd1 vccd1 _5188_/B sky130_fd_sc_hd__buf_6
Xfanout348 _3683_/X vssd1 vssd1 vccd1 vccd1 _6959_/A sky130_fd_sc_hd__buf_4
Xfanout337 _3803_/X vssd1 vssd1 vccd1 vccd1 _6969_/A sky130_fd_sc_hd__buf_4
Xfanout326 _3977_/X vssd1 vssd1 vccd1 vccd1 _6923_/A sky130_fd_sc_hd__buf_4
X_7065_ _7065_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7065_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout359 _3681_/X vssd1 vssd1 vccd1 vccd1 _4079_/B1 sky130_fd_sc_hd__buf_8
X_4277_ _4277_/A _4278_/B vssd1 vssd1 vccd1 vccd1 _4277_/Y sky130_fd_sc_hd__nor2_1
X_6016_ _6016_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6017_/B sky130_fd_sc_hd__or2_1
XANTENNA__5275__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7967_ _8500_/CLK hold62/X vssd1 vssd1 vccd1 vccd1 _7967_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_34_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8143_/CLK sky130_fd_sc_hd__clkbuf_16
X_7898_ _8419_/CLK _7898_/D vssd1 vssd1 vccd1 vccd1 _7898_/Q sky130_fd_sc_hd__dfxtp_1
X_6918_ _7024_/A _6918_/A2 _6970_/A3 _6917_/X vssd1 vssd1 vccd1 vccd1 _6918_/X sky130_fd_sc_hd__a31o_1
X_6849_ _6849_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6849_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4881__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5735__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1570_A _7370_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4633__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5830__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8519_ _8519_/CLK _8519_/D vssd1 vssd1 vccd1 vccd1 _8519_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3761__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6160__A0 _6140_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold380 _7330_/Q vssd1 vssd1 vccd1 vccd1 _5427_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold391 _5454_/X vssd1 vssd1 vccd1 vccd1 _7643_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6466__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5370__A _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5266__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5018__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1080 _6620_/X vssd1 vssd1 vccd1 vccd1 _8174_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6215__A1 _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1091 _8281_/Q vssd1 vssd1 vccd1 vccd1 _6726_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6913__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6766__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8461_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output103_A _7298_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5529__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4200_ _4435_/B _4200_/B vssd1 vssd1 vccd1 vccd1 _4432_/A sky130_fd_sc_hd__nand2b_1
X_5180_ _5180_/A1 _5182_/A2 _5182_/B1 _5179_/X vssd1 vssd1 vccd1 vccd1 _7402_/D sky130_fd_sc_hd__o211a_1
XANTENNA__4595__S _4641_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4131_ _3896_/A _4130_/X _4129_/Y vssd1 vssd1 vccd1 vccd1 _4132_/B sky130_fd_sc_hd__o21a_1
X_4062_ _4062_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _4062_/X sky130_fd_sc_hd__or2_1
XANTENNA__5257__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6757__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7821_ _8445_/CLK _7821_/D vssd1 vssd1 vccd1 vccd1 _7821_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6823__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7752_ _8370_/CLK _7752_/D vssd1 vssd1 vccd1 vccd1 _7752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_16_clk _7871_/CLK vssd1 vssd1 vccd1 vccd1 _8469_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_74_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4964_ _4963_/X _4960_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8256_/D sky130_fd_sc_hd__mux2_1
XANTENNA__7000__A _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4863__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6703_ _6908_/C _6704_/B vssd1 vssd1 vccd1 vccd1 _6703_/Y sky130_fd_sc_hd__nor2_4
X_3915_ _4746_/B _3669_/Y _4082_/B1 _6847_/A _3914_/X vssd1 vssd1 vccd1 vccd1 _5820_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_58_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5439__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4895_ _8343_/Q _7819_/Q _7485_/Q _7453_/Q _4895_/S0 _4896_/S1 vssd1 vssd1 vccd1
+ vccd1 _4895_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_62_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7683_ _8450_/CLK _7683_/D vssd1 vssd1 vccd1 vccd1 _7683_/Q sky130_fd_sc_hd__dfxtp_1
X_3846_ _3846_/A _3846_/B vssd1 vssd1 vccd1 vccd1 _6406_/A sky130_fd_sc_hd__nand2_1
X_6634_ _7023_/A _6634_/A2 _6666_/A3 _6633_/X vssd1 vssd1 vccd1 vccd1 _6634_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5193__A1 _6849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4615__S1 _4737_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3777_ _4067_/A_N _7957_/Q vssd1 vssd1 vccd1 vccd1 _3777_/X sky130_fd_sc_hd__and2b_1
X_6565_ _6917_/A _6559_/B _6591_/B1 _6565_/B2 vssd1 vssd1 vccd1 vccd1 _6565_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_132_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8304_ _8462_/CLK _8304_/D vssd1 vssd1 vccd1 vccd1 _8304_/Q sky130_fd_sc_hd__dfxtp_1
X_5516_ _8235_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7705_/D sky130_fd_sc_hd__and3_1
X_6496_ _6520_/A _6496_/B vssd1 vssd1 vccd1 vccd1 _6496_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout301_A _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3743__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5447_ _5447_/A _7073_/A _5449_/C vssd1 vssd1 vccd1 vccd1 _5447_/X sky130_fd_sc_hd__and3_1
X_8235_ _8235_/CLK _8235_/D vssd1 vssd1 vccd1 vccd1 _8235_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__6693__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8166_ _8421_/CLK _8166_/D vssd1 vssd1 vccd1 vccd1 _8166_/Q sky130_fd_sc_hd__dfxtp_1
X_5378_ _6553_/A _6553_/B vssd1 vssd1 vccd1 vccd1 _6973_/B sky130_fd_sc_hd__and2b_1
X_8097_ _8419_/CLK _8131_/D vssd1 vssd1 vccd1 vccd1 _8097_/Q sky130_fd_sc_hd__dfxtp_1
X_4329_ _8492_/Q _4329_/B vssd1 vssd1 vccd1 vccd1 _4329_/Y sky130_fd_sc_hd__nand2_1
X_7117_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7117_/Y sky130_fd_sc_hd__inv_2
Xfanout178 _7073_/A vssd1 vssd1 vccd1 vccd1 _5453_/B sky130_fd_sc_hd__buf_4
Xfanout189 _3945_/Y vssd1 vssd1 vccd1 vccd1 _5804_/A sky130_fd_sc_hd__buf_4
Xfanout167 hold1510/X vssd1 vssd1 vccd1 vccd1 _5538_/B sky130_fd_sc_hd__buf_4
X_7048_ _7048_/A _7055_/B vssd1 vssd1 vccd1 vccd1 _7048_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5248__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4518__B _5408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6986__A_N _7354_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4551__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6748__A2 _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4854__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5708__A0 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6920__A2 _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4790__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5531__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5239__A2 _5258_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4542__S0 _4611_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6643__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3700_ _7663_/Q _7940_/Q vssd1 vssd1 vccd1 vccd1 _3700_/Y sky130_fd_sc_hd__nand2_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680_ _4679_/X _4676_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7522_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_126_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6350_ _6350_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6352_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5301_ _6777_/A _5300_/B _5300_/Y hold264/X vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5733__A_N _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6124__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6281_ _6281_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6282_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _8475_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6675__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8020_ _8020_/CLK _8020_/D vssd1 vssd1 vccd1 vccd1 _8020_/Q sky130_fd_sc_hd__dfxtp_1
X_5232_ _6917_/A _5258_/A2 _5258_/B1 hold859/X vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__a22o_1
X_5163_ _5461_/A _5540_/C vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__or2_1
Xhold1805 _7352_/Q vssd1 vssd1 vccd1 vccd1 hold1805/X sky130_fd_sc_hd__dlygate4sd3_1
X_4114_ _4090_/A _4113_/X _4112_/Y vssd1 vssd1 vccd1 vccd1 _4115_/B sky130_fd_sc_hd__o21a_1
Xhold1816 _7889_/Q vssd1 vssd1 vccd1 vccd1 hold1816/X sky130_fd_sc_hd__dlygate4sd3_1
X_5094_ input8/X _5144_/A2 _5146_/B1 _5093_/X vssd1 vssd1 vccd1 vccd1 _7359_/D sky130_fd_sc_hd__o211a_1
X_4045_ _4045_/A _4045_/B _4109_/A _4045_/D vssd1 vssd1 vccd1 vccd1 _4045_/X sky130_fd_sc_hd__or4_1
XANTENNA__5650__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7804_ _8136_/CLK _7804_/D vssd1 vssd1 vccd1 vccd1 _7804_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4836__S1 _7358_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5996_ _5996_/A _5996_/B vssd1 vssd1 vccd1 vccd1 _5996_/X sky130_fd_sc_hd__xor2_1
XANTENNA_fanout349_A _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5169__B _5465_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7735_ _7907_/CLK _7735_/D vssd1 vssd1 vccd1 vccd1 _7735_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4947_ _8190_/Q _8222_/Q _8286_/Q _7794_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4947_/X sky130_fd_sc_hd__mux4_1
X_7666_ _8421_/CLK _7666_/D vssd1 vssd1 vccd1 vccd1 _7666_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_117_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4878_ _8470_/Q _8402_/Q _8434_/Q _8308_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4878_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_62_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3964__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6363__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6617_ _6923_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6617_/X sky130_fd_sc_hd__and2_1
X_3829_ _3829_/A1 _4073_/A2 _3826_/X _4073_/B2 vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3716__A2 _4068_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7597_ _8090_/CLK _7597_/D vssd1 vssd1 vccd1 vccd1 _7597_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6548_ _6548_/A _6548_/B vssd1 vssd1 vccd1 vccd1 _8030_/D sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_81_clk_A clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6479_ _6550_/A _6479_/B vssd1 vssd1 vccd1 vccd1 _6479_/X sky130_fd_sc_hd__and2_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6666__A1 _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8218_ _8218_/CLK _8218_/D vssd1 vssd1 vccd1 vccd1 _8218_/Q sky130_fd_sc_hd__dfxtp_1
X_8149_ _8413_/CLK _8149_/D vssd1 vssd1 vccd1 vccd1 _8149_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_96_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4524__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4963__S _4991_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5641__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_34_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_49_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5095__A _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5526__C _5541_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6106__B1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5865__C1 _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5542__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6409__A1 _6352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_107_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3891__A1 _3890_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4873__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5632__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7218__96 _8419_/CLK vssd1 vssd1 vccd1 vccd1 _8131_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6290__C1 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6356__B1_N _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6268__S0 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5850_ _5850_/A _5850_/B vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__or2_1
XANTENNA__6042__C1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4818__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4801_ _8459_/Q _8391_/Q _8423_/Q _8297_/Q _4896_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4801_/X sky130_fd_sc_hd__mux4_1
X_5781_ _6140_/A _6115_/A _5782_/S vssd1 vssd1 vccd1 vccd1 _5781_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4732_ _4730_/X _4731_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__mux2_1
X_7520_ _7520_/CLK _7520_/D vssd1 vssd1 vccd1 vccd1 _7520_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_29_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6345__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4663_ _8186_/Q _8218_/Q _8282_/Q _7790_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4663_/X sky130_fd_sc_hd__mux4_1
X_7451_ _8471_/CLK _7451_/D vssd1 vssd1 vccd1 vccd1 _7451_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5699__A2 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6402_ _6390_/A _6387_/X _6389_/B vssd1 vssd1 vccd1 vccd1 _6402_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__6896__A1 _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4594_ _8466_/Q _8398_/Q _8430_/Q _8304_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4594_/X sky130_fd_sc_hd__mux4_1
X_7382_ _8510_/CLK _7382_/D vssd1 vssd1 vccd1 vccd1 _7382_/Q sky130_fd_sc_hd__dfxtp_1
Xhold913 _8474_/Q vssd1 vssd1 vccd1 vccd1 _7016_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold902 _5324_/X vssd1 vssd1 vccd1 vccd1 _7555_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold924 _5278_/X vssd1 vssd1 vccd1 vccd1 _7482_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 _8481_/Q vssd1 vssd1 vccd1 vccd1 _7023_/B sky130_fd_sc_hd__dlygate4sd3_1
X_6333_ _6334_/A _6334_/B vssd1 vssd1 vccd1 vccd1 _6333_/Y sky130_fd_sc_hd__nand2_1
Xhold946 _5359_/X vssd1 vssd1 vccd1 vccd1 _7586_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6829__A _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold979 _7481_/Q vssd1 vssd1 vccd1 vccd1 hold979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 _5259_/X vssd1 vssd1 vccd1 vccd1 _7467_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _7551_/Q vssd1 vssd1 vccd1 vccd1 hold957/X sky130_fd_sc_hd__dlygate4sd3_1
X_6264_ _6247_/A _6246_/A _6245_/A vssd1 vssd1 vccd1 vccd1 _6266_/B sky130_fd_sc_hd__a21o_1
XANTENNA__6648__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8003_ _8034_/CLK _8003_/D vssd1 vssd1 vccd1 vccd1 _8003_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5452__B _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5215_ _6959_/A _5221_/A2 _5221_/B1 hold759/X vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5320__A1 _6947_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_15_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout299_A _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6195_ _6140_/A _6157_/A _6175_/A _6191_/A _5782_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _6195_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5146_ _5146_/A1 _4425_/B _5146_/B1 _5145_/X vssd1 vssd1 vccd1 vccd1 _7385_/D sky130_fd_sc_hd__o211a_1
Xhold1635 _7681_/Q vssd1 vssd1 vccd1 vccd1 _4084_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1613 _4189_/X vssd1 vssd1 vccd1 vccd1 _4190_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1602 _4173_/Y vssd1 vssd1 vccd1 vccd1 _4174_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1624 _4293_/Y vssd1 vssd1 vccd1 vccd1 _4295_/A sky130_fd_sc_hd__dlygate4sd3_1
X_5077_ _5545_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5077_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout466_A _6911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1657 _7696_/Q vssd1 vssd1 vccd1 vccd1 _3816_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1646 _4351_/X vssd1 vssd1 vccd1 vccd1 _4352_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1668 _4302_/Y vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5084__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5623__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6820__A1 _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4028_ _4028_/A1 _4073_/A2 _6931_/A _4073_/B2 _4027_/X vssd1 vssd1 vccd1 vccd1 _4028_/X
+ sky130_fd_sc_hd__a221o_2
Xhold1679 _7687_/Q vssd1 vssd1 vccd1 vccd1 _3795_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5979_ _4021_/A _5731_/Y _6413_/B1 _4020_/A _6011_/A2 vssd1 vssd1 vccd1 vccd1 _5979_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6584__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7718_ _8486_/CLK _7718_/D vssd1 vssd1 vccd1 vccd1 _7718_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold1650_A _7055_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7649_ _8091_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 _7649_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4993__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3862__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4033__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A1 _6929_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__S _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7064__A1 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6474__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4693__S _7048_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5614__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6921__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6575__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3928__A2 _6421_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5537__B _5538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6878__A1 _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold209 _5457_/X vssd1 vssd1 vccd1 vccd1 _7646_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6649__A _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5553__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__A1 _3939_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5000_ _6534_/A _5000_/B vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__and2_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3864__A1 _4764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6802__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5066__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5605__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6951_ _6951_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6951_/X sky130_fd_sc_hd__and2_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5902_ _6270_/A _5901_/X _5900_/B vssd1 vssd1 vccd1 vccd1 _5902_/Y sky130_fd_sc_hd__a21oi_1
X_6882_ _7017_/A _6882_/A2 _6906_/A3 _6881_/X vssd1 vssd1 vccd1 vccd1 _6882_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_48_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6566__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5833_ _6334_/A _6352_/A _6370_/A _6388_/A _5744_/S _5859_/S vssd1 vssd1 vccd1 vccd1
+ _5834_/B sky130_fd_sc_hd__mux4_1
XANTENNA__6831__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3919__A2 _3917_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5728__A _5734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7503_ _7503_/CLK _7503_/D vssd1 vssd1 vccd1 vccd1 _7503_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5447__B _7073_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5764_ _5763_/A _5763_/B _5971_/B vssd1 vssd1 vccd1 vccd1 _5765_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5695_ _5846_/A _5820_/A _5765_/A _3934_/B _5772_/S _5804_/A vssd1 vssd1 vccd1 vccd1
+ _5695_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8483_ _8483_/CLK _8483_/D vssd1 vssd1 vccd1 vccd1 _8483_/Q sky130_fd_sc_hd__dfxtp_1
X_4715_ _4714_/X _4711_/X _7046_/A vssd1 vssd1 vccd1 vccd1 _7527_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7434_ _8448_/CLK _7434_/D vssd1 vssd1 vccd1 vccd1 _7434_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4646_ _8344_/Q _7820_/Q _7486_/Q _7454_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4646_/X sky130_fd_sc_hd__mux4_1
XANTENNA_fanout214_A _5456_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4778__S _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4577_ _8141_/Q _7540_/Q _7412_/Q _7572_/Q _7072_/B2 _7050_/A vssd1 vssd1 vccd1 vccd1
+ _4577_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6559__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7365_ _8461_/CLK _7365_/D vssd1 vssd1 vccd1 vccd1 _7365_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4975__S0 _7063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold710 _5652_/X vssd1 vssd1 vccd1 vccd1 _7832_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold721 _8460_/Q vssd1 vssd1 vccd1 vccd1 _7002_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 _7006_/X vssd1 vssd1 vccd1 vccd1 _8464_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 _5233_/X vssd1 vssd1 vccd1 vccd1 _7441_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 _8470_/Q vssd1 vssd1 vccd1 vccd1 _7012_/B sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ _6318_/A _6318_/B vssd1 vssd1 vccd1 vccd1 _6319_/A sky130_fd_sc_hd__nand2_1
X_7296_ _8368_/CLK _7296_/D _7106_/Y vssd1 vssd1 vccd1 vccd1 _7296_/Q sky130_fd_sc_hd__dfrtp_2
Xhold787 _7474_/Q vssd1 vssd1 vccd1 vccd1 hold787/X sky130_fd_sc_hd__dlygate4sd3_1
X_3662__1 _8388_/CLK vssd1 vssd1 vccd1 vccd1 _7500_/CLK sky130_fd_sc_hd__inv_2
Xhold776 _5230_/X vssd1 vssd1 vccd1 vccd1 _7438_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5829__C1 _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold765 _7781_/Q vssd1 vssd1 vccd1 vccd1 hold765/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6247_ _6247_/A _6247_/B vssd1 vssd1 vccd1 vccd1 _6247_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold798 _6731_/X vssd1 vssd1 vccd1 vccd1 _8286_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4727__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6178_ _6140_/A _6175_/A _6115_/A _6157_/A _5860_/S _5744_/S vssd1 vssd1 vccd1 vccd1
+ _6178_/X sky130_fd_sc_hd__mux4_1
Xhold1410 _4267_/X vssd1 vssd1 vccd1 vccd1 _5567_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1443 hold1806/X vssd1 vssd1 vccd1 vccd1 _7074_/A sky130_fd_sc_hd__buf_2
X_5129_ _5444_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5129_/X sky130_fd_sc_hd__or2_1
Xhold1421 _4356_/X vssd1 vssd1 vccd1 vccd1 _4357_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1432 hold1802/X vssd1 vssd1 vccd1 vccd1 _4766_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3855__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1476 _7293_/Q vssd1 vssd1 vccd1 vccd1 _5142_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1465 _7312_/Q vssd1 vssd1 vccd1 vccd1 _5180_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 _7302_/Q vssd1 vssd1 vccd1 vccd1 _5160_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold1498 _7288_/Q vssd1 vssd1 vccd1 vccd1 _5132_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1487 hold1501/X vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1698_A _4073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6021__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6741__B _6741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5780__A1 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6469__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4966__S0 _4990_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6188__B _6405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5048__B1 _5166_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3767__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5548__A _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6651__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5068__C_N _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4023__B2 _8014_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5220__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5771__A1 _6105_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5480_ _7501_/Q _7088_/A _7088_/B vssd1 vssd1 vccd1 vccd1 _7669_/D sky130_fd_sc_hd__and3_1
XFILLER_0_53_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4500_ _5152_/A1 _4413_/B _5454_/C vssd1 vssd1 vccd1 vccd1 _7298_/D sky130_fd_sc_hd__mux2_1
X_4431_ _5020_/A1 _4430_/Y _5451_/C vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_1 _7694_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6720__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4362_ _3648_/Y _7734_/Q _7735_/Q _3647_/Y _4359_/Y vssd1 vssd1 vccd1 vccd1 _4362_/Y
+ sky130_fd_sc_hd__o221ai_1
XFILLER_0_6_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7081_ _5081_/A _6975_/C _7080_/X _7044_/A vssd1 vssd1 vccd1 vccd1 _7082_/C sky130_fd_sc_hd__a22o_1
XANTENNA__6079__A2 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6101_ _5936_/B _6100_/X _6342_/S vssd1 vssd1 vccd1 vccd1 _6101_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4709__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4293_ _4291_/Y _4293_/B vssd1 vssd1 vccd1 vccd1 _4293_/Y sky130_fd_sc_hd__nand2b_1
X_6032_ _6032_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6035_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__5826__A2 _6380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5287__B1 _5294_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7238__116 _8450_/CLK vssd1 vssd1 vccd1 vccd1 _8248_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__7003__A _7019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6236__C1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7983_ _8369_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 _7983_/Q sky130_fd_sc_hd__dfxtp_1
X_6934_ _7007_/A _6934_/A2 _6943_/B _6933_/X vssd1 vssd1 vccd1 vccd1 _6934_/X sky130_fd_sc_hd__a31o_1
XANTENNA_fanout164_A _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6003__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6865_ _6931_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6865_/X sky130_fd_sc_hd__and2_1
XANTENNA__5211__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6796_ _7007_/A _6796_/A2 _6779_/B _6795_/X vssd1 vssd1 vccd1 vccd1 _6796_/X sky130_fd_sc_hd__a31o_1
X_7202__80 _8469_/CLK vssd1 vssd1 vccd1 vccd1 _8115_/CLK sky130_fd_sc_hd__inv_2
X_5816_ _5811_/X _5815_/X _6412_/S vssd1 vssd1 vccd1 vccd1 _5816_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout429_A _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4081__B _4081_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5747_ _5745_/X _5746_/X _5950_/S vssd1 vssd1 vccd1 vccd1 _5748_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_45_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_8466_ _8466_/CLK _8466_/D vssd1 vssd1 vccd1 vccd1 _8466_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7417_ _8473_/CLK _7417_/D vssd1 vssd1 vccd1 vccd1 _7417_/Q sky130_fd_sc_hd__dfxtp_1
X_5678_ _6550_/A hold27/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__and2_1
XFILLER_0_130_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3706__A _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8397_ _8465_/CLK _8397_/D vssd1 vssd1 vccd1 vccd1 _8397_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6711__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4948__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4629_ _8471_/Q _8403_/Q _8435_/Q _8309_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4629_/X sky130_fd_sc_hd__mux4_1
Xhold551 _8271_/Q vssd1 vssd1 vccd1 vccd1 hold551/X sky130_fd_sc_hd__dlygate4sd3_1
X_7348_ _7977_/CLK _7348_/D vssd1 vssd1 vccd1 vccd1 _7348_/Q sky130_fd_sc_hd__dfxtp_1
Xhold562 _5352_/X vssd1 vssd1 vccd1 vccd1 _7579_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _5609_/X vssd1 vssd1 vccd1 vccd1 _7793_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _7448_/Q vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _8207_/Q vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6110__B1_N _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold584 _6723_/X vssd1 vssd1 vccd1 vccd1 _8278_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7279_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7279_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5921__A _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5278__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3828__A1 _4773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3828__B2 _6967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1251 _8186_/Q vssd1 vssd1 vccd1 vccd1 _6644_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1240 _6874_/X vssd1 vssd1 vccd1 vccd1 _8403_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 hold1814/X vssd1 vssd1 vccd1 vccd1 _7077_/A sky130_fd_sc_hd__clkbuf_2
Xhold1284 _8445_/Q vssd1 vssd1 vccd1 vccd1 _6960_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1262 _6970_/X vssd1 vssd1 vccd1 vccd1 _8450_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1295 _6816_/X vssd1 vssd1 vccd1 vccd1 _8345_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4971__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5202__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4005__A1 _4004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5087__B _5451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5753__A1 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3939__A_N _4083_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6702__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5534__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6927__A _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput93 _8108_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[7] sky130_fd_sc_hd__buf_12
Xoutput71 _8117_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[16] sky130_fd_sc_hd__buf_12
XFILLER_0_128_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5269__B1 _5295_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput82 _8127_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[26] sky130_fd_sc_hd__buf_12
XFILLER_0_37_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6769__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6233__A2 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4980_ _8162_/Q _7561_/Q _7433_/Q _7593_/Q _4983_/S0 _7061_/A vssd1 vssd1 vccd1 vccd1
+ _4980_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_128_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ _4744_/B _3676_/A _4082_/B1 _6777_/A _3930_/X vssd1 vssd1 vccd1 vccd1 _3934_/B
+ sky130_fd_sc_hd__o221a_2
XFILLER_0_46_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3862_ _8087_/Q _3861_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__mux2_1
X_6650_ _7024_/A _6650_/A2 _6666_/A3 _6649_/X vssd1 vssd1 vccd1 vccd1 _6650_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5744__A1 _6175_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6581_ _6949_/A _6559_/B _6591_/B1 _6581_/B2 vssd1 vssd1 vccd1 vccd1 _6581_/X sky130_fd_sc_hd__a22o_1
X_5601_ _6939_/A _5616_/A2 _5616_/B1 hold457/X vssd1 vssd1 vccd1 vccd1 _5601_/X sky130_fd_sc_hd__a22o_1
X_5532_ _8251_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7721_/D sky130_fd_sc_hd__and3_1
X_3793_ _4763_/B _4071_/A2 _4071_/B1 _6947_/A _3792_/X vssd1 vssd1 vccd1 vccd1 _6191_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_42_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8320_ _8483_/CLK _8320_/D vssd1 vssd1 vccd1 vccd1 _8320_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8251_ _8251_/CLK _8251_/D vssd1 vssd1 vccd1 vccd1 _8251_/Q sky130_fd_sc_hd__dfxtp_1
X_5463_ _5463_/A _5465_/B _5463_/C vssd1 vssd1 vccd1 vccd1 _5463_/X sky130_fd_sc_hd__and3_1
XFILLER_0_100_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5394_ _6553_/A _6975_/C vssd1 vssd1 vccd1 vccd1 _5547_/B sky130_fd_sc_hd__nand2_1
X_8182_ _8402_/CLK _8182_/D vssd1 vssd1 vccd1 vccd1 _8182_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4414_ _4255_/Y _5454_/C _4413_/X _4412_/X vssd1 vssd1 vccd1 vccd1 _8372_/D sky130_fd_sc_hd__a31o_1
XFILLER_0_111_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4345_ _4335_/Y _4339_/B _4337_/B vssd1 vssd1 vccd1 vccd1 _4345_/X sky130_fd_sc_hd__o21a_1
Xfanout305 _5582_/Y vssd1 vssd1 vccd1 vccd1 _5616_/A2 sky130_fd_sc_hd__buf_8
XFILLER_0_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout316 _5186_/Y vssd1 vssd1 vccd1 vccd1 _5221_/A2 sky130_fd_sc_hd__buf_6
Xfanout338 _6815_/A vssd1 vssd1 vccd1 vccd1 _6947_/A sky130_fd_sc_hd__buf_4
Xfanout327 _3965_/X vssd1 vssd1 vccd1 vccd1 _6917_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6837__A _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout349 _6413_/B1 vssd1 vssd1 vccd1 vccd1 _6398_/B1 sky130_fd_sc_hd__buf_4
X_7064_ _7071_/B _7063_/Y _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8504_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__5460__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4276_ _4407_/A _4404_/B vssd1 vssd1 vccd1 vccd1 _4276_/Y sky130_fd_sc_hd__nand2_1
X_6015_ _6016_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout379_A _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout281_A _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7966_ _8030_/CLK _7966_/D vssd1 vssd1 vccd1 vccd1 _7966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_134_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7179__57 _8011_/CLK vssd1 vssd1 vccd1 vccd1 _8059_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__5188__A _6741_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7897_ _8504_/CLK _7897_/D vssd1 vssd1 vccd1 vccd1 _7897_/Q sky130_fd_sc_hd__dfxtp_1
X_6917_ _6917_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6917_/X sky130_fd_sc_hd__and2_1
X_6848_ _7010_/A _6848_/A2 _6845_/B _6847_/X vssd1 vssd1 vccd1 vccd1 _6848_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_119_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6779_ _6845_/A _6779_/B vssd1 vssd1 vccd1 vccd1 _6779_/Y sky130_fd_sc_hd__nor2_1
X_8518_ _8519_/CLK _8518_/D vssd1 vssd1 vccd1 vccd1 _8518_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5735__B2 _5789_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5830__S1 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8449_ _8485_/CLK _8449_/D vssd1 vssd1 vccd1 vccd1 _8449_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6160__A1 _6157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold370 _8208_/Q vssd1 vssd1 vccd1 vccd1 hold370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 _5427_/X vssd1 vssd1 vccd1 vccd1 _7616_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _7776_/Q vssd1 vssd1 vccd1 vccd1 hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5370__B _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1081 _8459_/Q vssd1 vssd1 vccd1 vccd1 _7001_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6215__A2 _6191_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1092 _6726_/X vssd1 vssd1 vccd1 vccd1 _8281_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1070 _7026_/X vssd1 vssd1 vccd1 vccd1 _8484_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6482__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4206__S _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5529__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7193__71 _8473_/CLK vssd1 vssd1 vccd1 vccd1 _8106_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5545__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6151__A1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4876__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5561__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4130_ _6206_/A _6209_/A _3896_/D _3892_/Y _6226_/A vssd1 vssd1 vccd1 vccd1 _4130_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__6657__A _6963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4061_ _6053_/A vssd1 vssd1 vccd1 vccd1 _4061_/Y sky130_fd_sc_hd__inv_2
X_7820_ _8346_/CLK _7820_/D vssd1 vssd1 vccd1 vccd1 _7820_/Q sky130_fd_sc_hd__dfxtp_1
X_7751_ _8370_/CLK _7751_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
X_4963_ _4962_/X _4961_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__mux2_1
X_3914_ _3914_/A _4081_/B vssd1 vssd1 vccd1 vccd1 _3914_/X sky130_fd_sc_hd__or2_1
X_7682_ _8451_/CLK _7682_/D vssd1 vssd1 vccd1 vccd1 _7682_/Q sky130_fd_sc_hd__dfxtp_1
X_6702_ _6971_/A _6669_/B _6702_/B1 hold841/X vssd1 vssd1 vccd1 vccd1 _6702_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3976__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5439__C _5470_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4894_ _4893_/X _4890_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8246_/D sky130_fd_sc_hd__mux2_1
X_6633_ _6939_/A _6665_/B vssd1 vssd1 vccd1 vccd1 _6633_/X sky130_fd_sc_hd__and2_1
XFILLER_0_117_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3845_ _4118_/A _6126_/A vssd1 vssd1 vccd1 vccd1 _3846_/B sky130_fd_sc_hd__or2_1
XFILLER_0_27_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6564_ _6849_/A _6560_/B _6560_/Y hold280/X vssd1 vssd1 vccd1 vccd1 _6564_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_104_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3776_ _6157_/A _6154_/A vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8303_ _8465_/CLK _8303_/D vssd1 vssd1 vccd1 vccd1 _8303_/Q sky130_fd_sc_hd__dfxtp_1
X_6495_ _6498_/A hold3/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__and2_1
XANTENNA__5455__B _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5515_ _8234_/Q _5538_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _7704_/D sky130_fd_sc_hd__and3_1
X_5446_ _5446_/A _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8234_ _8234_/CLK _8234_/D vssd1 vssd1 vccd1 vccd1 _8234_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5471__A _7052_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5377_ _5408_/C _5388_/C vssd1 vssd1 vccd1 vccd1 _6553_/B sky130_fd_sc_hd__nor2_1
X_8165_ _8515_/CLK _8165_/D vssd1 vssd1 vccd1 vccd1 _8165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6693__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4328_ _8492_/Q _4329_/B vssd1 vssd1 vccd1 vccd1 _4328_/Y sky130_fd_sc_hd__nor2_1
X_8096_ _8096_/CLK _8130_/D vssd1 vssd1 vccd1 vccd1 _8096_/Q sky130_fd_sc_hd__dfxtp_1
X_7116_ _7273_/A vssd1 vssd1 vccd1 vccd1 _7116_/Y sky130_fd_sc_hd__inv_2
Xfanout179 hold1510/X vssd1 vssd1 vccd1 vccd1 _7073_/A sky130_fd_sc_hd__buf_6
Xfanout168 hold1510/X vssd1 vssd1 vccd1 vccd1 _5541_/B sky130_fd_sc_hd__clkbuf_4
X_7047_ _7031_/Y _7046_/Y _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8496_/D sky130_fd_sc_hd__a21oi_1
X_4259_ _4249_/Y _4253_/B _4250_/Y vssd1 vssd1 vccd1 vccd1 _4260_/B sky130_fd_sc_hd__o21a_1
XANTENNA__5653__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4551__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7949_ _8510_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 _7949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__B1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1680_A _3795_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5708__A1 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3719__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6381__A1 _6412_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6133__A1 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6684__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5381__A _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6477__A _6550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4790__S1 _4867_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5644__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4542__S1 _4640_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7101__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5556__A _6494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4460__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5300_ _6706_/A _5300_/B vssd1 vssd1 vccd1 vccd1 _5300_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_59_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6280_ _6281_/A _6281_/B vssd1 vssd1 vccd1 vccd1 _6280_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5231_ _6849_/A _5227_/B _5227_/Y hold254/X vssd1 vssd1 vccd1 vccd1 _5231_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6387__A _6388_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6675__A2 _6701_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5883__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5162_ _5162_/A1 _5067_/S _5172_/B1 _5161_/X vssd1 vssd1 vccd1 vccd1 _7393_/D sky130_fd_sc_hd__o211a_1
X_5093_ _5477_/A _5546_/C vssd1 vssd1 vccd1 vccd1 _5093_/X sky130_fd_sc_hd__or2_1
Xhold1806 _7372_/Q vssd1 vssd1 vccd1 vccd1 hold1806/X sky130_fd_sc_hd__dlygate4sd3_1
X_4113_ _4061_/Y _6056_/A _4090_/D _4086_/Y _6075_/A vssd1 vssd1 vccd1 vccd1 _4113_/X
+ sky130_fd_sc_hd__o32a_1
Xhold1817 _7888_/Q vssd1 vssd1 vccd1 vccd1 hold1817/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5635__B1 _5653_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4044_ _4044_/A _4044_/B vssd1 vssd1 vccd1 vccd1 _4045_/D sky130_fd_sc_hd__and2_1
XFILLER_0_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7803_ _8326_/CLK _7803_/D vssd1 vssd1 vccd1 vccd1 _7803_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__7011__A _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7734_ _8456_/CLK _7734_/D vssd1 vssd1 vccd1 vccd1 _7734_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _5976_/A _5975_/A _5973_/Y vssd1 vssd1 vccd1 vccd1 _5996_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_91_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout244_A _3676_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7149__27 _8353_/CLK vssd1 vssd1 vccd1 vccd1 _7526_/CLK sky130_fd_sc_hd__inv_2
X_4946_ _4944_/X _4945_/X _7059_/A vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__mux2_1
X_7665_ _8456_/CLK _7665_/D vssd1 vssd1 vccd1 vccd1 _7665_/Q sky130_fd_sc_hd__dfxtp_1
X_4877_ _8180_/Q _8212_/Q _8276_/Q _7784_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4877_/X sky130_fd_sc_hd__mux4_1
X_6616_ _7008_/A _6616_/A2 _6605_/B _6615_/X vssd1 vssd1 vccd1 vccd1 _6616_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_105_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7596_ _8515_/CLK _7596_/D vssd1 vssd1 vccd1 vccd1 _7596_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout411_A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3828_ _4773_/B _4071_/A2 _4071_/B1 _6967_/A _3827_/X vssd1 vssd1 vccd1 vccd1 _6370_/A
+ sky130_fd_sc_hd__o221a_4
XANTENNA__5166__A2 _4416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6547_ _7008_/A _6547_/B vssd1 vssd1 vccd1 vccd1 _8029_/D sky130_fd_sc_hd__and2_1
XFILLER_0_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__6902__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3759_ _3759_/A _3759_/B vssd1 vssd1 vccd1 vccd1 _6137_/A sky130_fd_sc_hd__nand2_2
X_6478_ _7005_/A _6478_/B vssd1 vssd1 vccd1 vccd1 _6478_/X sky130_fd_sc_hd__and2_1
XFILLER_0_100_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8217_ _8475_/CLK _8217_/D vssd1 vssd1 vccd1 vccd1 _8217_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6297__A _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5429_ _5429_/A _5465_/B _5465_/C vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__and3_1
X_8148_ _8450_/CLK _8148_/D vssd1 vssd1 vccd1 vccd1 _8148_/Q sky130_fd_sc_hd__dfxtp_1
X_8079_ _8079_/CLK _8113_/D vssd1 vssd1 vccd1 vccd1 _8079_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5626__B1 _5652_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__S1 _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5376__A _5408_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7163__41 _8283_/CLK vssd1 vssd1 vccd1 vccd1 _8043_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6919__B _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5542__C _5542_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6409__A2 _6126_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5617__B1 _5617_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4455__A _7024_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6268__S1 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4800_ _8169_/Q _8201_/Q _8265_/Q _7773_/Q _4895_/S0 _4867_/S1 vssd1 vssd1 vccd1
+ vccd1 _4800_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6670__A _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5780_ _6016_/A _5993_/A _6056_/A _6035_/A _5772_/S _5797_/S vssd1 vssd1 vccd1 vccd1
+ _5780_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_84_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4731_ _8163_/Q _7562_/Q _7434_/Q _7594_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4731_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5148__A2 _4425_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7450_ _8154_/CLK _7450_/D vssd1 vssd1 vccd1 vccd1 _7450_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4662_ _4660_/X _4661_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5699__A3 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6401_ _6391_/Y _6396_/X _6397_/Y _6399_/X _6400_/Y vssd1 vssd1 vccd1 vccd1 _7898_/D
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_3_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4593_ _8176_/Q _8208_/Q _8272_/Q _7780_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4593_/X sky130_fd_sc_hd__mux4_1
X_7381_ _8370_/CLK _7381_/D vssd1 vssd1 vccd1 vccd1 _7381_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 _8486_/Q vssd1 vssd1 vccd1 vccd1 _7028_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 _7023_/X vssd1 vssd1 vccd1 vccd1 _8481_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6332_ _6334_/A _6334_/B vssd1 vssd1 vccd1 vccd1 _6335_/A sky130_fd_sc_hd__and2_1
Xhold925 _8205_/Q vssd1 vssd1 vccd1 vccd1 hold925/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6829__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold914 _7016_/X vssd1 vssd1 vccd1 vccd1 _8474_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 _5320_/X vssd1 vssd1 vccd1 vccd1 _7551_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6263_ _6263_/A _6263_/B vssd1 vssd1 vccd1 vccd1 _6266_/A sky130_fd_sc_hd__nor2_1
Xhold947 _7800_/Q vssd1 vssd1 vccd1 vccd1 hold947/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold969 _8282_/Q vssd1 vssd1 vccd1 vccd1 hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7006__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8002_ _8515_/CLK hold82/X vssd1 vssd1 vccd1 vccd1 _8002_/Q sky130_fd_sc_hd__dfxtp_1
X_5214_ _6891_/A _5188_/B _5220_/B1 hold603/X vssd1 vssd1 vccd1 vccd1 _5214_/X sky130_fd_sc_hd__a22o_1
X_6194_ _6194_/A _6194_/B vssd1 vssd1 vccd1 vccd1 _6194_/X sky130_fd_sc_hd__xor2_1
XANTENNA__5320__A2 _5299_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5145_ _5452_/A _5453_/C vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__or2_1
Xhold1614 _4190_/X vssd1 vssd1 vccd1 vccd1 _5556_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1603 _4174_/Y vssd1 vssd1 vccd1 vccd1 _4176_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5608__B1 _5616_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1625 _4295_/X vssd1 vssd1 vccd1 vccd1 _5571_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5076_ input29/X _5099_/B _5148_/B1 _5075_/X vssd1 vssd1 vccd1 vccd1 _7350_/D sky130_fd_sc_hd__o211a_1
Xhold1669 _7680_/Q vssd1 vssd1 vccd1 vccd1 _4059_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1636 _4084_/X vssd1 vssd1 vccd1 vccd1 _6434_/B sky130_fd_sc_hd__buf_1
Xhold1647 _4352_/X vssd1 vssd1 vccd1 vccd1 _5579_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1658 _3816_/X vssd1 vssd1 vccd1 vccd1 _6449_/B sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__4365__A _5476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4027_ _4755_/B _4072_/B vssd1 vssd1 vccd1 vccd1 _4027_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout459_A _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5978_ _6008_/A _5694_/Y _5718_/X _5955_/Y _5881_/C vssd1 vssd1 vccd1 vccd1 _5978_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6584__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7717_ _8473_/CLK _7717_/D vssd1 vssd1 vccd1 vccd1 _7717_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5380__A_N _7065_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4929_ _4928_/X _4925_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8251_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1476_A _7293_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4304__S _5503_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7648_ _8378_/CLK _7648_/D vssd1 vssd1 vccd1 vccd1 _7648_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7579_ _8431_/CLK _7579_/D vssd1 vssd1 vccd1 vccd1 _7579_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4993__S1 _4997_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6195__S0 _5782_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5311__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4974__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6272__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6024__A0 _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6490__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6575__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5818__B _6094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4050__A2 _3676_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__S0 _4734_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5537__C _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6327__B2 _6130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output88_A _8132_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6649__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5302__A2 _5332_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6665__A _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3864__A2 _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6950_ _7018_/A _6950_/A2 _6970_/A3 _6949_/X vssd1 vssd1 vccd1 vccd1 _6950_/X sky130_fd_sc_hd__a31o_1
X_5901_ _5952_/A _5753_/Y _5836_/B vssd1 vssd1 vccd1 vccd1 _5901_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_80_clk_A clkbuf_4_7_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6881_ _6947_/A _6905_/B vssd1 vssd1 vccd1 vccd1 _6881_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6566__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5832_ _5830_/X _5831_/X _5950_/S vssd1 vssd1 vccd1 vccd1 _5832_/X sky130_fd_sc_hd__mux2_1
X_5763_ _5763_/A _5763_/B _5971_/B vssd1 vssd1 vccd1 vccd1 _5765_/B sky130_fd_sc_hd__or3_1
XANTENNA__5728__B _6380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7502_ _7502_/CLK _7502_/D vssd1 vssd1 vccd1 vccd1 _7502_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4714_ _4713_/X _4712_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4714_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_95_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5447__C _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5694_ _6128_/A _6129_/B vssd1 vssd1 vccd1 vccd1 _5694_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_71_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8482_ _8483_/CLK _8482_/D vssd1 vssd1 vccd1 vccd1 _8482_/Q sky130_fd_sc_hd__dfxtp_1
X_4645_ _4644_/X _4641_/X _5474_/A vssd1 vssd1 vccd1 vccd1 _7517_/D sky130_fd_sc_hd__mux2_1
X_7433_ _8427_/CLK _7433_/D vssd1 vssd1 vccd1 vccd1 _7433_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4576_ _8334_/Q _7810_/Q _7476_/Q _7444_/Q _7072_/B2 _5472_/A vssd1 vssd1 vccd1 vccd1
+ _4576_/X sky130_fd_sc_hd__mux4_1
Xhold711 _7595_/Q vssd1 vssd1 vccd1 vccd1 hold711/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold700 _5356_/X vssd1 vssd1 vccd1 vccd1 _7583_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7364_ _8476_/CLK _7364_/D vssd1 vssd1 vccd1 vccd1 _7364_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold733 _8303_/Q vssd1 vssd1 vccd1 vccd1 hold733/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6559__B _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold744 _7012_/X vssd1 vssd1 vccd1 vccd1 _8470_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4975__S1 _4976_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6315_ _6315_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6318_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold755 _8292_/Q vssd1 vssd1 vccd1 vccd1 hold755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold722 _7002_/X vssd1 vssd1 vccd1 vccd1 _8460_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5463__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold788 _5270_/X vssd1 vssd1 vccd1 vccd1 _7474_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7295_ _8370_/CLK _7295_/D _7105_/Y vssd1 vssd1 vccd1 vccd1 _7295_/Q sky130_fd_sc_hd__dfrtp_4
Xhold777 _7557_/Q vssd1 vssd1 vccd1 vccd1 hold777/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold766 _5597_/X vssd1 vssd1 vccd1 vccd1 _7781_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold799 _8322_/Q vssd1 vssd1 vccd1 vccd1 hold799/X sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ _6246_/A _6246_/B vssd1 vssd1 vccd1 vccd1 _6247_/B sky130_fd_sc_hd__nand2_1
XANTENNA__4727__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1400 _4422_/A vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__buf_1
X_6177_ _6177_/A _6177_/B vssd1 vssd1 vccd1 vccd1 _6177_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5128_ _5128_/A1 _5182_/A2 _5182_/B1 _5127_/X vssd1 vssd1 vccd1 vccd1 _7376_/D sky130_fd_sc_hd__o211a_1
Xhold1422 _4357_/Y vssd1 vssd1 vccd1 vccd1 _5580_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3855__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1433 _8379_/Q vssd1 vssd1 vccd1 vccd1 _5046_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 hold1801/X vssd1 vssd1 vccd1 vccd1 _4768_/B sky130_fd_sc_hd__clkbuf_2
Xhold1466 hold1808/X vssd1 vssd1 vccd1 vccd1 _4755_/B sky130_fd_sc_hd__buf_1
Xhold1444 _7032_/Y vssd1 vssd1 vccd1 vccd1 _7033_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6254__B1 _6398_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1477 _7307_/Q vssd1 vssd1 vccd1 vccd1 _5170_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 _7643_/Q vssd1 vssd1 vccd1 vccd1 _4243_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_48_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1499 hold1813/X vssd1 vssd1 vccd1 vccd1 _4760_/B sky130_fd_sc_hd__buf_1
X_5059_ _5439_/A _5470_/C vssd1 vssd1 vccd1 vccd1 _5059_/X sky130_fd_sc_hd__or2_1
Xhold1488 _7311_/Q vssd1 vssd1 vccd1 vccd1 _5178_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5919__A _5921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4663__S0 _4706_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5780__A2 _6056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_106_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3791__A1 _3790_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5654__A _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7133__11 _8332_/CLK vssd1 vssd1 vccd1 vccd1 _7510_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_133_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4966__S1 _4969_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6485__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6796__A1 _7007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5599__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6340__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4023__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4654__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4452__B _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5220__A1 _6969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_14_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_14_0_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4879__S _4998_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _4430_/A _4430_/B vssd1 vssd1 vccd1 vccd1 _4430_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_2 _7885_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4361_ _7052_/A _7732_/Q _7734_/Q _3648_/Y _4360_/X vssd1 vssd1 vccd1 vccd1 _4361_/X
+ sky130_fd_sc_hd__a221o_1
X_6100_ _6024_/X _6099_/X _6393_/A vssd1 vssd1 vccd1 vccd1 _6100_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_7080_ _5389_/X _5402_/B _7055_/A vssd1 vssd1 vccd1 vccd1 _7080_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_67_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5287__A1 _6955_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4709__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4292_ _8497_/Q _4292_/B vssd1 vssd1 vccd1 vccd1 _4292_/Y sky130_fd_sc_hd__nand2_1
X_6031_ _4008_/B _6063_/A _6023_/Y _6031_/B2 _6911_/A vssd1 vssd1 vccd1 vccd1 _6031_/Y
+ sky130_fd_sc_hd__a221oi_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3837__A2 _8034_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7982_ _8079_/CLK _7982_/D vssd1 vssd1 vccd1 vccd1 _7982_/Q sky130_fd_sc_hd__dfxtp_1
X_6933_ _6933_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6933_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6864_ _7008_/A _6864_/A2 _6842_/X _6863_/X vssd1 vssd1 vccd1 vccd1 _6864_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5739__A _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5815_ _6128_/A _5815_/B _5815_/C vssd1 vssd1 vccd1 vccd1 _5815_/X sky130_fd_sc_hd__or3_1
XANTENNA__5458__B _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5211__A1 _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6795_ _6927_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6795_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5746_ _6281_/A _6244_/A _6262_/A _6226_/A _5860_/S _3928_/X vssd1 vssd1 vccd1 vccd1
+ _5746_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_45_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4789__S _4929_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8465_ _8465_/CLK _8465_/D vssd1 vssd1 vccd1 vccd1 _8465_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5677_ _7027_/A hold17/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__and2_1
XANTENNA__5474__A _5474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7416_ _8143_/CLK _7416_/D vssd1 vssd1 vccd1 vccd1 _7416_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4628_ _8181_/Q _8213_/Q _8277_/Q _7785_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4628_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_130_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold530 _6674_/X vssd1 vssd1 vccd1 vccd1 _8201_/D sky130_fd_sc_hd__dlygate4sd3_1
X_8396_ _8464_/CLK _8396_/D vssd1 vssd1 vccd1 vccd1 _8396_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6711__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4948__S1 _7061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold552 _6716_/X vssd1 vssd1 vccd1 vccd1 _8271_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 _7473_/Q vssd1 vssd1 vccd1 vccd1 hold541/X sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _8461_/Q _8393_/Q _8425_/Q _8299_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4559_/X sky130_fd_sc_hd__mux4_1
X_7347_ _8501_/CLK _7347_/D vssd1 vssd1 vccd1 vccd1 _7347_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold563 _7494_/Q vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold596 _5240_/X vssd1 vssd1 vccd1 vccd1 _7448_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _8302_/Q vssd1 vssd1 vccd1 vccd1 hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _6680_/X vssd1 vssd1 vccd1 vccd1 _8207_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold1439_A _7289_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5278__A1 _6937_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7278_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7278_/Y sky130_fd_sc_hd__inv_2
X_6229_ _6229_/A _6229_/B vssd1 vssd1 vccd1 vccd1 _6229_/X sky130_fd_sc_hd__xor2_1
XANTENNA__3828__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1241 _8438_/Q vssd1 vssd1 vccd1 vccd1 _6946_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 _6644_/X vssd1 vssd1 vccd1 vccd1 _8186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1230 _6940_/X vssd1 vssd1 vccd1 vccd1 _8435_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6778__A1 _6706_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4029__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6322__S0 _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1285 _6960_/X vssd1 vssd1 vccd1 vccd1 _8445_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _7038_/Y vssd1 vssd1 vccd1 vccd1 _7039_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1263 _8195_/Q vssd1 vssd1 vccd1 vccd1 _6662_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1296 _8192_/Q vssd1 vssd1 vccd1 vccd1 _6656_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4884__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4516__A_N _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4636__S0 _3649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5753__A2 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6950__A1 _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6702__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput94 _8109_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[8] sky130_fd_sc_hd__buf_12
XANTENNA__6927__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5269__A1 _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput72 _8118_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[17] sky130_fd_sc_hd__buf_12
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput83 _8128_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[27] sky130_fd_sc_hd__buf_12
XFILLER_0_128_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7104__A _7264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4046__A_N _3923_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6769__A1 _6961_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6233__A3 _6226_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3930_ _7700_/Q _4081_/B vssd1 vssd1 vccd1 vccd1 _3930_/X sky130_fd_sc_hd__or2_1
XANTENNA__5559__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4875__S0 _4997_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4463__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3861_ _7991_/Q _4068_/A2 _4068_/B1 _8023_/Q _3860_/X vssd1 vssd1 vccd1 vccd1 _3861_/X
+ sky130_fd_sc_hd__a221o_2
X_5600_ _6937_/A _5584_/B _5617_/B1 hold655/X vssd1 vssd1 vccd1 vccd1 _5600_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_73_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6580_ _6947_/A _6559_/B _6591_/B1 _6580_/B2 vssd1 vssd1 vccd1 vccd1 _6580_/X sky130_fd_sc_hd__a22o_1
X_3792_ _7719_/Q _4070_/B vssd1 vssd1 vccd1 vccd1 _3792_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5531_ _8250_/Q _5538_/B _5538_/C vssd1 vssd1 vccd1 vccd1 _7720_/D sky130_fd_sc_hd__and3_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8250_ _8250_/CLK _8250_/D vssd1 vssd1 vccd1 vccd1 _8250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_112_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5462_ _5462_/A _5503_/B _5462_/C vssd1 vssd1 vccd1 vccd1 _5462_/X sky130_fd_sc_hd__and3_1
X_5393_ _6553_/A _6975_/C vssd1 vssd1 vccd1 vccd1 _7071_/A sky130_fd_sc_hd__and2_1
XFILLER_0_50_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8181_ _8431_/CLK _8181_/D vssd1 vssd1 vccd1 vccd1 _8181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4413_ _4416_/A _4413_/B vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__or2_1
X_4344_ _4342_/Y _4344_/B vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout328 _3954_/X vssd1 vssd1 vccd1 vccd1 _6921_/A sky130_fd_sc_hd__buf_4
Xfanout306 _5582_/Y vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__buf_6
Xfanout317 _4080_/X vssd1 vssd1 vccd1 vccd1 _6935_/A sky130_fd_sc_hd__buf_4
X_7063_ _7063_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7063_/Y sky130_fd_sc_hd__nand2_1
Xfanout339 _3779_/X vssd1 vssd1 vccd1 vccd1 _6945_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6837__B _6837_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6014_ _6016_/A _6016_/B vssd1 vssd1 vccd1 vccd1 _6017_/A sky130_fd_sc_hd__nand2_1
XANTENNA__7014__A _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4275_ _4274_/X _4403_/A _5540_/B vssd1 vssd1 vccd1 vccd1 _4404_/B sky130_fd_sc_hd__mux2_1
XANTENNA__6853__A _6853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout274_A _3669_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7965_ _8096_/CLK hold34/X vssd1 vssd1 vccd1 vccd1 _7965_/Q sky130_fd_sc_hd__dfxtp_1
X_6916_ _7010_/A _6916_/A2 _6943_/B _6915_/X vssd1 vssd1 vccd1 vccd1 _6916_/X sky130_fd_sc_hd__a31o_1
X_7896_ _8500_/CLK _7896_/D vssd1 vssd1 vccd1 vccd1 _7896_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout441_A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6847_ _6847_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6847_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5188__B _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5196__B1 _5221_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6778_ _6706_/A _6778_/A2 _6779_/B _6777_/X vssd1 vssd1 vccd1 vccd1 _6778_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_119_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5735__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4618__S0 _4696_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6932__A1 _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8517_ _8517_/CLK _8517_/D vssd1 vssd1 vccd1 vccd1 _8517_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5729_ _5730_/A _5730_/B vssd1 vssd1 vccd1 vccd1 _5738_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3746__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold1556_A _3917_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8448_ _8448_/CLK _8448_/D vssd1 vssd1 vccd1 vccd1 _8448_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_111_clk clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _8353_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_102_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6696__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8379_ _8379_/CLK _8379_/D _7273_/Y vssd1 vssd1 vccd1 vccd1 _8379_/Q sky130_fd_sc_hd__dfrtp_1
Xhold371 _6681_/X vssd1 vssd1 vccd1 vccd1 _8208_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _7535_/Q vssd1 vssd1 vccd1 vccd1 hold360/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold393 _5592_/X vssd1 vssd1 vccd1 vccd1 _7776_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _7383_/Q vssd1 vssd1 vccd1 vccd1 _5450_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5120__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1060 _6772_/X vssd1 vssd1 vccd1 vccd1 _8323_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1082 _7001_/X vssd1 vssd1 vccd1 vccd1 _8459_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 _8465_/Q vssd1 vssd1 vccd1 vccd1 _7007_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6215__A3 _6209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1093 _7475_/Q vssd1 vssd1 vccd1 vccd1 _5271_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3682__B1 _4068_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5959__C1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4857__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5545__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_102_clk clkbuf_4_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _8427_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6687__B1 _6702_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output70_A _8116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6657__B _6661_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4458__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4060_ _4221_/A _4059_/X _4085_/S vssd1 vssd1 vccd1 vccd1 _6053_/A sky130_fd_sc_hd__mux2_2
X_7750_ _8368_/CLK _7750_/D vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _8482_/Q _8414_/Q _8446_/Q _8320_/Q _4990_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4962_/X sky130_fd_sc_hd__mux4_1
X_3913_ _8069_/Q _3912_/X _4080_/S vssd1 vssd1 vccd1 vccd1 _6913_/A sky130_fd_sc_hd__mux2_2
X_7681_ _8328_/CLK _7681_/D vssd1 vssd1 vccd1 vccd1 _7681_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3976__B2 _8010_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4893_ _4892_/X _4891_/X _4991_/S vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__mux2_1
X_6701_ _6969_/A _6701_/A2 _6701_/B1 _6701_/B2 vssd1 vssd1 vccd1 vccd1 _6701_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_104_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6632_ _7019_/A _6632_/A2 _6605_/B _6631_/X vssd1 vssd1 vccd1 vccd1 _6632_/X sky130_fd_sc_hd__a31o_1
X_3844_ _4118_/A _6126_/A vssd1 vssd1 vccd1 vccd1 _3846_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5178__B1 _5182_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6914__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6563_ _6847_/A _6560_/B _6560_/Y hold304/X vssd1 vssd1 vccd1 vccd1 _6563_/X sky130_fd_sc_hd__o22a_1
X_3775_ _6157_/A _6154_/A vssd1 vssd1 vccd1 vccd1 _3775_/X sky130_fd_sc_hd__or2_1
XANTENNA__7009__A _7023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_8302_ _8428_/CLK _8302_/D vssd1 vssd1 vccd1 vccd1 _8302_/Q sky130_fd_sc_hd__dfxtp_1
X_5514_ _8233_/Q _5528_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7703_/D sky130_fd_sc_hd__and3_1
X_6494_ _6494_/A hold71/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__and2_1
XFILLER_0_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_8233_ _8233_/CLK _8233_/D vssd1 vssd1 vccd1 vccd1 _8233_/Q sky130_fd_sc_hd__dfxtp_1
X_5445_ _5445_/A _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5445_/X sky130_fd_sc_hd__and3_1
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6678__B1 _6701_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5350__B1 _5368_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8164_ _8487_/CLK _8164_/D vssd1 vssd1 vccd1 vccd1 _8164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5752__A _5804_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5471__B _7090_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5376_ _5408_/B _5391_/A vssd1 vssd1 vccd1 vccd1 _5388_/C sky130_fd_sc_hd__nand2_1
XANTENNA__3900__A1 _3899_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7115_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7115_/Y sky130_fd_sc_hd__inv_2
X_8095_ _8500_/CLK _8129_/D vssd1 vssd1 vccd1 vccd1 _8095_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout391_A _7362_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4327_ _4390_/A _4390_/B _4327_/C _4385_/B vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__and4_2
XANTENNA__5102__B1 _5148_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7046_ _7046_/A _7046_/B vssd1 vssd1 vccd1 vccd1 _7046_/Y sky130_fd_sc_hd__nand2_1
Xfanout169 _7030_/B vssd1 vssd1 vccd1 vccd1 _5503_/B sky130_fd_sc_hd__buf_4
X_4258_ _4256_/Y _4258_/B vssd1 vssd1 vccd1 vccd1 _4258_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__5653__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4189_ _4183_/A _4180_/Y _4182_/B vssd1 vssd1 vccd1 vccd1 _4189_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4839__S0 _4895_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7948_ _8365_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 _7948_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3967__B2 _4073_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7879_ _8086_/CLK _7879_/D vssd1 vssd1 vccd1 vccd1 _7879_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3719__A1 _4770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3719__B2 _3717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4977__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5662__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5341__B1 _5367_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold190 _7599_/Q vssd1 vssd1 vccd1 vccd1 _6420_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4447__A2 _7030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6493__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5644__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3958__B2 _4084_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4887__S _4999_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5230_ _6847_/A _5226_/B _5259_/B1 hold775/X vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6124__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3791__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5572__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5332__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8529__470 vssd1 vssd1 vccd1 vccd1 _8529__470/HI _8529_/A sky130_fd_sc_hd__conb_1
XANTENNA__5883__B2 _6251_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3804__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5161_ hold43/X _5463_/C vssd1 vssd1 vccd1 vccd1 _5161_/X sky130_fd_sc_hd__or2_1
Xhold1807 _7878_/Q vssd1 vssd1 vccd1 vccd1 hold1807/X sky130_fd_sc_hd__dlygate4sd3_1
X_4112_ _6096_/A _6094_/A vssd1 vssd1 vccd1 vccd1 _4112_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1818 _7896_/Q vssd1 vssd1 vccd1 vccd1 hold1818/X sky130_fd_sc_hd__dlygate4sd3_1
X_5092_ input7/X _5067_/S _5172_/B1 _5091_/X vssd1 vssd1 vccd1 vccd1 _7358_/D sky130_fd_sc_hd__o211a_1
X_4043_ _5993_/A _5990_/A vssd1 vssd1 vccd1 vccd1 _4044_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7802_ _7805_/CLK _7802_/D vssd1 vssd1 vccd1 vccd1 _7802_/Q sky130_fd_sc_hd__dfxtp_1
X_5994_ _5994_/A _5994_/B vssd1 vssd1 vccd1 vccd1 _5996_/A sky130_fd_sc_hd__nor2_1
X_7733_ _8456_/CLK _7733_/D vssd1 vssd1 vccd1 vccd1 _7733_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4945_ _8157_/Q _7556_/Q _7428_/Q _7588_/Q _4983_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4945_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4071__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7664_ _8456_/CLK _7664_/D vssd1 vssd1 vccd1 vccd1 _7664_/Q sky130_fd_sc_hd__dfxtp_1
X_4876_ _4874_/X _4875_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout237_A _5099_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6615_ _6921_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6615_/X sky130_fd_sc_hd__and2_1
X_7595_ _8487_/CLK _7595_/D vssd1 vssd1 vccd1 vccd1 _7595_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6363__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5466__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3827_ _3827_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3827_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout404_A hold1746/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6546_ _6706_/A _6546_/B vssd1 vssd1 vccd1 vccd1 _8028_/D sky130_fd_sc_hd__and2_1
XFILLER_0_131_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3758_ _3968_/A _4250_/A vssd1 vssd1 vccd1 vccd1 _3759_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3689_ _7836_/Q _7662_/Q vssd1 vssd1 vccd1 vccd1 _3689_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_113_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6477_ _6550_/A hold92/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__and2_1
XANTENNA__6666__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5323__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_8216_ _8346_/CLK _8216_/D vssd1 vssd1 vccd1 vccd1 _8216_/Q sky130_fd_sc_hd__dfxtp_1
X_5428_ _5428_/A _5540_/B _5456_/C vssd1 vssd1 vccd1 vccd1 _5428_/X sky130_fd_sc_hd__and3_1
XFILLER_0_100_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8147_ _8469_/CLK _8147_/D vssd1 vssd1 vccd1 vccd1 _8147_/Q sky130_fd_sc_hd__dfxtp_1
X_5359_ _6953_/A _5367_/A2 _5367_/B1 hold945/X vssd1 vssd1 vccd1 vccd1 _5359_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3885__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8078_ _8086_/CLK _8112_/D vssd1 vssd1 vccd1 vccd1 _8078_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4429__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7029_ _7029_/A _7029_/B vssd1 vssd1 vccd1 vccd1 _7029_/X sky130_fd_sc_hd__and2_1
XANTENNA__5626__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5657__A _5667_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5376__B _5391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5392__A _7346_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6106__A2 _5732_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3905__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6488__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5314__B1 _5332_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6409__A3 _6370_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6935__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5617__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7112__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6290__A1 _6270_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6951__A _6951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__A0 _8505_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5567__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _8356_/Q _7832_/Q _7498_/Q _7466_/Q _3649_/A _4731_/S1 vssd1 vssd1 vccd1 vccd1
+ _4730_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4471__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6345__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4661_ _8153_/Q _7552_/Q _7424_/Q _7584_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4661_/X sky130_fd_sc_hd__mux4_1
X_7380_ _7977_/CLK _7380_/D vssd1 vssd1 vccd1 vccd1 _7380_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_71_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6400_ _6400_/A1 _6292_/A _7279_/A vssd1 vssd1 vccd1 vccd1 _6400_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4592_ _4590_/X _4591_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4592_/X sky130_fd_sc_hd__mux2_1
X_6331_ _6331_/A _6405_/B vssd1 vssd1 vccd1 vccd1 _6334_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6896__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold904 _7028_/X vssd1 vssd1 vccd1 vccd1 _8486_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _8145_/Q vssd1 vssd1 vccd1 vccd1 hold937/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 _7545_/Q vssd1 vssd1 vccd1 vccd1 hold915/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3815__A _4772_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold926 _6678_/X vssd1 vssd1 vccd1 vccd1 _8205_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold959 _7571_/Q vssd1 vssd1 vccd1 vccd1 hold959/X sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ _6262_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6263_/B sky130_fd_sc_hd__nor2_1
Xhold948 _5616_/X vssd1 vssd1 vccd1 vccd1 _7800_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6648__A3 _6666_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5305__B1 _5331_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5856__A1 _5870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_8001_ _8030_/CLK _8001_/D vssd1 vssd1 vccd1 vccd1 _8001_/Q sky130_fd_sc_hd__dfxtp_1
X_6193_ _6177_/A _6176_/A _6174_/Y vssd1 vssd1 vccd1 vccd1 _6194_/B sky130_fd_sc_hd__a21o_1
X_5213_ _6955_/A _5188_/B _5220_/B1 hold609/X vssd1 vssd1 vccd1 vccd1 _5213_/X sky130_fd_sc_hd__a22o_1
X_5144_ _5144_/A1 _5144_/A2 _5146_/B1 _5143_/X vssd1 vssd1 vccd1 vccd1 _7384_/D sky130_fd_sc_hd__o211a_1
XANTENNA__7058__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6845__B _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1626 _7637_/Q vssd1 vssd1 vccd1 vccd1 _4202_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1615 _4192_/A vssd1 vssd1 vccd1 vccd1 _4509_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1604 _4176_/X vssd1 vssd1 vccd1 vccd1 _5554_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5608__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5075_ _5544_/A _5523_/C vssd1 vssd1 vccd1 vccd1 _5075_/X sky130_fd_sc_hd__or2_1
Xhold1648 hold1818/X vssd1 vssd1 vccd1 vccd1 _4772_/B sky130_fd_sc_hd__clkbuf_2
Xhold1659 _7360_/Q vssd1 vssd1 vccd1 vccd1 hold1659/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1637 _7364_/Q vssd1 vssd1 vccd1 vccd1 hold1637/X sky130_fd_sc_hd__buf_2
XANTENNA__5084__A2 _5144_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7209__87 _8451_/CLK vssd1 vssd1 vccd1 vccd1 _8122_/CLK sky130_fd_sc_hd__inv_2
XANTENNA__6820__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4026_ _4755_/B _4071_/A2 _4071_/B1 _4024_/X _4025_/X vssd1 vssd1 vccd1 vccd1 _6035_/A
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6861__A _6927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_91_clk clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 _8379_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5477__A _5477_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5977_ _5976_/A _5976_/B _6030_/A1 vssd1 vssd1 vccd1 vccd1 _5977_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6584__A2 _6559_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4928_ _4927_/X _4926_/X _4998_/S vssd1 vssd1 vccd1 vccd1 _4928_/X sky130_fd_sc_hd__mux2_1
X_7716_ _8319_/CLK _7716_/D vssd1 vssd1 vccd1 vccd1 _7716_/Q sky130_fd_sc_hd__dfxtp_1
X_7647_ _8071_/CLK _7647_/D vssd1 vssd1 vccd1 vccd1 _7647_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold1469_A _7292_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4859_ _4858_/X _4855_/X _4999_/S vssd1 vssd1 vccd1 vccd1 _8241_/D sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_7_clk_A clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7578_ _8154_/CLK _7578_/D vssd1 vssd1 vccd1 vccd1 _7578_/Q sky130_fd_sc_hd__dfxtp_1
X_6529_ _6552_/A _6529_/B vssd1 vssd1 vccd1 vccd1 _8011_/D sky130_fd_sc_hd__and2_1
XANTENNA_hold1636_A _4084_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6195__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7049__B1 _7064_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6024__A1 _5974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_82_clk clkbuf_4_6_0_clk/X vssd1 vssd1 vccd1 vccd1 _8071_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_128_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6575__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4681__S1 _4734_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6327__A2 _6414_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6878__A3 _6845_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__7107__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6665__B _6665_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4466__A _6999_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6802__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5066__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5900_ _6129_/B _5900_/B _5900_/C vssd1 vssd1 vccd1 vccd1 _5900_/X sky130_fd_sc_hd__or3_1
XFILLER_0_49_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_73_clk clkbuf_4_12_0_clk/X vssd1 vssd1 vccd1 vccd1 _8454_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6880_ _7028_/A _6880_/A2 _6906_/A3 _6879_/X vssd1 vssd1 vccd1 vccd1 _6880_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6566__A2 _6592_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4026__B1 _4071_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5831_ _6298_/A _6318_/A _6262_/A _6281_/A _5744_/S _5860_/S vssd1 vssd1 vccd1 vccd1
+ _5831_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_119_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5762_ _6163_/A _5762_/B vssd1 vssd1 vccd1 vccd1 _5762_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7501_ _7501_/CLK _7501_/D vssd1 vssd1 vccd1 vccd1 _7501_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4713_ _8483_/Q _8415_/Q _8447_/Q _8321_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4713_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5693_ _5881_/C _6008_/B vssd1 vssd1 vccd1 vccd1 _5786_/B sky130_fd_sc_hd__nor2_2
X_8481_ _8481_/CLK _8481_/D vssd1 vssd1 vccd1 vccd1 _8481_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4644_ _4643_/X _4642_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4644_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_7432_ _8354_/CLK _7432_/D vssd1 vssd1 vccd1 vccd1 _7432_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7363_ _8326_/CLK _7363_/D vssd1 vssd1 vccd1 vccd1 _7363_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold712 _5368_/X vssd1 vssd1 vccd1 vccd1 _7595_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold701 _7464_/Q vssd1 vssd1 vccd1 vccd1 hold701/X sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ _4574_/X _4571_/X _7365_/Q vssd1 vssd1 vccd1 vccd1 _7507_/D sky130_fd_sc_hd__mux2_1
X_7294_ _8368_/CLK _7294_/D _7104_/Y vssd1 vssd1 vccd1 vccd1 _7294_/Q sky130_fd_sc_hd__dfrtp_4
Xhold723 _8134_/Q vssd1 vssd1 vccd1 vccd1 hold723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 _6752_/X vssd1 vssd1 vccd1 vccd1 _8303_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6314_ _6297_/Y _6301_/B _6299_/B vssd1 vssd1 vccd1 vccd1 _6320_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold745 _7495_/Q vssd1 vssd1 vccd1 vccd1 hold745/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__7017__A _7017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold767 _8262_/Q vssd1 vssd1 vccd1 vccd1 hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _5326_/X vssd1 vssd1 vccd1 vccd1 _7557_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6245_ _6245_/A vssd1 vssd1 vccd1 vccd1 _6246_/B sky130_fd_sc_hd__inv_2
Xhold756 _6737_/X vssd1 vssd1 vccd1 vccd1 _8292_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold789 _7592_/Q vssd1 vssd1 vccd1 vccd1 hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold1401 _4418_/X vssd1 vssd1 vccd1 vccd1 _4420_/B1 sky130_fd_sc_hd__dlygate4sd3_1
X_6176_ _6176_/A _6176_/B vssd1 vssd1 vccd1 vccd1 _6177_/B sky130_fd_sc_hd__nand2_1
X_5127_ _5443_/A _7030_/C vssd1 vssd1 vccd1 vccd1 _5127_/X sky130_fd_sc_hd__or2_1
Xhold1423 _4358_/X vssd1 vssd1 vccd1 vccd1 _4372_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _4393_/X vssd1 vssd1 vccd1 vccd1 _8379_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1412 _8381_/Q vssd1 vssd1 vccd1 vccd1 _5050_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1467 _7286_/Q vssd1 vssd1 vccd1 vccd1 _5128_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 _7033_/Y vssd1 vssd1 vccd1 vccd1 _8489_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _5058_/A1 _5069_/S _5182_/B1 _5057_/X vssd1 vssd1 vccd1 vccd1 _7341_/D sky130_fd_sc_hd__o211a_1
Xhold1456 _4243_/Y vssd1 vssd1 vccd1 vccd1 _4244_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 _7836_/Q vssd1 vssd1 vccd1 vccd1 _6457_/A0 sky130_fd_sc_hd__dlygate4sd3_1
X_4009_ _3923_/B _7947_/Q vssd1 vssd1 vccd1 vccd1 _4009_/X sky130_fd_sc_hd__and2b_1
Xhold1478 hold1819/X vssd1 vssd1 vccd1 vccd1 _7079_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_64_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _8364_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5000__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4663__S1 _4733_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5780__A3 _6035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5670__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4985__S _7057_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5048__A2 _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6340__S1 _5860_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output119_A _7313_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_55_clk clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 _8079_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4654__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5220__A2 _5188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _7898_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _7052_/A _7732_/Q _7735_/Q _3647_/Y vssd1 vssd1 vccd1 vccd1 _4360_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6720__A2 _6705_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5580__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4291_ _8497_/Q _4292_/B vssd1 vssd1 vccd1 vccd1 _4291_/Y sky130_fd_sc_hd__nor2_1
X_6030_ _6030_/A1 _6018_/Y _6029_/X _6163_/A vssd1 vssd1 vccd1 vccd1 _6030_/X sky130_fd_sc_hd__o22a_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5287__A2 _5294_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4590__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3812__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6236__A1 _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7981_ _8510_/CLK _7981_/D vssd1 vssd1 vccd1 vccd1 _7981_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clkbuf_4_13_0_clk/X vssd1 vssd1 vccd1 vccd1 _8517_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_6932_ _7023_/A _6932_/A2 _6970_/A3 _6931_/X vssd1 vssd1 vccd1 vccd1 _6932_/X sky130_fd_sc_hd__a31o_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6863_ _6929_/A _6901_/B vssd1 vssd1 vccd1 vccd1 _6863_/X sky130_fd_sc_hd__and2_1
XFILLER_0_76_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5814_ _6008_/A _5814_/B vssd1 vssd1 vccd1 vccd1 _5815_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_8_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5211__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6794_ _6706_/A _6794_/A2 _6779_/B _6793_/X vssd1 vssd1 vccd1 vccd1 _6794_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5745_ _6157_/A _6175_/A _6191_/A _6209_/A _5744_/S _5859_/S vssd1 vssd1 vccd1 vccd1
+ _5745_/X sky130_fd_sc_hd__mux4_1
X_8464_ _8464_/CLK _8464_/D vssd1 vssd1 vccd1 vccd1 _8464_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout317_A _4080_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5676_ _6550_/A _5676_/B vssd1 vssd1 vccd1 vccd1 _5676_/X sky130_fd_sc_hd__and2_1
XFILLER_0_115_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5474__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7415_ _8475_/CLK _7415_/D vssd1 vssd1 vccd1 vccd1 _7415_/Q sky130_fd_sc_hd__dfxtp_1
X_4627_ _4625_/X _4626_/X _5103_/A vssd1 vssd1 vccd1 vccd1 _4627_/X sky130_fd_sc_hd__mux2_1
X_8395_ _8463_/CLK _8395_/D vssd1 vssd1 vccd1 vccd1 _8395_/Q sky130_fd_sc_hd__dfxtp_1
Xhold520 _5294_/X vssd1 vssd1 vccd1 vccd1 _7498_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6711__A2 _6737_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold542 _5269_/X vssd1 vssd1 vccd1 vccd1 _7473_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _8171_/Q _8203_/Q _8267_/Q _7775_/Q _4696_/S0 _4740_/S1 vssd1 vssd1 vccd1
+ vccd1 _4558_/X sky130_fd_sc_hd__mux4_1
Xhold531 _7562_/Q vssd1 vssd1 vccd1 vccd1 hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _7594_/Q vssd1 vssd1 vccd1 vccd1 hold553/X sky130_fd_sc_hd__dlygate4sd3_1
X_7346_ _8020_/CLK _7346_/D vssd1 vssd1 vccd1 vccd1 _7346_/Q sky130_fd_sc_hd__dfxtp_2
Xhold597 _7478_/Q vssd1 vssd1 vccd1 vccd1 hold597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 _6751_/X vssd1 vssd1 vccd1 vccd1 _8302_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _5174_/A1 _4383_/B _5468_/C vssd1 vssd1 vccd1 vccd1 _7309_/D sky130_fd_sc_hd__mux2_1
Xhold575 _8305_/Q vssd1 vssd1 vccd1 vccd1 hold575/X sky130_fd_sc_hd__dlygate4sd3_1
X_7277_ _7279_/A vssd1 vssd1 vccd1 vccd1 _7277_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_40_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold564 _5290_/X vssd1 vssd1 vccd1 vccd1 _7494_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5278__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6228_ _6211_/A _6210_/A _6208_/Y vssd1 vssd1 vccd1 vccd1 _6229_/B sky130_fd_sc_hd__a21o_1
X_6159_ _6159_/A _6159_/B vssd1 vssd1 vccd1 vccd1 _6159_/X sky130_fd_sc_hd__xor2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1220 _6618_/X vssd1 vssd1 vccd1 vccd1 _8173_/D sky130_fd_sc_hd__dlygate4sd3_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1242 _6946_/X vssd1 vssd1 vccd1 vccd1 _8438_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 _8418_/Q vssd1 vssd1 vccd1 vccd1 _6904_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6322__S1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1275 _7039_/Y vssd1 vssd1 vccd1 vccd1 _8492_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 _8350_/Q vssd1 vssd1 vccd1 vccd1 _6826_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 _6662_/X vssd1 vssd1 vccd1 vccd1 _8195_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_37_clk clkbuf_4_11_0_clk/X vssd1 vssd1 vccd1 vccd1 _8458_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1286 _8194_/Q vssd1 vssd1 vccd1 vccd1 _6660_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1297 _6656_/X vssd1 vssd1 vccd1 vccd1 _8192_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4884__S1 _4990_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5202__A2 _5221_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5833__S0 _5744_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4636__S1 _4731_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5665__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6702__A2 _6669_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6496__A _6520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 _8129_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[28] sky130_fd_sc_hd__buf_12
XANTENNA__5269__A2 _5262_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput73 _8119_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[18] sky130_fd_sc_hd__buf_12
Xoutput95 _8110_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[9] sky130_fd_sc_hd__buf_12
XANTENNA_clkbuf_leaf_94_clk_A clkbuf_4_4_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4572__S0 _4727_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6943__B _6943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6769__A2 _6773_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4744__A _7006_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 _8465_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4875__S1 _4952_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7120__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3860_ _4067_/A_N _7959_/Q vssd1 vssd1 vccd1 vccd1 _3860_/X sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_32_clk_A clkbuf_4_10_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3791_ _8086_/Q _3790_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _6815_/A sky130_fd_sc_hd__mux2_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5530_ _8249_/Q _5541_/B _5541_/C vssd1 vssd1 vccd1 vccd1 _7719_/D sky130_fd_sc_hd__and3_1
XFILLER_0_42_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5575__A _6551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5461_ _5461_/A _5540_/B _5540_/C vssd1 vssd1 vccd1 vccd1 _5461_/X sky130_fd_sc_hd__and3_1
XFILLER_0_26_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_A clkbuf_4_14_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4412_ _4412_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4412_/X sky130_fd_sc_hd__and2_1
X_7244__122 _8195_/CLK vssd1 vssd1 vccd1 vccd1 _8254_/CLK sky130_fd_sc_hd__inv_2
X_5392_ _7346_/Q _5392_/B _5408_/B vssd1 vssd1 vccd1 vccd1 _5392_/X sky130_fd_sc_hd__or3b_1
X_8180_ _8402_/CLK _8180_/D vssd1 vssd1 vccd1 vccd1 _8180_/Q sky130_fd_sc_hd__dfxtp_1
X_4343_ _8490_/Q _4343_/B vssd1 vssd1 vccd1 vccd1 _4344_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout329 _6913_/A vssd1 vssd1 vccd1 vccd1 _6847_/A sky130_fd_sc_hd__clkbuf_8
Xfanout307 _5333_/Y vssd1 vssd1 vccd1 vccd1 _5367_/A2 sky130_fd_sc_hd__buf_6
X_7062_ _7071_/B _7061_/Y _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8503_/D sky130_fd_sc_hd__a21oi_1
Xfanout318 _4069_/X vssd1 vssd1 vccd1 vccd1 _6939_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4274_ _4274_/A _4274_/B vssd1 vssd1 vccd1 vccd1 _4274_/X sky130_fd_sc_hd__xor2_1
X_6013_ _6013_/A _6094_/B vssd1 vssd1 vccd1 vccd1 _6016_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4563__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_105_clk_A clkbuf_4_1_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6853__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5968__B1 _7258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_19_clk clkbuf_4_8_0_clk/X vssd1 vssd1 vccd1 vccd1 _8481_/CLK sky130_fd_sc_hd__clkbuf_16
X_7964_ _8096_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 _7964_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6915_ _6915_/A _6963_/B vssd1 vssd1 vccd1 vccd1 _6915_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout267_A _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7030__A _7031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5469__B _5470_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7895_ _8504_/CLK _7895_/D vssd1 vssd1 vccd1 vccd1 _7895_/Q sky130_fd_sc_hd__dfxtp_1
X_6846_ _6999_/A _6846_/A2 _6845_/B _6845_/Y vssd1 vssd1 vccd1 vccd1 _6846_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout434_A _6660_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5196__A1 _6921_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6777_ _6777_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6777_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4618__S1 _4740_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8516_ _8519_/CLK _8516_/D vssd1 vssd1 vccd1 vccd1 _8516_/Q sky130_fd_sc_hd__dfxtp_1
X_3989_ _7705_/Q _4081_/B vssd1 vssd1 vccd1 vccd1 _3989_/X sky130_fd_sc_hd__or2_1
X_5728_ _5734_/A _6380_/A vssd1 vssd1 vccd1 vccd1 _5728_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3746__A2 _6448_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5659_ _6494_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5659_/X sky130_fd_sc_hd__and2_1
XANTENNA__6696__A1 _6959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8447_ _8483_/CLK _8447_/D vssd1 vssd1 vccd1 vccd1 _8447_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6160__A3 _6115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_8378_ _8378_/CLK _8378_/D _7272_/Y vssd1 vssd1 vccd1 vccd1 _8378_/Q sky130_fd_sc_hd__dfrtp_1
Xhold361 _5304_/X vssd1 vssd1 vccd1 vccd1 _7535_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold350 _7341_/Q vssd1 vssd1 vccd1 vccd1 _5438_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7329_ _8379_/CLK _7329_/D vssd1 vssd1 vccd1 vccd1 _7329_/Q sky130_fd_sc_hd__dfxtp_1
Xhold383 _5450_/X vssd1 vssd1 vccd1 vccd1 _7639_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 _7493_/Q vssd1 vssd1 vccd1 vccd1 hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _7456_/Q vssd1 vssd1 vccd1 vccd1 hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5120__A1 input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_13_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_4_13_0_clk/X sky130_fd_sc_hd__clkbuf_8
Xhold1050 _5268_/X vssd1 vssd1 vccd1 vccd1 _7472_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _7007_/X vssd1 vssd1 vccd1 vccd1 _8465_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1061 _7470_/Q vssd1 vssd1 vccd1 vccd1 _5266_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5959__B1 _6413_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1094 _5271_/X vssd1 vssd1 vccd1 vccd1 _7475_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3682__B2 _8028_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1083 _7408_/Q vssd1 vssd1 vccd1 vccd1 _5194_/B2 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6620__A1 _4775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4857__S1 _4987_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7228__106 _8464_/CLK vssd1 vssd1 vccd1 vccd1 _8238_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6687__A1 _6941_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4793__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__7115__A _7267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4545__S0 _4640_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4474__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4961_ _8192_/Q _8224_/Q _8288_/Q _7796_/Q _4990_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4961_/X sky130_fd_sc_hd__mux4_1
X_7680_ _8339_/CLK _7680_/D vssd1 vssd1 vccd1 vccd1 _7680_/Q sky130_fd_sc_hd__dfxtp_1
X_3912_ _7973_/Q _4079_/A2 _4079_/B1 _8005_/Q _3911_/X vssd1 vssd1 vccd1 vccd1 _3912_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_80_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4892_ _8472_/Q _8404_/Q _8436_/Q _8310_/Q _4987_/S0 _4987_/S1 vssd1 vssd1 vccd1
+ vccd1 _4892_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3976__A2 _4079_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6700_ _6967_/A _6701_/A2 _6701_/B1 _6700_/B2 vssd1 vssd1 vccd1 vccd1 _6700_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6631_ _6937_/A _6661_/B vssd1 vssd1 vccd1 vccd1 _6631_/X sky130_fd_sc_hd__and2_1
X_3843_ _6126_/A vssd1 vssd1 vccd1 vccd1 _5955_/A sky130_fd_sc_hd__inv_2
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6562_ _3939_/C _6592_/A2 _6592_/B1 hold723/X vssd1 vssd1 vccd1 vccd1 _6562_/X sky130_fd_sc_hd__a22o_1
X_3774_ _3968_/A _3774_/A2 _3773_/X vssd1 vssd1 vccd1 vccd1 _6154_/A sky130_fd_sc_hd__a21bo_2
X_8301_ _8427_/CLK _8301_/D vssd1 vssd1 vccd1 vccd1 _8301_/Q sky130_fd_sc_hd__dfxtp_1
X_7184__62 _8460_/CLK vssd1 vssd1 vccd1 vccd1 _8064_/CLK sky130_fd_sc_hd__inv_2
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5513_ _8232_/Q _5542_/B _5542_/C vssd1 vssd1 vccd1 vccd1 _7702_/D sky130_fd_sc_hd__and3_1
XFILLER_0_89_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6493_ _6539_/A _6493_/B vssd1 vssd1 vccd1 vccd1 _6493_/X sky130_fd_sc_hd__and2_1
XFILLER_0_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7126__4 _8339_/CLK vssd1 vssd1 vccd1 vccd1 _7503_/CLK sky130_fd_sc_hd__inv_2
X_8232_ _8232_/CLK _8232_/D vssd1 vssd1 vccd1 vccd1 _8232_/Q sky130_fd_sc_hd__dfxtp_1
X_5444_ _5444_/A _7082_/A _7082_/B vssd1 vssd1 vccd1 vccd1 _5444_/X sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_8_clk clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _8319_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__6678__A1 _6923_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8163_ _8484_/CLK _8163_/D vssd1 vssd1 vccd1 vccd1 _8163_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4784__S0 _5475_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5375_ _7082_/A _7082_/B _6981_/A vssd1 vssd1 vccd1 vccd1 _6600_/A sky130_fd_sc_hd__and3_1
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__7025__A _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7114_ _7267_/A vssd1 vssd1 vccd1 vccd1 _7114_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4326_ _5575_/B _5052_/A1 _5465_/B vssd1 vssd1 vccd1 vccd1 _4385_/B sky130_fd_sc_hd__mux2_1
X_8094_ _8382_/CLK _8128_/D vssd1 vssd1 vccd1 vccd1 _8094_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout384_A _7050_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout159 _5370_/Y vssd1 vssd1 vccd1 vccd1 _7064_/B1 sky130_fd_sc_hd__buf_4
X_7045_ _7031_/Y _7045_/A2 _7064_/B1 vssd1 vssd1 vccd1 vccd1 _8495_/D sky130_fd_sc_hd__a21oi_1
X_4257_ _8502_/Q _4257_/B vssd1 vssd1 vccd1 vccd1 _4257_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__6850__A1 _7010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5653__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4188_ _4186_/Y _4188_/B vssd1 vssd1 vccd1 vccd1 _4190_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__4839__S1 _4896_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7947_ _8365_/CLK _7947_/D vssd1 vssd1 vccd1 vccd1 _7947_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_7878_ _8464_/CLK _7878_/D vssd1 vssd1 vccd1 vccd1 _7878_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__A2 _4073_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6829_ _6961_/A _6837_/B vssd1 vssd1 vccd1 vccd1 _6829_/X sky130_fd_sc_hd__and2_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3680__A_N _4067_/A_N vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3719__A2 _4071_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5341__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold180 _7849_/Q vssd1 vssd1 vccd1 vccd1 _6470_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold191 _6420_/X vssd1 vssd1 vccd1 vccd1 _7902_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4527__S0 _7072_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5644__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3958__A2 _4084_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4080__A1 _4079_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6357__A0 _6298_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4233__S _5453_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6014__A _6016_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6109__B1 _6108_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6949__A _6949_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5332__A1 _6971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4469__A _7018_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5883__A2 _6398_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5160_ _5160_/A1 _4416_/B _5166_/B1 _5159_/X vssd1 vssd1 vccd1 vccd1 _7392_/D sky130_fd_sc_hd__o211a_1
XANTENNA__7085__B2 _5473_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4111_ _4105_/X _4109_/X _4110_/Y _4092_/C vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__a31o_1
Xhold1808 _7879_/Q vssd1 vssd1 vccd1 vccd1 hold1808/X sky130_fd_sc_hd__dlygate4sd3_1
X_5091_ _7061_/A _5465_/C vssd1 vssd1 vccd1 vccd1 _5091_/X sky130_fd_sc_hd__or2_1
XANTENNA__5635__A2 _5620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4042_ _5993_/A _5990_/A vssd1 vssd1 vccd1 vccd1 _4044_/A sky130_fd_sc_hd__or2_1
Xhold1819 _7367_/Q vssd1 vssd1 vccd1 vccd1 hold1819/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5096__B1 _5172_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6832__A1 _7025_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6045__C1 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5993_ _5993_/A _5993_/B vssd1 vssd1 vccd1 vccd1 _5994_/B sky130_fd_sc_hd__nor2_1
X_7801_ _8451_/CLK _7801_/D vssd1 vssd1 vccd1 vccd1 _7801_/Q sky130_fd_sc_hd__dfxtp_1
X_7732_ _8079_/CLK _7732_/D vssd1 vssd1 vccd1 vccd1 _7732_/Q sky130_fd_sc_hd__dfxtp_1
X_4944_ _8350_/Q _7826_/Q _7492_/Q _7460_/Q _4983_/S0 _4969_/S1 vssd1 vssd1 vccd1
+ vccd1 _4944_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7663_ _8079_/CLK _7663_/D vssd1 vssd1 vccd1 vccd1 _7663_/Q sky130_fd_sc_hd__dfxtp_1
X_4875_ _8147_/Q _7546_/Q _7418_/Q _7578_/Q _4997_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4875_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_47_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5020__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6614_ _7015_/A _6614_/A2 _6605_/B _6613_/X vssd1 vssd1 vccd1 vccd1 _6614_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7594_ _8467_/CLK _7594_/D vssd1 vssd1 vccd1 vccd1 _7594_/Q sky130_fd_sc_hd__dfxtp_1
X_3826_ _8096_/Q _3825_/X _4069_/S vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6859__A _6925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3982__S _4074_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4374__A2 _5182_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3757_ _4074_/S _3757_/B vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__nand2_1
X_6545_ _6545_/A _6545_/B vssd1 vssd1 vccd1 vccd1 _8027_/D sky130_fd_sc_hd__and2_1
XFILLER_0_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3688_ _7662_/Q _7836_/Q vssd1 vssd1 vccd1 vccd1 _3688_/X sky130_fd_sc_hd__and2b_1
X_8215_ _8461_/CLK _8215_/D vssd1 vssd1 vccd1 vccd1 _8215_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5482__B _5542_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6476_ _7027_/A _6476_/B vssd1 vssd1 vccd1 vccd1 _6476_/X sky130_fd_sc_hd__and2_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5323__A1 _6953_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5427_ _5427_/A _7030_/B _5463_/C vssd1 vssd1 vccd1 vccd1 _5427_/X sky130_fd_sc_hd__and3_1
X_8146_ _8328_/CLK _8146_/D vssd1 vssd1 vccd1 vccd1 _8146_/Q sky130_fd_sc_hd__dfxtp_1
X_5358_ _6951_/A _5335_/B _5368_/B1 hold441/X vssd1 vssd1 vccd1 vccd1 _5358_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8077_ _8464_/CLK _8111_/D vssd1 vssd1 vccd1 vccd1 _8077_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3885__B2 _8024_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4309_ _4298_/Y _4302_/B _4300_/B vssd1 vssd1 vccd1 vccd1 _4310_/B sky130_fd_sc_hd__o21a_1
XANTENNA__6593__C_N _7069_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5289_ _6959_/A _5262_/B _5295_/B1 hold372/X vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__a22o_1
X_7028_ _7028_/A _7028_/B vssd1 vssd1 vccd1 vccd1 _7028_/X sky130_fd_sc_hd__and2_1
XANTENNA__5626__A2 _5652_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6587__B1 _6591_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6339__B1 _6391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4053__S _4085_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4996__S0 _4996_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4988__S _4988_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3905__B _8516_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5865__A2 _6063_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5078__B1 _5146_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5617__A2 _5584_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6814__A1 _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6290__A2 _6309_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4920__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6578__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6951__B _6963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4752__A _6498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4053__A1 _4052_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5250__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4660_ _8346_/Q _7822_/Q _7488_/Q _7456_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4660_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4591_ _8143_/Q _7542_/Q _7414_/Q _7574_/Q _4640_/S0 _4639_/S1 vssd1 vssd1 vccd1
+ vccd1 _4591_/X sky130_fd_sc_hd__mux4_1
X_7154__32 _8487_/CLK vssd1 vssd1 vccd1 vccd1 _7531_/CLK sky130_fd_sc_hd__inv_2
X_6330_ _3725_/A _6292_/A _6329_/X _7279_/A vssd1 vssd1 vccd1 vccd1 _7894_/D sky130_fd_sc_hd__a211oi_1
XANTENNA__6750__B1 _6773_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4987__S0 _4987_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold927 _7453_/Q vssd1 vssd1 vccd1 vccd1 hold927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 _5314_/X vssd1 vssd1 vccd1 vccd1 _7545_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold905 _8213_/Q vssd1 vssd1 vccd1 vccd1 hold905/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold938 _6573_/X vssd1 vssd1 vccd1 vccd1 _8145_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3815__B _4072_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6261_ _6262_/A _6262_/B vssd1 vssd1 vccd1 vccd1 _6261_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5305__A1 _6917_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold949 _7558_/Q vssd1 vssd1 vccd1 vccd1 hold949/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5856__A2 _5892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6192_ _6192_/A _6192_/B vssd1 vssd1 vccd1 vccd1 _6194_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3867__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5212_ _6953_/A _5188_/B _5220_/B1 hold849/X vssd1 vssd1 vccd1 vccd1 _5212_/X sky130_fd_sc_hd__a22o_1
X_8000_ _8385_/CLK _8000_/D vssd1 vssd1 vccd1 vccd1 _8000_/Q sky130_fd_sc_hd__dfxtp_1
X_5143_ _5451_/A _5451_/C vssd1 vssd1 vccd1 vccd1 _5143_/X sky130_fd_sc_hd__or2_1
XANTENNA__7058__A1 _7071_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1605 _7345_/Q vssd1 vssd1 vccd1 vccd1 _5404_/A sky130_fd_sc_hd__buf_2
XANTENNA__5069__A0 input26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1616 _7675_/Q vssd1 vssd1 vccd1 vccd1 _3981_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3831__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5608__A2 _5616_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1649 _7344_/Q vssd1 vssd1 vccd1 vccd1 _5404_/B sky130_fd_sc_hd__clkbuf_2
Xhold1627 _4202_/Y vssd1 vssd1 vccd1 vccd1 _4203_/B sky130_fd_sc_hd__dlygate4sd3_1
X_5074_ input28/X _5085_/B _5140_/B1 _5073_/Y vssd1 vssd1 vccd1 vccd1 _7349_/D sky130_fd_sc_hd__o211a_1
Xhold1638 _7048_/Y vssd1 vssd1 vccd1 vccd1 _7049_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4025_ _7711_/Q _4070_/B vssd1 vssd1 vccd1 vccd1 _4025_/X sky130_fd_sc_hd__or2_1
XANTENNA__6569__B1 _6592_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6861__B _6901_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3977__S _4069_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5241__B1 _5259_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5976_ _5976_/A _5976_/B vssd1 vssd1 vccd1 vccd1 _5976_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5477__B _7088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4927_ _8477_/Q _8409_/Q _8441_/Q _8315_/Q _4996_/S0 _4952_/S1 vssd1 vssd1 vccd1
+ vccd1 _4927_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_47_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7715_ _8484_/CLK _7715_/D vssd1 vssd1 vccd1 vccd1 _7715_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4858_ _4857_/X _4856_/X _4988_/S vssd1 vssd1 vccd1 vccd1 _4858_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7646_ _8501_/CLK _7646_/D vssd1 vssd1 vccd1 vccd1 _7646_/Q sky130_fd_sc_hd__dfxtp_1
X_3809_ _6388_/A _6386_/A vssd1 vssd1 vccd1 vccd1 _3811_/A sky130_fd_sc_hd__or2_1
X_4789_ _4788_/X _4785_/X _4929_/S vssd1 vssd1 vccd1 vccd1 _8231_/D sky130_fd_sc_hd__mux2_1
X_7577_ _8473_/CLK _7577_/D vssd1 vssd1 vccd1 vccd1 _7577_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6528_ _7018_/A _6528_/B vssd1 vssd1 vccd1 vccd1 _8010_/D sky130_fd_sc_hd__and2_1
X_6459_ _6498_/A hold75/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__and2_1
X_8129_ _8129_/CLK _8129_/D vssd1 vssd1 vccd1 vccd1 _8129_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4048__S _4080_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6272__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4902__S0 _5089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5668__A _6552_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6024__A2 _5993_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5232__B1 _5258_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6499__A _6534_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6732__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4969__S0 _4983_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__A _7029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__7123__A _7279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5578__A _6539_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5830_ _6191_/A _6209_/A _6226_/A _6244_/A _5744_/S _5859_/S vssd1 vssd1 vccd1 vccd1
+ _5830_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5761_ _5881_/C _5755_/X _5760_/Y _6008_/B vssd1 vssd1 vccd1 vccd1 _5762_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_7500_ _7500_/CLK _7500_/D vssd1 vssd1 vccd1 vccd1 _7500_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_8480_ _8480_/CLK _8480_/D vssd1 vssd1 vccd1 vccd1 _8480_/Q sky130_fd_sc_hd__dfxtp_1
X_4712_ _8193_/Q _8225_/Q _8289_/Q _7797_/Q _4727_/S0 _4727_/S1 vssd1 vssd1 vccd1
+ vccd1 _4712_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5692_ _5723_/B _5727_/C vssd1 vssd1 vccd1 vccd1 _6129_/B sky130_fd_sc_hd__or2_4
XFILLER_0_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_7431_ _8160_/CLK _7431_/D vssd1 vssd1 vccd1 vccd1 _7431_/Q sky130_fd_sc_hd__dfxtp_1
X_4643_ _8473_/Q _8405_/Q _8437_/Q _8311_/Q _4696_/S0 _4737_/S1 vssd1 vssd1 vccd1
+ vccd1 _4643_/X sky130_fd_sc_hd__mux4_1
XANTENNA__6723__B1 _6738_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold702 _5256_/X vssd1 vssd1 vccd1 vccd1 _7464_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7362_ _8448_/CLK _7362_/D vssd1 vssd1 vccd1 vccd1 _7362_/Q sky130_fd_sc_hd__dfxtp_4
X_4574_ _4573_/X _4572_/X _7048_/A vssd1 vssd1 vccd1 vccd1 _4574_/X sky130_fd_sc_hd__mux2_1
X_7293_ _8507_/CLK _7293_/D _7103_/Y vssd1 vssd1 vccd1 vccd1 _7293_/Q sky130_fd_sc_hd__dfrtp_4
Xhold724 _6562_/X vssd1 vssd1 vccd1 vccd1 _8134_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6313_ _3714_/B _6292_/A _6312_/X _6347_/B1 vssd1 vssd1 vccd1 vccd1 _7893_/D sky130_fd_sc_hd__a211oi_2
Xhold735 _7434_/Q vssd1 vssd1 vccd1 vccd1 hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 _7556_/Q vssd1 vssd1 vccd1 vccd1 hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _5291_/X vssd1 vssd1 vccd1 vccd1 _7495_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 _6707_/X vssd1 vssd1 vccd1 vccd1 _8262_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold757 _8203_/Q vssd1 vssd1 vccd1 vccd1 hold757/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 _7786_/Q vssd1 vssd1 vccd1 vccd1 hold779/X sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ _6244_/A _6244_/B vssd1 vssd1 vccd1 vccd1 _6245_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout297_A _6557_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6175_ _6175_/A _6175_/B vssd1 vssd1 vccd1 vccd1 _6176_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold1402 hold1405/X vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__clkbuf_2
X_5126_ _5126_/A1 _4448_/B _5140_/B1 _5125_/X vssd1 vssd1 vccd1 vccd1 _7375_/D sky130_fd_sc_hd__o211a_1
Xhold1424 _7656_/Q vssd1 vssd1 vccd1 vccd1 _4336_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1413 _4327_/C vssd1 vssd1 vccd1 vccd1 _4387_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 _7291_/Q vssd1 vssd1 vccd1 vccd1 _5138_/A1 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1446 _7285_/Q vssd1 vssd1 vccd1 vccd1 _5126_/A1 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6254__A2 _6414_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5057_ _5438_/A _5470_/C vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__or2_1
Xhold1435 _7645_/Q vssd1 vssd1 vccd1 vccd1 _4257_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 _4244_/Y vssd1 vssd1 vccd1 vccd1 _4246_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4008_ _4008_/A _4008_/B vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__and2_1
XFILLER_0_79_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout464_A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1479 _7042_/Y vssd1 vssd1 vccd1 vccd1 _7043_/A2 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5214__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5959_ _3985_/A _6398_/A2 _6413_/B1 _5943_/A _6063_/A vssd1 vssd1 vccd1 vccd1 _5959_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold1481_A _7299_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_7629_ _8500_/CLK _7629_/D vssd1 vssd1 vccd1 vccd1 _7629_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__6714__B1 _6737_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold1746_A _7359_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5951__A _6411_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6796__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4506__S _5449_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5205__B1 _5220_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3646__A _7273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6181__A1 _5740_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__7118__A _7281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output93_A _8108_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 _3999_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _4401_/A _4397_/B vssd1 vssd1 vccd1 vccd1 _4398_/A sky130_fd_sc_hd__and2_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4590__S1 _4639_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clkbuf_4_2_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7980_ _8364_/CLK hold95/X vssd1 vssd1 vccd1 vccd1 _7980_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6931_ _6931_/A _6969_/B vssd1 vssd1 vccd1 vccd1 _6931_/X sky130_fd_sc_hd__and2_1
X_6862_ _7007_/A _6862_/A2 _6845_/B _6861_/X vssd1 vssd1 vccd1 vccd1 _6862_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_107_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5101__A _5472_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5813_ _5952_/A _5812_/X _5803_/Y vssd1 vssd1 vccd1 vccd1 _5814_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6793_ _6925_/A _6839_/B vssd1 vssd1 vccd1 vccd1 _6793_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5744_ _6157_/A _6175_/A _5744_/S vssd1 vssd1 vccd1 vccd1 _5744_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_8463_ _8463_/CLK _8463_/D vssd1 vssd1 vccd1 vccd1 _8463_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5675_ _7027_/A _5675_/B vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__and2_1
X_8394_ _8426_/CLK _8394_/D vssd1 vssd1 vccd1 vccd1 _8394_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5474__C _7088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_7414_ _8343_/CLK _7414_/D vssd1 vssd1 vccd1 vccd1 _7414_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout212_A _5538_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4626_ _8148_/Q _7547_/Q _7419_/Q _7579_/Q _4706_/S0 _4733_/S1 vssd1 vssd1 vccd1
+ vccd1 _4626_/X sky130_fd_sc_hd__mux4_1
XANTENNA__7028__A _7028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold510 _6759_/X vssd1 vssd1 vccd1 vccd1 _8310_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7345_ _7903_/CLK _7345_/D vssd1 vssd1 vccd1 vccd1 _7345_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_130_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold543 _7404_/Q vssd1 vssd1 vccd1 vccd1 hold543/X sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ _4555_/X _4556_/X _4742_/S vssd1 vssd1 vccd1 vccd1 _4557_/X sky130_fd_sc_hd__mux2_1
Xhold532 _5331_/X vssd1 vssd1 vccd1 vccd1 _7562_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _5367_/X vssd1 vssd1 vccd1 vccd1 _7594_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold521 _7488_/Q vssd1 vssd1 vccd1 vccd1 hold521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _7816_/Q vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _8217_/Q vssd1 vssd1 vccd1 vccd1 hold587/X sky130_fd_sc_hd__dlygate4sd3_1
X_4488_ _5176_/A1 _4341_/C _5468_/C vssd1 vssd1 vccd1 vccd1 _7310_/D sky130_fd_sc_hd__mux2_1
Xhold576 _6754_/X vssd1 vssd1 vccd1 vccd1 _8305_/D sky130_fd_sc_hd__dlygate4sd3_1
X_7276_ _7281_/A vssd1 vssd1 vccd1 vccd1 _7276_/Y sky130_fd_sc_hd__inv_2
Xhold598 _5274_/X vssd1 vssd1 vccd1 vccd1 _7478_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5490__B _5541_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6227_ _6227_/A _6227_/B vssd1 vssd1 vccd1 vccd1 _6229_/A sky130_fd_sc_hd__nor2_1
X_6158_ _6142_/A _6141_/A _6139_/Y vssd1 vssd1 vccd1 vccd1 _6159_/B sky130_fd_sc_hd__a21o_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _8398_/Q vssd1 vssd1 vccd1 vccd1 _6864_/A2 sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _7079_/A _7030_/C vssd1 vssd1 vccd1 vccd1 _5109_/X sky130_fd_sc_hd__or2_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1210 _6888_/X vssd1 vssd1 vccd1 vccd1 _8410_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 _8181_/Q vssd1 vssd1 vccd1 vccd1 _6634_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 _6904_/X vssd1 vssd1 vccd1 vccd1 _8418_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6778__A3 _6779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5710__S _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6089_ _6128_/A _6088_/X _6362_/C _5899_/B vssd1 vssd1 vccd1 vccd1 _6089_/X sky130_fd_sc_hd__a2bb2o_1
Xhold1265 _8414_/Q vssd1 vssd1 vccd1 vccd1 _6896_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _8392_/Q vssd1 vssd1 vccd1 vccd1 _6852_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1254 _6826_/X vssd1 vssd1 vccd1 vccd1 _8350_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold1298 _8169_/Q vssd1 vssd1 vccd1 vccd1 _6610_/A2 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1287 _6660_/X vssd1 vssd1 vccd1 vccd1 _8194_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4326__S _5465_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5946__A _5946_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5833__S1 _5859_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6950__A3 _6970_/A3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6777__A _6777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5681__A _6524_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput74 _8120_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[19] sky130_fd_sc_hd__buf_12
Xoutput85 _8130_/Q vssd1 vssd1 vccd1 vccd1 o_data_addr_M[29] sky130_fd_sc_hd__buf_12
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput96 _8099_/Q vssd1 vssd1 vccd1 vccd1 o_mem_write_M sky130_fd_sc_hd__buf_12
XANTENNA__4572__S1 _4727_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4760__A _7026_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3790_ _7990_/Q _4068_/A2 _4068_/B1 _8022_/Q _3789_/X vssd1 vssd1 vccd1 vccd1 _3790_/X
+ sky130_fd_sc_hd__a221o_2
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5067__S _5067_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5460_ hold43/X _5465_/B _5463_/C vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__and3_1
X_4411_ _5034_/A1 _4416_/B _4409_/X _4410_/Y vssd1 vssd1 vccd1 vccd1 _8373_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5391_ _5391_/A _5408_/C _5408_/B vssd1 vssd1 vccd1 vccd1 _6975_/C sky130_fd_sc_hd__nor3b_4
XFILLER_0_50_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3912__B1 _4079_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ _8490_/Q _4343_/B vssd1 vssd1 vccd1 vccd1 _4342_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout319 _4057_/X vssd1 vssd1 vccd1 vccd1 _6933_/A sky130_fd_sc_hd__buf_4
Xfanout308 _5333_/Y vssd1 vssd1 vccd1 vccd1 _5335_/B sky130_fd_sc_hd__clkbuf_8
X_7061_ _7061_/A _7069_/B vssd1 vssd1 vccd1 vccd1 _7061_/Y sky130_fd_sc_hd__nand2_1
X_4273_ _4263_/Y _4267_/B _4265_/B vssd1 vssd1 vccd1 vccd1 _4274_/B sky130_fd_sc_hd__o21a_1
X_6012_ _5992_/Y _5996_/B _5994_/B vssd1 vssd1 vccd1 vccd1 _6018_/A sky130_fd_sc_hd__a21o_1
.ends

