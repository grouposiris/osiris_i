magic
tech sky130A
magscale 1 2
timestamp 1731114205
<< obsli1 >>
rect 2760 2703 32200 32113
<< obsm1 >>
rect 14 2672 34854 32360
<< metal2 >>
rect 662 33544 718 34344
rect 1950 33544 2006 34344
rect 3882 33544 3938 34344
rect 5170 33544 5226 34344
rect 6458 33544 6514 34344
rect 8390 33544 8446 34344
rect 9678 33544 9734 34344
rect 11610 33544 11666 34344
rect 12898 33544 12954 34344
rect 14186 33544 14242 34344
rect 16118 33544 16174 34344
rect 17406 33544 17462 34344
rect 18694 33544 18750 34344
rect 20626 33544 20682 34344
rect 21914 33544 21970 34344
rect 23846 33544 23902 34344
rect 25134 33544 25190 34344
rect 26422 33544 26478 34344
rect 28354 33544 28410 34344
rect 29642 33544 29698 34344
rect 31574 33544 31630 34344
rect 32862 33544 32918 34344
rect 34150 33544 34206 34344
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 4526 0 4582 800
rect 5814 0 5870 800
rect 7102 0 7158 800
rect 9034 0 9090 800
rect 10322 0 10378 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19338 0 19394 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28998 0 29054 800
rect 30286 0 30342 800
rect 32218 0 32274 800
rect 33506 0 33562 800
rect 34794 0 34850 800
<< obsm2 >>
rect 20 33488 606 34105
rect 774 33488 1894 34105
rect 2062 33488 3826 34105
rect 3994 33488 5114 34105
rect 5282 33488 6402 34105
rect 6570 33488 8334 34105
rect 8502 33488 9622 34105
rect 9790 33488 11554 34105
rect 11722 33488 12842 34105
rect 13010 33488 14130 34105
rect 14298 33488 16062 34105
rect 16230 33488 17350 34105
rect 17518 33488 18638 34105
rect 18806 33488 20570 34105
rect 20738 33488 21858 34105
rect 22026 33488 23790 34105
rect 23958 33488 25078 34105
rect 25246 33488 26366 34105
rect 26534 33488 28298 34105
rect 28466 33488 29586 34105
rect 29754 33488 31518 34105
rect 31686 33488 32806 34105
rect 32974 33488 34094 34105
rect 34262 33488 34848 34105
rect 20 856 34848 33488
rect 130 734 1250 856
rect 1418 734 2538 856
rect 2706 734 4470 856
rect 4638 734 5758 856
rect 5926 734 7046 856
rect 7214 734 8978 856
rect 9146 734 10266 856
rect 10434 734 12198 856
rect 12366 734 13486 856
rect 13654 734 14774 856
rect 14942 734 16706 856
rect 16874 734 17994 856
rect 18162 734 19282 856
rect 19450 734 21214 856
rect 21382 734 22502 856
rect 22670 734 24434 856
rect 24602 734 25722 856
rect 25890 734 27010 856
rect 27178 734 28942 856
rect 29110 734 30230 856
rect 30398 734 32162 856
rect 32330 734 33450 856
rect 33618 734 34738 856
<< metal3 >>
rect 0 34008 800 34128
rect 34168 33328 34968 33448
rect 0 31968 800 32088
rect 34168 31968 34968 32088
rect 0 30608 800 30728
rect 34168 30608 34968 30728
rect 0 28568 800 28688
rect 34168 28568 34968 28688
rect 0 27208 800 27328
rect 34168 27208 34968 27328
rect 0 25848 800 25968
rect 34168 25168 34968 25288
rect 0 23808 800 23928
rect 34168 23808 34968 23928
rect 0 22448 800 22568
rect 34168 22448 34968 22568
rect 0 20408 800 20528
rect 34168 20408 34968 20528
rect 0 19048 800 19168
rect 34168 19048 34968 19168
rect 0 17688 800 17808
rect 34168 17008 34968 17128
rect 0 15648 800 15768
rect 34168 15648 34968 15768
rect 0 14288 800 14408
rect 34168 14288 34968 14408
rect 0 12928 800 13048
rect 34168 12248 34968 12368
rect 0 10888 800 11008
rect 34168 10888 34968 11008
rect 0 9528 800 9648
rect 34168 9528 34968 9648
rect 0 7488 800 7608
rect 34168 7488 34968 7608
rect 0 6128 800 6248
rect 34168 6128 34968 6248
rect 0 4768 800 4888
rect 34168 4088 34968 4208
rect 0 2728 800 2848
rect 34168 2728 34968 2848
rect 0 1368 800 1488
rect 34168 1368 34968 1488
<< obsm3 >>
rect 880 33928 34168 34101
rect 800 33528 34168 33928
rect 800 33248 34088 33528
rect 800 32168 34168 33248
rect 880 31888 34088 32168
rect 800 30808 34168 31888
rect 880 30528 34088 30808
rect 800 28768 34168 30528
rect 880 28488 34088 28768
rect 800 27408 34168 28488
rect 880 27128 34088 27408
rect 800 26048 34168 27128
rect 880 25768 34168 26048
rect 800 25368 34168 25768
rect 800 25088 34088 25368
rect 800 24008 34168 25088
rect 880 23728 34088 24008
rect 800 22648 34168 23728
rect 880 22368 34088 22648
rect 800 20608 34168 22368
rect 880 20328 34088 20608
rect 800 19248 34168 20328
rect 880 18968 34088 19248
rect 800 17888 34168 18968
rect 880 17608 34168 17888
rect 800 17208 34168 17608
rect 800 16928 34088 17208
rect 800 15848 34168 16928
rect 880 15568 34088 15848
rect 800 14488 34168 15568
rect 880 14208 34088 14488
rect 800 13128 34168 14208
rect 880 12848 34168 13128
rect 800 12448 34168 12848
rect 800 12168 34088 12448
rect 800 11088 34168 12168
rect 880 10808 34088 11088
rect 800 9728 34168 10808
rect 880 9448 34088 9728
rect 800 7688 34168 9448
rect 880 7408 34088 7688
rect 800 6328 34168 7408
rect 880 6048 34088 6328
rect 800 4968 34168 6048
rect 880 4688 34168 4968
rect 800 4288 34168 4688
rect 800 4008 34088 4288
rect 800 2928 34168 4008
rect 880 2648 34088 2928
rect 800 1568 34168 2648
rect 880 1395 34088 1568
<< metal4 >>
rect 6280 2672 6600 32144
rect 6940 2672 7260 32144
rect 13640 2672 13960 32144
rect 14300 2672 14620 32144
rect 21000 2672 21320 32144
rect 21660 2672 21980 32144
rect 28360 2672 28680 32144
rect 29020 2672 29340 32144
<< obsm4 >>
rect 11099 5475 13560 31925
rect 14040 5475 14220 31925
rect 14700 5475 20920 31925
rect 21400 5475 21580 31925
rect 22060 5475 24597 31925
<< labels >>
rlabel metal3 s 0 17688 800 17808 6 clk
port 1 nsew signal input
rlabel metal3 s 34168 28568 34968 28688 6 i_start_rx
port 2 nsew signal input
rlabel metal3 s 34168 6128 34968 6248 6 i_uart_rx
port 3 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 o_uart_tx
port 4 nsew signal output
rlabel metal3 s 34168 27208 34968 27328 6 rst
port 5 nsew signal input
rlabel metal4 s 6280 2672 6600 32144 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 13640 2672 13960 32144 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 21000 2672 21320 32144 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 28360 2672 28680 32144 6 vccd1
port 6 nsew power bidirectional
rlabel metal4 s 6940 2672 7260 32144 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 14300 2672 14620 32144 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 21660 2672 21980 32144 6 vssd1
port 7 nsew ground bidirectional
rlabel metal4 s 29020 2672 29340 32144 6 vssd1
port 7 nsew ground bidirectional
rlabel metal3 s 34168 20408 34968 20528 6 wb_ack_i
port 8 nsew signal input
rlabel metal2 s 16118 33544 16174 34344 6 wb_adr_o[0]
port 9 nsew signal output
rlabel metal2 s 14186 33544 14242 34344 6 wb_adr_o[10]
port 10 nsew signal output
rlabel metal3 s 34168 12248 34968 12368 6 wb_adr_o[11]
port 11 nsew signal output
rlabel metal2 s 1950 33544 2006 34344 6 wb_adr_o[12]
port 12 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 wb_adr_o[13]
port 13 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 wb_adr_o[14]
port 14 nsew signal output
rlabel metal2 s 12254 0 12310 800 6 wb_adr_o[15]
port 15 nsew signal output
rlabel metal3 s 34168 25168 34968 25288 6 wb_adr_o[1]
port 16 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 wb_adr_o[2]
port 17 nsew signal output
rlabel metal3 s 34168 22448 34968 22568 6 wb_adr_o[3]
port 18 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wb_adr_o[4]
port 19 nsew signal output
rlabel metal2 s 32862 33544 32918 34344 6 wb_adr_o[5]
port 20 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 wb_adr_o[6]
port 21 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 wb_adr_o[7]
port 22 nsew signal output
rlabel metal2 s 23846 33544 23902 34344 6 wb_adr_o[8]
port 23 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 wb_adr_o[9]
port 24 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wb_cyc_o
port 25 nsew signal output
rlabel metal2 s 21914 33544 21970 34344 6 wb_dat_i[0]
port 26 nsew signal input
rlabel metal3 s 34168 23808 34968 23928 6 wb_dat_i[10]
port 27 nsew signal input
rlabel metal2 s 6458 33544 6514 34344 6 wb_dat_i[11]
port 28 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 wb_dat_i[12]
port 29 nsew signal input
rlabel metal3 s 34168 14288 34968 14408 6 wb_dat_i[13]
port 30 nsew signal input
rlabel metal2 s 18694 33544 18750 34344 6 wb_dat_i[14]
port 31 nsew signal input
rlabel metal3 s 34168 2728 34968 2848 6 wb_dat_i[15]
port 32 nsew signal input
rlabel metal2 s 25134 33544 25190 34344 6 wb_dat_i[16]
port 33 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 wb_dat_i[17]
port 34 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 wb_dat_i[18]
port 35 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 wb_dat_i[19]
port 36 nsew signal input
rlabel metal2 s 17406 33544 17462 34344 6 wb_dat_i[1]
port 37 nsew signal input
rlabel metal3 s 34168 33328 34968 33448 6 wb_dat_i[20]
port 38 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 wb_dat_i[21]
port 39 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wb_dat_i[22]
port 40 nsew signal input
rlabel metal3 s 34168 10888 34968 11008 6 wb_dat_i[23]
port 41 nsew signal input
rlabel metal2 s 662 33544 718 34344 6 wb_dat_i[24]
port 42 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wb_dat_i[25]
port 43 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wb_dat_i[26]
port 44 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 wb_dat_i[27]
port 45 nsew signal input
rlabel metal3 s 34168 30608 34968 30728 6 wb_dat_i[28]
port 46 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 wb_dat_i[29]
port 47 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wb_dat_i[2]
port 48 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 wb_dat_i[30]
port 49 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wb_dat_i[31]
port 50 nsew signal input
rlabel metal3 s 34168 9528 34968 9648 6 wb_dat_i[3]
port 51 nsew signal input
rlabel metal3 s 34168 4088 34968 4208 6 wb_dat_i[4]
port 52 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wb_dat_i[5]
port 53 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 wb_dat_i[6]
port 54 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wb_dat_i[7]
port 55 nsew signal input
rlabel metal2 s 9678 33544 9734 34344 6 wb_dat_i[8]
port 56 nsew signal input
rlabel metal3 s 34168 7488 34968 7608 6 wb_dat_i[9]
port 57 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 wb_dat_o[0]
port 58 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wb_dat_o[10]
port 59 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 wb_dat_o[11]
port 60 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 wb_dat_o[12]
port 61 nsew signal output
rlabel metal2 s 12898 33544 12954 34344 6 wb_dat_o[13]
port 62 nsew signal output
rlabel metal2 s 16762 0 16818 800 6 wb_dat_o[14]
port 63 nsew signal output
rlabel metal2 s 18 0 74 800 6 wb_dat_o[15]
port 64 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wb_dat_o[16]
port 65 nsew signal output
rlabel metal2 s 11610 33544 11666 34344 6 wb_dat_o[17]
port 66 nsew signal output
rlabel metal2 s 20626 33544 20682 34344 6 wb_dat_o[18]
port 67 nsew signal output
rlabel metal2 s 31574 33544 31630 34344 6 wb_dat_o[19]
port 68 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 wb_dat_o[1]
port 69 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wb_dat_o[20]
port 70 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 wb_dat_o[21]
port 71 nsew signal output
rlabel metal2 s 34150 33544 34206 34344 6 wb_dat_o[22]
port 72 nsew signal output
rlabel metal2 s 26422 33544 26478 34344 6 wb_dat_o[23]
port 73 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wb_dat_o[24]
port 74 nsew signal output
rlabel metal3 s 34168 31968 34968 32088 6 wb_dat_o[25]
port 75 nsew signal output
rlabel metal3 s 34168 1368 34968 1488 6 wb_dat_o[26]
port 76 nsew signal output
rlabel metal2 s 5170 33544 5226 34344 6 wb_dat_o[27]
port 77 nsew signal output
rlabel metal3 s 34168 17008 34968 17128 6 wb_dat_o[28]
port 78 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 wb_dat_o[29]
port 79 nsew signal output
rlabel metal2 s 10322 0 10378 800 6 wb_dat_o[2]
port 80 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 wb_dat_o[30]
port 81 nsew signal output
rlabel metal3 s 34168 19048 34968 19168 6 wb_dat_o[31]
port 82 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wb_dat_o[3]
port 83 nsew signal output
rlabel metal2 s 29642 33544 29698 34344 6 wb_dat_o[4]
port 84 nsew signal output
rlabel metal2 s 28354 33544 28410 34344 6 wb_dat_o[5]
port 85 nsew signal output
rlabel metal2 s 3882 33544 3938 34344 6 wb_dat_o[6]
port 86 nsew signal output
rlabel metal2 s 8390 33544 8446 34344 6 wb_dat_o[7]
port 87 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wb_dat_o[8]
port 88 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 wb_dat_o[9]
port 89 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 wb_stb_o
port 90 nsew signal output
rlabel metal3 s 34168 15648 34968 15768 6 wb_we_o
port 91 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 34968 34344
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3558088
string GDS_FILE /home/roliveira/Desktop/osiris_i_rtl_folder/osiris_i/openlane/uart_wbs_bridge/runs/metal/results/signoff/uart_wbs_bridge.magic.gds
string GDS_START 683116
<< end >>

