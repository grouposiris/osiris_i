magic
tech sky130A
magscale 1 2
timestamp 1731048028
<< viali >>
rect 4353 34085 4387 34119
rect 14105 34085 14139 34119
rect 21097 34085 21131 34119
rect 28825 34085 28859 34119
rect 3065 34017 3099 34051
rect 5089 34017 5123 34051
rect 6009 34017 6043 34051
rect 8033 34017 8067 34051
rect 9045 34017 9079 34051
rect 10609 34017 10643 34051
rect 12541 34017 12575 34051
rect 13369 34017 13403 34051
rect 15577 34017 15611 34051
rect 15761 34017 15795 34051
rect 18429 34017 18463 34051
rect 22109 34017 22143 34051
rect 22661 34017 22695 34051
rect 24133 34017 24167 34051
rect 26065 34017 26099 34051
rect 30021 34017 30055 34051
rect 31217 34017 31251 34051
rect 6377 33949 6411 33983
rect 9689 33949 9723 33983
rect 10885 33949 10919 33983
rect 11713 33949 11747 33983
rect 15209 33949 15243 33983
rect 18797 33949 18831 33983
rect 24409 33949 24443 33983
rect 26525 33949 26559 33983
rect 31769 33949 31803 33983
rect 3249 33813 3283 33847
rect 8217 33813 8251 33847
rect 12265 33813 12299 33847
rect 12449 33813 12483 33847
rect 14657 33813 14691 33847
rect 15393 33813 15427 33847
rect 15945 33813 15979 33847
rect 22845 33813 22879 33847
rect 3525 33473 3559 33507
rect 5917 33473 5951 33507
rect 12725 33473 12759 33507
rect 13829 33473 13863 33507
rect 26985 33473 27019 33507
rect 30297 33473 30331 33507
rect 31769 33473 31803 33507
rect 4721 33405 4755 33439
rect 5457 33405 5491 33439
rect 8677 33405 8711 33439
rect 10793 33405 10827 33439
rect 13001 33405 13035 33439
rect 13553 33405 13587 33439
rect 15577 33405 15611 33439
rect 18797 33405 18831 33439
rect 18889 33405 18923 33439
rect 21373 33405 21407 33439
rect 26525 33405 26559 33439
rect 31033 33405 31067 33439
rect 31401 33405 31435 33439
rect 8953 33337 8987 33371
rect 10701 33337 10735 33371
rect 13093 33337 13127 33371
rect 13277 33337 13311 33371
rect 15485 33337 15519 33371
rect 5089 33269 5123 33303
rect 10425 33269 10459 33303
rect 11253 33269 11287 33303
rect 15301 33269 15335 33303
rect 18705 33269 18739 33303
rect 19073 33269 19107 33303
rect 21557 33269 21591 33303
rect 9045 33065 9079 33099
rect 11621 33065 11655 33099
rect 14013 33065 14047 33099
rect 3249 32997 3283 33031
rect 4721 32997 4755 33031
rect 10149 32997 10183 33031
rect 11345 32997 11379 33031
rect 11897 32997 11931 33031
rect 15761 32997 15795 33031
rect 30297 32997 30331 33031
rect 4445 32929 4479 32963
rect 5733 32929 5767 32963
rect 6929 32929 6963 32963
rect 9965 32929 9999 32963
rect 10057 32929 10091 32963
rect 10287 32929 10321 32963
rect 11161 32929 11195 32963
rect 11253 32929 11287 32963
rect 11437 32929 11471 32963
rect 11822 32919 11856 32953
rect 11989 32929 12023 32963
rect 12127 32929 12161 32963
rect 12449 32929 12483 32963
rect 13369 32929 13403 32963
rect 13553 32929 13587 32963
rect 13645 32929 13679 32963
rect 14010 32929 14044 32963
rect 14565 32929 14599 32963
rect 14749 32929 14783 32963
rect 15485 32929 15519 32963
rect 15577 32929 15611 32963
rect 15853 32929 15887 32963
rect 19073 32929 19107 32963
rect 29285 32929 29319 32963
rect 32137 32929 32171 32963
rect 32321 32929 32355 32963
rect 6193 32861 6227 32895
rect 9689 32861 9723 32895
rect 9781 32861 9815 32895
rect 10425 32861 10459 32895
rect 12265 32861 12299 32895
rect 13001 32861 13035 32895
rect 14473 32861 14507 32895
rect 14657 32861 14691 32895
rect 16129 32861 16163 32895
rect 18889 32861 18923 32895
rect 19349 32861 19383 32895
rect 31677 32861 31711 32895
rect 32781 32861 32815 32895
rect 13185 32793 13219 32827
rect 13829 32793 13863 32827
rect 15577 32793 15611 32827
rect 18061 32793 18095 32827
rect 7297 32725 7331 32759
rect 10977 32725 11011 32759
rect 14381 32725 14415 32759
rect 14841 32725 14875 32759
rect 16773 32725 16807 32759
rect 18337 32725 18371 32759
rect 10609 32521 10643 32555
rect 12449 32521 12483 32555
rect 13369 32521 13403 32555
rect 14105 32521 14139 32555
rect 14657 32521 14691 32555
rect 17245 32521 17279 32555
rect 5549 32453 5583 32487
rect 13921 32453 13955 32487
rect 15393 32453 15427 32487
rect 23949 32453 23983 32487
rect 3249 32385 3283 32419
rect 5273 32385 5307 32419
rect 6009 32385 6043 32419
rect 6193 32385 6227 32419
rect 6561 32385 6595 32419
rect 12265 32385 12299 32419
rect 17509 32385 17543 32419
rect 17601 32385 17635 32419
rect 17877 32385 17911 32419
rect 23121 32385 23155 32419
rect 23305 32385 23339 32419
rect 24593 32385 24627 32419
rect 28549 32385 28583 32419
rect 30297 32385 30331 32419
rect 33793 32385 33827 32419
rect 4445 32317 4479 32351
rect 8953 32317 8987 32351
rect 9321 32317 9355 32351
rect 10977 32317 11011 32351
rect 12081 32317 12115 32351
rect 12357 32317 12391 32351
rect 12541 32317 12575 32351
rect 13277 32317 13311 32351
rect 13369 32317 13403 32351
rect 14381 32317 14415 32351
rect 14657 32317 14691 32351
rect 14841 32317 14875 32351
rect 15577 32317 15611 32351
rect 19625 32317 19659 32351
rect 19993 32317 20027 32351
rect 24961 32317 24995 32351
rect 32781 32317 32815 32351
rect 10793 32249 10827 32283
rect 12909 32249 12943 32283
rect 14289 32249 14323 32283
rect 23489 32249 23523 32283
rect 28733 32249 28767 32283
rect 29653 32249 29687 32283
rect 4629 32181 4663 32215
rect 5917 32181 5951 32215
rect 8401 32181 8435 32215
rect 9229 32181 9263 32215
rect 11897 32181 11931 32215
rect 13553 32181 13587 32215
rect 14105 32181 14139 32215
rect 15761 32181 15795 32215
rect 19349 32181 19383 32215
rect 23581 32181 23615 32215
rect 24041 32181 24075 32215
rect 24869 32181 24903 32215
rect 28273 32181 28307 32215
rect 28825 32181 28859 32215
rect 29193 32181 29227 32215
rect 9781 31977 9815 32011
rect 10149 31977 10183 32011
rect 18337 31977 18371 32011
rect 19441 31977 19475 32011
rect 25237 31977 25271 32011
rect 30389 31977 30423 32011
rect 5181 31909 5215 31943
rect 6837 31909 6871 31943
rect 8309 31909 8343 31943
rect 11095 31909 11129 31943
rect 11621 31909 11655 31943
rect 14717 31909 14751 31943
rect 14933 31909 14967 31943
rect 15209 31909 15243 31943
rect 15393 31909 15427 31943
rect 18797 31909 18831 31943
rect 23765 31909 23799 31943
rect 28917 31909 28951 31943
rect 33425 31909 33459 31943
rect 4445 31841 4479 31875
rect 4905 31841 4939 31875
rect 6929 31841 6963 31875
rect 8033 31841 8067 31875
rect 10793 31841 10827 31875
rect 10885 31841 10919 31875
rect 10977 31841 11011 31875
rect 11345 31841 11379 31875
rect 11437 31841 11471 31875
rect 15301 31841 15335 31875
rect 18705 31841 18739 31875
rect 27629 31841 27663 31875
rect 27905 31841 27939 31875
rect 32229 31841 32263 31875
rect 3249 31773 3283 31807
rect 6653 31773 6687 31807
rect 11253 31773 11287 31807
rect 16957 31773 16991 31807
rect 17785 31773 17819 31807
rect 18981 31773 19015 31807
rect 23489 31773 23523 31807
rect 28641 31773 28675 31807
rect 30665 31773 30699 31807
rect 31861 31773 31895 31807
rect 32137 31773 32171 31807
rect 14565 31705 14599 31739
rect 10609 31637 10643 31671
rect 11529 31637 11563 31671
rect 14749 31637 14783 31671
rect 17233 31637 17267 31671
rect 26985 31637 27019 31671
rect 27813 31637 27847 31671
rect 4813 31433 4847 31467
rect 15301 31433 15335 31467
rect 15485 31433 15519 31467
rect 18337 31433 18371 31467
rect 31309 31433 31343 31467
rect 3065 31297 3099 31331
rect 5917 31297 5951 31331
rect 10425 31297 10459 31331
rect 16589 31297 16623 31331
rect 16865 31297 16899 31331
rect 18797 31297 18831 31331
rect 22293 31297 22327 31331
rect 26525 31297 26559 31331
rect 26801 31297 26835 31331
rect 28273 31297 28307 31331
rect 30021 31297 30055 31331
rect 33793 31297 33827 31331
rect 5089 31229 5123 31263
rect 5549 31229 5583 31263
rect 7757 31229 7791 31263
rect 11161 31229 11195 31263
rect 12173 31229 12207 31263
rect 15393 31229 15427 31263
rect 16497 31229 16531 31263
rect 18429 31229 18463 31263
rect 28365 31229 28399 31263
rect 30757 31229 30791 31263
rect 31401 31229 31435 31263
rect 32505 31229 32539 31263
rect 32781 31229 32815 31263
rect 3341 31161 3375 31195
rect 4997 31161 5031 31195
rect 11897 31161 11931 31195
rect 22569 31161 22603 31195
rect 29193 31161 29227 31195
rect 31769 31161 31803 31195
rect 9045 31093 9079 31127
rect 9781 31093 9815 31127
rect 11345 31093 11379 31127
rect 12081 31093 12115 31127
rect 12265 31093 12299 31127
rect 12449 31093 12483 31127
rect 16313 31093 16347 31127
rect 24041 31093 24075 31127
rect 29469 31093 29503 31127
rect 30205 31093 30239 31127
rect 31861 31093 31895 31127
rect 6377 30889 6411 30923
rect 8401 30889 8435 30923
rect 11713 30889 11747 30923
rect 16589 30889 16623 30923
rect 17325 30889 17359 30923
rect 23489 30889 23523 30923
rect 27629 30889 27663 30923
rect 33609 30889 33643 30923
rect 3985 30821 4019 30855
rect 4721 30821 4755 30855
rect 8861 30821 8895 30855
rect 9505 30821 9539 30855
rect 11161 30821 11195 30855
rect 16773 30821 16807 30855
rect 29285 30821 29319 30855
rect 31677 30821 31711 30855
rect 32137 30821 32171 30855
rect 33885 30821 33919 30855
rect 8309 30753 8343 30787
rect 8769 30753 8803 30787
rect 9229 30753 9263 30787
rect 11069 30753 11103 30787
rect 11529 30753 11563 30787
rect 11805 30753 11839 30787
rect 12633 30753 12667 30787
rect 13369 30753 13403 30787
rect 14841 30753 14875 30787
rect 16865 30753 16899 30787
rect 17693 30753 17727 30787
rect 17785 30753 17819 30787
rect 18521 30753 18555 30787
rect 24777 30753 24811 30787
rect 27537 30753 27571 30787
rect 29009 30753 29043 30787
rect 31401 30753 31435 30787
rect 31769 30753 31803 30787
rect 33793 30753 33827 30787
rect 5273 30685 5307 30719
rect 9045 30685 9079 30719
rect 12725 30685 12759 30719
rect 12817 30685 12851 30719
rect 15117 30685 15151 30719
rect 17877 30685 17911 30719
rect 18429 30685 18463 30719
rect 19717 30685 19751 30719
rect 24041 30685 24075 30719
rect 25513 30685 25547 30719
rect 27721 30685 27755 30719
rect 30757 30685 30791 30719
rect 31861 30685 31895 30719
rect 11345 30617 11379 30651
rect 4997 30549 5031 30583
rect 5825 30549 5859 30583
rect 8217 30549 8251 30583
rect 10977 30549 11011 30583
rect 12265 30549 12299 30583
rect 13277 30549 13311 30583
rect 17141 30549 17175 30583
rect 19165 30549 19199 30583
rect 24225 30549 24259 30583
rect 24961 30549 24995 30583
rect 26985 30549 27019 30583
rect 27169 30549 27203 30583
rect 28917 30549 28951 30583
rect 30849 30549 30883 30583
rect 3801 30345 3835 30379
rect 5457 30345 5491 30379
rect 14933 30345 14967 30379
rect 23581 30345 23615 30379
rect 32965 30345 32999 30379
rect 3709 30277 3743 30311
rect 23765 30277 23799 30311
rect 30205 30277 30239 30311
rect 4445 30209 4479 30243
rect 5273 30209 5307 30243
rect 6101 30209 6135 30243
rect 7941 30209 7975 30243
rect 11989 30209 12023 30243
rect 12265 30209 12299 30243
rect 23029 30209 23063 30243
rect 23121 30209 23155 30243
rect 24041 30209 24075 30243
rect 24317 30209 24351 30243
rect 29561 30209 29595 30243
rect 29745 30209 29779 30243
rect 4169 30141 4203 30175
rect 5825 30141 5859 30175
rect 6929 30141 6963 30175
rect 7205 30141 7239 30175
rect 11161 30141 11195 30175
rect 15577 30141 15611 30175
rect 15761 30141 15795 30175
rect 15945 30141 15979 30175
rect 16221 30141 16255 30175
rect 16865 30141 16899 30175
rect 23857 30141 23891 30175
rect 26249 30141 26283 30175
rect 26893 30141 26927 30175
rect 28549 30141 28583 30175
rect 29377 30141 29411 30175
rect 30481 30141 30515 30175
rect 31217 30141 31251 30175
rect 33701 30141 33735 30175
rect 33977 30141 34011 30175
rect 3157 30073 3191 30107
rect 8217 30073 8251 30107
rect 16129 30073 16163 30107
rect 26157 30073 26191 30107
rect 31033 30073 31067 30107
rect 31493 30073 31527 30107
rect 3249 30005 3283 30039
rect 4261 30005 4295 30039
rect 4629 30005 4663 30039
rect 5917 30005 5951 30039
rect 6285 30005 6319 30039
rect 7113 30005 7147 30039
rect 9689 30005 9723 30039
rect 10149 30005 10183 30039
rect 10609 30005 10643 30039
rect 13737 30005 13771 30039
rect 16313 30005 16347 30039
rect 23213 30005 23247 30039
rect 25789 30005 25823 30039
rect 26985 30005 27019 30039
rect 27445 30005 27479 30039
rect 27721 30005 27755 30039
rect 27905 30005 27939 30039
rect 28733 30005 28767 30039
rect 29837 30005 29871 30039
rect 8861 29801 8895 29835
rect 9781 29801 9815 29835
rect 12173 29801 12207 29835
rect 13185 29801 13219 29835
rect 14105 29801 14139 29835
rect 14473 29801 14507 29835
rect 15485 29801 15519 29835
rect 16037 29801 16071 29835
rect 16497 29801 16531 29835
rect 24869 29801 24903 29835
rect 25329 29801 25363 29835
rect 27721 29801 27755 29835
rect 28641 29801 28675 29835
rect 31125 29801 31159 29835
rect 32689 29801 32723 29835
rect 33149 29801 33183 29835
rect 6009 29733 6043 29767
rect 11897 29733 11931 29767
rect 14197 29733 14231 29767
rect 18337 29733 18371 29767
rect 29285 29733 29319 29767
rect 4445 29665 4479 29699
rect 6285 29665 6319 29699
rect 8769 29665 8803 29699
rect 10425 29665 10459 29699
rect 10609 29665 10643 29699
rect 10701 29665 10735 29699
rect 11989 29665 12023 29699
rect 12081 29665 12115 29699
rect 12265 29665 12299 29699
rect 12357 29665 12391 29699
rect 13369 29665 13403 29699
rect 13829 29665 13863 29699
rect 14289 29665 14323 29699
rect 15209 29665 15243 29699
rect 15393 29665 15427 29699
rect 15577 29665 15611 29699
rect 16129 29665 16163 29699
rect 17601 29665 17635 29699
rect 24961 29665 24995 29699
rect 28825 29665 28859 29699
rect 28917 29665 28951 29699
rect 29009 29665 29043 29699
rect 29193 29665 29227 29699
rect 31493 29665 31527 29699
rect 31585 29665 31619 29699
rect 31953 29665 31987 29699
rect 32597 29665 32631 29699
rect 33057 29665 33091 29699
rect 4077 29597 4111 29631
rect 4537 29597 4571 29631
rect 6929 29597 6963 29631
rect 9873 29597 9907 29631
rect 10057 29597 10091 29631
rect 13001 29597 13035 29631
rect 13461 29597 13495 29631
rect 15945 29597 15979 29631
rect 18981 29597 19015 29631
rect 24777 29597 24811 29631
rect 25881 29597 25915 29631
rect 26157 29597 26191 29631
rect 27629 29597 27663 29631
rect 28273 29597 28307 29631
rect 31677 29597 31711 29631
rect 33241 29597 33275 29631
rect 9413 29529 9447 29563
rect 13921 29529 13955 29563
rect 17417 29529 17451 29563
rect 24133 29529 24167 29563
rect 6377 29461 6411 29495
rect 10241 29461 10275 29495
rect 13369 29461 13403 29495
rect 15025 29461 15059 29495
rect 23673 29461 23707 29495
rect 24501 29461 24535 29495
rect 30573 29461 30607 29495
rect 3065 29257 3099 29291
rect 6193 29257 6227 29291
rect 11989 29257 12023 29291
rect 14105 29257 14139 29291
rect 15117 29257 15151 29291
rect 17601 29257 17635 29291
rect 19441 29257 19475 29291
rect 23765 29257 23799 29291
rect 26617 29257 26651 29291
rect 29469 29257 29503 29291
rect 32413 29257 32447 29291
rect 6469 29189 6503 29223
rect 12265 29189 12299 29223
rect 13645 29189 13679 29223
rect 4537 29121 4571 29155
rect 5549 29121 5583 29155
rect 5733 29121 5767 29155
rect 7297 29121 7331 29155
rect 9045 29121 9079 29155
rect 12633 29121 12667 29155
rect 13921 29121 13955 29155
rect 14473 29121 14507 29155
rect 14841 29121 14875 29155
rect 14958 29121 14992 29155
rect 15853 29121 15887 29155
rect 16129 29121 16163 29155
rect 21281 29121 21315 29155
rect 23029 29121 23063 29155
rect 23121 29121 23155 29155
rect 24409 29121 24443 29155
rect 27721 29121 27755 29155
rect 27997 29121 28031 29155
rect 29561 29121 29595 29155
rect 4813 29053 4847 29087
rect 5089 29053 5123 29087
rect 9505 29053 9539 29087
rect 11621 29053 11655 29087
rect 11713 29053 11747 29087
rect 12081 29053 12115 29087
rect 13829 29053 13863 29087
rect 14749 29053 14783 29087
rect 17693 29053 17727 29087
rect 19717 29053 19751 29087
rect 23857 29053 23891 29087
rect 24777 29053 24811 29087
rect 27261 29053 27295 29087
rect 30941 29053 30975 29087
rect 31861 29053 31895 29087
rect 32045 29053 32079 29087
rect 32505 29053 32539 29087
rect 32597 29053 32631 29087
rect 5825 28985 5859 29019
rect 7573 28985 7607 29019
rect 10609 28985 10643 29019
rect 14289 28985 14323 29019
rect 17969 28985 18003 29019
rect 19625 28985 19659 29019
rect 21557 28985 21591 29019
rect 30297 28985 30331 29019
rect 33793 28985 33827 29019
rect 4997 28917 5031 28951
rect 9689 28917 9723 28951
rect 10793 28917 10827 28951
rect 10885 28917 10919 28951
rect 10977 28917 11011 28951
rect 11161 28917 11195 28951
rect 13277 28917 13311 28951
rect 24685 28917 24719 28951
rect 26433 28917 26467 28951
rect 27537 28917 27571 28951
rect 30205 28917 30239 28951
rect 31309 28917 31343 28951
rect 32137 28917 32171 28951
rect 8309 28713 8343 28747
rect 8493 28713 8527 28747
rect 10701 28713 10735 28747
rect 14473 28713 14507 28747
rect 15025 28713 15059 28747
rect 16129 28713 16163 28747
rect 17141 28713 17175 28747
rect 18337 28713 18371 28747
rect 21557 28713 21591 28747
rect 23029 28713 23063 28747
rect 27445 28713 27479 28747
rect 28825 28713 28859 28747
rect 30941 28713 30975 28747
rect 10333 28645 10367 28679
rect 10451 28645 10485 28679
rect 12357 28645 12391 28679
rect 15393 28645 15427 28679
rect 16497 28645 16531 28679
rect 18153 28645 18187 28679
rect 19349 28645 19383 28679
rect 19441 28645 19475 28679
rect 22569 28645 22603 28679
rect 23489 28645 23523 28679
rect 27721 28645 27755 28679
rect 31309 28645 31343 28679
rect 3249 28577 3283 28611
rect 4445 28577 4479 28611
rect 5089 28577 5123 28611
rect 7757 28577 7791 28611
rect 7849 28577 7883 28611
rect 8217 28577 8251 28611
rect 9137 28577 9171 28611
rect 9965 28577 9999 28611
rect 10149 28577 10183 28611
rect 10241 28577 10275 28611
rect 10609 28577 10643 28611
rect 10701 28577 10735 28611
rect 10793 28577 10827 28611
rect 10977 28577 11011 28611
rect 11437 28577 11471 28611
rect 11529 28577 11563 28611
rect 11897 28577 11931 28611
rect 12633 28577 12667 28611
rect 14657 28577 14691 28611
rect 14749 28577 14783 28611
rect 14933 28577 14967 28611
rect 15117 28577 15151 28611
rect 16313 28577 16347 28611
rect 16405 28577 16439 28611
rect 17233 28577 17267 28611
rect 19257 28577 19291 28611
rect 19625 28577 19659 28611
rect 22477 28577 22511 28611
rect 22661 28577 22695 28611
rect 22845 28577 22879 28611
rect 23121 28577 23155 28611
rect 27629 28577 27663 28611
rect 27813 28577 27847 28611
rect 27997 28577 28031 28611
rect 28733 28577 28767 28611
rect 33793 28577 33827 28611
rect 5365 28509 5399 28543
rect 6837 28509 6871 28543
rect 6929 28509 6963 28543
rect 7573 28509 7607 28543
rect 9873 28509 9907 28543
rect 12449 28509 12483 28543
rect 13737 28509 13771 28543
rect 15301 28509 15335 28543
rect 16037 28509 16071 28543
rect 18981 28509 19015 28543
rect 22201 28509 22235 28543
rect 25237 28509 25271 28543
rect 25513 28509 25547 28543
rect 25605 28509 25639 28543
rect 25881 28509 25915 28543
rect 29193 28509 29227 28543
rect 29469 28509 29503 28543
rect 31033 28509 31067 28543
rect 33425 28509 33459 28543
rect 12081 28441 12115 28475
rect 12817 28441 12851 28475
rect 16681 28441 16715 28475
rect 19073 28441 19107 28475
rect 22293 28441 22327 28475
rect 27353 28441 27387 28475
rect 9229 28373 9263 28407
rect 11805 28373 11839 28407
rect 12633 28373 12667 28407
rect 13185 28373 13219 28407
rect 28273 28373 28307 28407
rect 32781 28373 32815 28407
rect 32873 28373 32907 28407
rect 33885 28373 33919 28407
rect 5273 28169 5307 28203
rect 7744 28169 7778 28203
rect 10609 28169 10643 28203
rect 12081 28169 12115 28203
rect 13001 28169 13035 28203
rect 13553 28169 13587 28203
rect 13645 28169 13679 28203
rect 14105 28169 14139 28203
rect 17509 28169 17543 28203
rect 24225 28169 24259 28203
rect 25421 28169 25455 28203
rect 26065 28169 26099 28203
rect 26801 28169 26835 28203
rect 29193 28169 29227 28203
rect 29929 28169 29963 28203
rect 31217 28169 31251 28203
rect 9965 28101 9999 28135
rect 10885 28101 10919 28135
rect 9229 28033 9263 28067
rect 10977 28033 11011 28067
rect 12909 28033 12943 28067
rect 13369 28033 13403 28067
rect 13921 28033 13955 28067
rect 14381 28033 14415 28067
rect 15761 28033 15795 28067
rect 27169 28033 27203 28067
rect 29101 28033 29135 28067
rect 29745 28033 29779 28067
rect 31769 28033 31803 28067
rect 32413 28033 32447 28067
rect 3985 27965 4019 27999
rect 4721 27965 4755 27999
rect 5641 27965 5675 27999
rect 7481 27965 7515 27999
rect 9781 27965 9815 27999
rect 10793 27965 10827 27999
rect 11069 27965 11103 27999
rect 11253 27965 11287 27999
rect 11437 27965 11471 27999
rect 12725 27965 12759 27999
rect 13277 27965 13311 27999
rect 13553 27965 13587 27999
rect 13829 27965 13863 27999
rect 14565 27965 14599 27999
rect 19625 27965 19659 27999
rect 21097 27965 21131 27999
rect 24777 27965 24811 27999
rect 26249 27965 26283 27999
rect 26433 27965 26467 27999
rect 26617 27965 26651 27999
rect 26709 27965 26743 27999
rect 27353 27965 27387 27999
rect 30481 27965 30515 27999
rect 30849 27965 30883 27999
rect 32137 27965 32171 27999
rect 7389 27897 7423 27931
rect 13001 27897 13035 27931
rect 14105 27897 14139 27931
rect 16037 27897 16071 27931
rect 22937 27897 22971 27931
rect 26341 27897 26375 27931
rect 27629 27897 27663 27931
rect 31585 27897 31619 27931
rect 31677 27897 31711 27931
rect 4537 27829 4571 27863
rect 12541 27829 12575 27863
rect 13093 27829 13127 27863
rect 14657 27829 14691 27863
rect 15025 27829 15059 27863
rect 17785 27829 17819 27863
rect 18981 27829 19015 27863
rect 21005 27829 21039 27863
rect 21925 27829 21959 27863
rect 22293 27829 22327 27863
rect 22753 27829 22787 27863
rect 25697 27829 25731 27863
rect 30757 27829 30791 27863
rect 33885 27829 33919 27863
rect 6745 27625 6779 27659
rect 8401 27625 8435 27659
rect 11069 27625 11103 27659
rect 11529 27625 11563 27659
rect 14381 27625 14415 27659
rect 16221 27625 16255 27659
rect 16773 27625 16807 27659
rect 17785 27625 17819 27659
rect 18153 27625 18187 27659
rect 20085 27625 20119 27659
rect 28181 27625 28215 27659
rect 28733 27625 28767 27659
rect 32505 27625 32539 27659
rect 33149 27625 33183 27659
rect 4537 27557 4571 27591
rect 7021 27557 7055 27591
rect 11437 27557 11471 27591
rect 12449 27557 12483 27591
rect 14013 27557 14047 27591
rect 14213 27557 14247 27591
rect 15393 27557 15427 27591
rect 17233 27557 17267 27591
rect 17693 27557 17727 27591
rect 18613 27557 18647 27591
rect 22937 27557 22971 27591
rect 23765 27557 23799 27591
rect 23857 27557 23891 27591
rect 25053 27557 25087 27591
rect 27629 27557 27663 27591
rect 29193 27557 29227 27591
rect 31309 27557 31343 27591
rect 33057 27557 33091 27591
rect 4813 27489 4847 27523
rect 5089 27489 5123 27523
rect 6929 27489 6963 27523
rect 7113 27489 7147 27523
rect 7297 27489 7331 27523
rect 8309 27489 8343 27523
rect 9505 27489 9539 27523
rect 10885 27489 10919 27523
rect 11345 27489 11379 27523
rect 11805 27489 11839 27523
rect 12081 27489 12115 27523
rect 12541 27489 12575 27523
rect 13461 27489 13495 27523
rect 13645 27489 13679 27523
rect 15209 27489 15243 27523
rect 16129 27489 16163 27523
rect 16681 27489 16715 27523
rect 23121 27489 23155 27523
rect 24961 27489 24995 27523
rect 26525 27489 26559 27523
rect 27537 27489 27571 27523
rect 27721 27489 27755 27523
rect 27905 27489 27939 27523
rect 28825 27489 28859 27523
rect 28917 27489 28951 27523
rect 29101 27489 29135 27523
rect 29285 27489 29319 27523
rect 31217 27489 31251 27523
rect 31861 27489 31895 27523
rect 33977 27489 34011 27523
rect 4997 27421 5031 27455
rect 5273 27421 5307 27455
rect 6009 27421 6043 27455
rect 10701 27421 10735 27455
rect 12265 27421 12299 27455
rect 13553 27421 13587 27455
rect 15945 27421 15979 27455
rect 17509 27421 17543 27455
rect 18337 27421 18371 27455
rect 21741 27421 21775 27455
rect 22017 27421 22051 27455
rect 23581 27421 23615 27455
rect 24317 27421 24351 27455
rect 25605 27421 25639 27455
rect 26341 27421 26375 27455
rect 29561 27421 29595 27455
rect 30113 27421 30147 27455
rect 30573 27421 30607 27455
rect 31953 27421 31987 27455
rect 32045 27421 32079 27455
rect 33241 27421 33275 27455
rect 24225 27353 24259 27387
rect 27353 27353 27387 27387
rect 29469 27353 29503 27387
rect 32689 27353 32723 27387
rect 3065 27285 3099 27319
rect 5825 27285 5859 27319
rect 6653 27285 6687 27319
rect 7665 27285 7699 27319
rect 9597 27285 9631 27319
rect 11897 27285 11931 27319
rect 14197 27285 14231 27319
rect 14657 27285 14691 27319
rect 20269 27285 20303 27319
rect 23213 27285 23247 27319
rect 25789 27285 25823 27319
rect 26709 27285 26743 27319
rect 27077 27285 27111 27319
rect 31125 27285 31159 27319
rect 31493 27285 31527 27319
rect 33793 27285 33827 27319
rect 3985 27081 4019 27115
rect 5457 27081 5491 27115
rect 6929 27081 6963 27115
rect 7849 27081 7883 27115
rect 10333 27081 10367 27115
rect 13829 27081 13863 27115
rect 14013 27081 14047 27115
rect 15853 27081 15887 27115
rect 18613 27081 18647 27115
rect 20913 27081 20947 27115
rect 22832 27081 22866 27115
rect 24317 27081 24351 27115
rect 24961 27081 24995 27115
rect 27813 27081 27847 27115
rect 32965 27081 32999 27115
rect 33517 27081 33551 27115
rect 11161 27013 11195 27047
rect 15209 27013 15243 27047
rect 28365 27013 28399 27047
rect 31033 27013 31067 27047
rect 4445 26945 4479 26979
rect 4537 26945 4571 26979
rect 5917 26945 5951 26979
rect 6009 26945 6043 26979
rect 11253 26945 11287 26979
rect 13277 26945 13311 26979
rect 14381 26945 14415 26979
rect 15025 26945 15059 26979
rect 17325 26945 17359 26979
rect 17601 26945 17635 26979
rect 22569 26945 22603 26979
rect 26065 26945 26099 26979
rect 29101 26945 29135 26979
rect 29285 26945 29319 26979
rect 31217 26945 31251 26979
rect 3065 26877 3099 26911
rect 3893 26877 3927 26911
rect 5825 26877 5859 26911
rect 6285 26877 6319 26911
rect 7205 26877 7239 26911
rect 8585 26877 8619 26911
rect 10734 26877 10768 26911
rect 11437 26877 11471 26911
rect 11529 26877 11563 26911
rect 11713 26877 11747 26911
rect 12541 26877 12575 26911
rect 14289 26877 14323 26911
rect 14565 26877 14599 26911
rect 14933 26877 14967 26911
rect 15485 26877 15519 26911
rect 15577 26877 15611 26911
rect 18705 26877 18739 26911
rect 21097 26877 21131 26911
rect 21189 26877 21223 26911
rect 21465 26877 21499 26911
rect 24409 26877 24443 26911
rect 24685 26877 24719 26911
rect 24777 26877 24811 26911
rect 25697 26877 25731 26911
rect 27905 26877 27939 26911
rect 28641 26877 28675 26911
rect 33241 26877 33275 26911
rect 13875 26843 13909 26877
rect 4353 26809 4387 26843
rect 8861 26809 8895 26843
rect 13645 26809 13679 26843
rect 14657 26809 14691 26843
rect 15301 26809 15335 26843
rect 21281 26809 21315 26843
rect 24593 26809 24627 26843
rect 26341 26809 26375 26843
rect 28733 26809 28767 26843
rect 29561 26809 29595 26843
rect 31493 26809 31527 26843
rect 33149 26809 33183 26843
rect 3249 26741 3283 26775
rect 5181 26741 5215 26775
rect 7113 26741 7147 26775
rect 7481 26741 7515 26775
rect 10609 26741 10643 26775
rect 10793 26741 10827 26775
rect 11897 26741 11931 26775
rect 11989 26741 12023 26775
rect 12725 26741 12759 26775
rect 15399 26741 15433 26775
rect 20729 26741 20763 26775
rect 22477 26741 22511 26775
rect 25145 26741 25179 26775
rect 28089 26741 28123 26775
rect 33885 26741 33919 26775
rect 4537 26537 4571 26571
rect 7113 26537 7147 26571
rect 9321 26537 9355 26571
rect 10701 26537 10735 26571
rect 12449 26537 12483 26571
rect 13829 26537 13863 26571
rect 15393 26537 15427 26571
rect 16497 26537 16531 26571
rect 17509 26537 17543 26571
rect 22937 26537 22971 26571
rect 26893 26537 26927 26571
rect 27169 26537 27203 26571
rect 29561 26537 29595 26571
rect 31493 26537 31527 26571
rect 6009 26469 6043 26503
rect 12357 26469 12391 26503
rect 12909 26469 12943 26503
rect 20913 26469 20947 26503
rect 24133 26469 24167 26503
rect 24777 26469 24811 26503
rect 4261 26401 4295 26435
rect 6285 26401 6319 26435
rect 10885 26401 10919 26435
rect 12817 26401 12851 26435
rect 13001 26401 13035 26435
rect 13645 26401 13679 26435
rect 14105 26401 14139 26435
rect 14565 26401 14599 26435
rect 14749 26401 14783 26435
rect 15577 26401 15611 26435
rect 16589 26401 16623 26435
rect 18981 26401 19015 26435
rect 21005 26401 21039 26435
rect 22201 26401 22235 26435
rect 24869 26401 24903 26435
rect 26801 26401 26835 26435
rect 27077 26401 27111 26435
rect 27261 26401 27295 26435
rect 28089 26401 28123 26435
rect 28365 26401 28399 26435
rect 28457 26401 28491 26435
rect 29929 26401 29963 26435
rect 30389 26401 30423 26435
rect 32045 26401 32079 26435
rect 32229 26401 32263 26435
rect 3249 26333 3283 26367
rect 6929 26333 6963 26367
rect 7665 26333 7699 26367
rect 9873 26333 9907 26367
rect 11345 26333 11379 26367
rect 12541 26333 12575 26367
rect 18153 26333 18187 26367
rect 19257 26333 19291 26367
rect 23489 26333 23523 26367
rect 24593 26333 24627 26367
rect 25881 26333 25915 26367
rect 26617 26333 26651 26367
rect 27997 26333 28031 26367
rect 29193 26333 29227 26367
rect 30021 26333 30055 26367
rect 30205 26333 30239 26367
rect 30941 26333 30975 26367
rect 33057 26333 33091 26367
rect 11897 26265 11931 26299
rect 11989 26265 12023 26299
rect 17417 26265 17451 26299
rect 20729 26265 20763 26299
rect 23305 26265 23339 26299
rect 25237 26265 25271 26299
rect 27813 26265 27847 26299
rect 6377 26197 6411 26231
rect 14197 26197 14231 26231
rect 14749 26197 14783 26231
rect 15853 26197 15887 26231
rect 17049 26197 17083 26231
rect 21557 26197 21591 26231
rect 25329 26197 25363 26231
rect 26065 26197 26099 26231
rect 27537 26197 27571 26231
rect 28641 26197 28675 26231
rect 7481 25993 7515 26027
rect 9597 25993 9631 26027
rect 13645 25993 13679 26027
rect 19257 25993 19291 26027
rect 25881 25993 25915 26027
rect 26065 25993 26099 26027
rect 27077 25993 27111 26027
rect 29377 25993 29411 26027
rect 18337 25925 18371 25959
rect 27353 25925 27387 25959
rect 6009 25857 6043 25891
rect 11713 25857 11747 25891
rect 17509 25857 17543 25891
rect 21557 25857 21591 25891
rect 23029 25857 23063 25891
rect 23857 25857 23891 25891
rect 24133 25857 24167 25891
rect 24409 25857 24443 25891
rect 27629 25857 27663 25891
rect 29653 25857 29687 25891
rect 3985 25789 4019 25823
rect 5733 25789 5767 25823
rect 7757 25789 7791 25823
rect 9873 25789 9907 25823
rect 10149 25789 10183 25823
rect 10701 25789 10735 25823
rect 10977 25789 11011 25823
rect 13553 25789 13587 25823
rect 13829 25789 13863 25823
rect 13921 25789 13955 25823
rect 14105 25789 14139 25823
rect 14749 25789 14783 25823
rect 15577 25789 15611 25823
rect 17785 25789 17819 25823
rect 18153 25789 18187 25823
rect 18429 25789 18463 25823
rect 18705 25789 18739 25823
rect 19073 25789 19107 25823
rect 20729 25789 20763 25823
rect 21097 25789 21131 25823
rect 21281 25789 21315 25823
rect 26249 25789 26283 25823
rect 26341 25789 26375 25823
rect 26617 25789 26651 25823
rect 26893 25789 26927 25823
rect 27077 25789 27111 25823
rect 7665 25721 7699 25755
rect 9597 25721 9631 25755
rect 11989 25721 12023 25755
rect 15761 25721 15795 25755
rect 17877 25721 17911 25755
rect 17969 25721 18003 25755
rect 18889 25721 18923 25755
rect 18981 25721 19015 25755
rect 26433 25721 26467 25755
rect 27905 25721 27939 25755
rect 3893 25653 3927 25687
rect 9781 25653 9815 25687
rect 10057 25653 10091 25687
rect 10701 25653 10735 25687
rect 13461 25653 13495 25687
rect 14197 25653 14231 25687
rect 14933 25653 14967 25687
rect 17601 25653 17635 25687
rect 19533 25653 19567 25687
rect 20085 25653 20119 25687
rect 21005 25653 21039 25687
rect 23213 25653 23247 25687
rect 30481 25653 30515 25687
rect 32137 25653 32171 25687
rect 3065 25449 3099 25483
rect 6101 25449 6135 25483
rect 12081 25449 12115 25483
rect 21465 25449 21499 25483
rect 21557 25449 21591 25483
rect 22017 25449 22051 25483
rect 22477 25449 22511 25483
rect 25237 25449 25271 25483
rect 25973 25449 26007 25483
rect 29101 25449 29135 25483
rect 6377 25381 6411 25415
rect 6469 25381 6503 25415
rect 7389 25381 7423 25415
rect 13645 25381 13679 25415
rect 14105 25381 14139 25415
rect 15761 25381 15795 25415
rect 19257 25381 19291 25415
rect 19349 25381 19383 25415
rect 23029 25381 23063 25415
rect 4813 25313 4847 25347
rect 6285 25313 6319 25347
rect 6653 25313 6687 25347
rect 8033 25313 8067 25347
rect 11805 25313 11839 25347
rect 11897 25313 11931 25347
rect 12081 25313 12115 25347
rect 13737 25313 13771 25347
rect 13829 25313 13863 25347
rect 15853 25313 15887 25347
rect 18153 25313 18187 25347
rect 18797 25313 18831 25347
rect 19073 25313 19107 25347
rect 19441 25313 19475 25347
rect 19717 25313 19751 25347
rect 21925 25313 21959 25347
rect 22569 25313 22603 25347
rect 22753 25313 22787 25347
rect 22937 25313 22971 25347
rect 23121 25313 23155 25347
rect 26617 25313 26651 25347
rect 28825 25313 28859 25347
rect 30297 25313 30331 25347
rect 4537 25245 4571 25279
rect 4905 25245 4939 25279
rect 5549 25245 5583 25279
rect 6745 25245 6779 25279
rect 8309 25245 8343 25279
rect 16405 25245 16439 25279
rect 17877 25245 17911 25279
rect 18981 25245 19015 25279
rect 19993 25245 20027 25279
rect 22109 25245 22143 25279
rect 23489 25245 23523 25279
rect 23765 25245 23799 25279
rect 25329 25245 25363 25279
rect 26433 25245 26467 25279
rect 26525 25245 26559 25279
rect 27077 25245 27111 25279
rect 27629 25245 27663 25279
rect 27813 25245 27847 25279
rect 28733 25245 28767 25279
rect 29837 25245 29871 25279
rect 15577 25177 15611 25211
rect 26985 25177 27019 25211
rect 5917 25109 5951 25143
rect 7665 25109 7699 25143
rect 9781 25109 9815 25143
rect 11621 25109 11655 25143
rect 18613 25109 18647 25143
rect 19625 25109 19659 25143
rect 23305 25109 23339 25143
rect 28457 25109 28491 25143
rect 29285 25109 29319 25143
rect 30205 25109 30239 25143
rect 4721 24905 4755 24939
rect 8585 24905 8619 24939
rect 9229 24905 9263 24939
rect 18429 24905 18463 24939
rect 18613 24905 18647 24939
rect 20545 24905 20579 24939
rect 24225 24905 24259 24939
rect 25421 24905 25455 24939
rect 26328 24905 26362 24939
rect 27813 24905 27847 24939
rect 4169 24769 4203 24803
rect 4261 24769 4295 24803
rect 6101 24769 6135 24803
rect 9873 24769 9907 24803
rect 16405 24769 16439 24803
rect 16681 24769 16715 24803
rect 16819 24769 16853 24803
rect 18061 24769 18095 24803
rect 19349 24769 19383 24803
rect 19901 24769 19935 24803
rect 22845 24769 22879 24803
rect 23581 24769 23615 24803
rect 29009 24769 29043 24803
rect 29285 24769 29319 24803
rect 3065 24701 3099 24735
rect 3341 24701 3375 24735
rect 4353 24701 4387 24735
rect 8493 24701 8527 24735
rect 10057 24701 10091 24735
rect 10241 24701 10275 24735
rect 10977 24701 11011 24735
rect 11069 24701 11103 24735
rect 11161 24701 11195 24735
rect 11253 24701 11287 24735
rect 11621 24701 11655 24735
rect 11805 24701 11839 24735
rect 15761 24701 15795 24735
rect 15945 24701 15979 24735
rect 16957 24701 16991 24735
rect 18705 24701 18739 24735
rect 18889 24701 18923 24735
rect 19073 24701 19107 24735
rect 21005 24701 21039 24735
rect 21557 24701 21591 24735
rect 24317 24701 24351 24735
rect 24409 24701 24443 24735
rect 25513 24701 25547 24735
rect 25881 24701 25915 24735
rect 26065 24701 26099 24735
rect 28825 24701 28859 24735
rect 7849 24633 7883 24667
rect 9597 24633 9631 24667
rect 10149 24633 10183 24667
rect 11437 24633 11471 24667
rect 23213 24633 23247 24667
rect 4997 24565 5031 24599
rect 6377 24565 6411 24599
rect 6929 24565 6963 24599
rect 7481 24565 7515 24599
rect 9689 24565 9723 24599
rect 10793 24565 10827 24599
rect 15577 24565 15611 24599
rect 17601 24565 17635 24599
rect 17969 24565 18003 24599
rect 18429 24565 18463 24599
rect 19717 24565 19751 24599
rect 22569 24565 22603 24599
rect 25789 24565 25823 24599
rect 28273 24565 28307 24599
rect 30757 24565 30791 24599
rect 5825 24361 5859 24395
rect 6653 24361 6687 24395
rect 12633 24361 12667 24395
rect 18153 24361 18187 24395
rect 29377 24361 29411 24395
rect 6837 24293 6871 24327
rect 7757 24293 7791 24327
rect 11897 24293 11931 24327
rect 17969 24293 18003 24327
rect 20637 24293 20671 24327
rect 28181 24293 28215 24327
rect 6101 24225 6135 24259
rect 6193 24225 6227 24259
rect 6469 24225 6503 24259
rect 7665 24225 7699 24259
rect 10333 24225 10367 24259
rect 10885 24225 10919 24259
rect 11558 24225 11592 24259
rect 12541 24225 12575 24259
rect 13185 24225 13219 24259
rect 15485 24225 15519 24259
rect 19349 24225 19383 24259
rect 23673 24225 23707 24259
rect 28641 24225 28675 24259
rect 29561 24225 29595 24259
rect 29653 24225 29687 24259
rect 29745 24225 29779 24259
rect 29883 24225 29917 24259
rect 30849 24225 30883 24259
rect 32229 24225 32263 24259
rect 4077 24157 4111 24191
rect 4353 24157 4387 24191
rect 6561 24157 6595 24191
rect 8033 24157 8067 24191
rect 8309 24157 8343 24191
rect 11069 24157 11103 24191
rect 13461 24157 13495 24191
rect 14933 24157 14967 24191
rect 15393 24157 15427 24191
rect 23029 24157 23063 24191
rect 26709 24157 26743 24191
rect 28457 24157 28491 24191
rect 30021 24157 30055 24191
rect 30665 24157 30699 24191
rect 33425 24157 33459 24191
rect 5917 24089 5951 24123
rect 7205 24089 7239 24123
rect 11253 24089 11287 24123
rect 17601 24089 17635 24123
rect 18889 24089 18923 24123
rect 6837 24021 6871 24055
rect 7573 24021 7607 24055
rect 9781 24021 9815 24055
rect 11621 24021 11655 24055
rect 11732 24021 11766 24055
rect 17141 24021 17175 24055
rect 17509 24021 17543 24055
rect 17969 24021 18003 24055
rect 18613 24021 18647 24055
rect 21925 24021 21959 24055
rect 22477 24021 22511 24055
rect 23581 24021 23615 24055
rect 26617 24021 26651 24055
rect 28825 24021 28859 24055
rect 5181 23817 5215 23851
rect 6101 23817 6135 23851
rect 6745 23817 6779 23851
rect 8217 23817 8251 23851
rect 9965 23817 9999 23851
rect 10333 23817 10367 23851
rect 11621 23817 11655 23851
rect 12909 23817 12943 23851
rect 14013 23817 14047 23851
rect 28273 23817 28307 23851
rect 29929 23817 29963 23851
rect 11437 23749 11471 23783
rect 18337 23749 18371 23783
rect 23673 23749 23707 23783
rect 29745 23749 29779 23783
rect 3525 23681 3559 23715
rect 5733 23681 5767 23715
rect 6101 23681 6135 23715
rect 7941 23681 7975 23715
rect 8033 23681 8067 23715
rect 9781 23681 9815 23715
rect 15577 23681 15611 23715
rect 22201 23681 22235 23715
rect 24041 23681 24075 23715
rect 25789 23681 25823 23715
rect 27629 23681 27663 23715
rect 3065 23613 3099 23647
rect 5089 23613 5123 23647
rect 6929 23613 6963 23647
rect 8309 23613 8343 23647
rect 8953 23613 8987 23647
rect 9045 23613 9079 23647
rect 9597 23613 9631 23647
rect 10057 23613 10091 23647
rect 10241 23613 10275 23647
rect 10701 23613 10735 23647
rect 11621 23613 11655 23647
rect 11713 23613 11747 23647
rect 11897 23613 11931 23647
rect 11989 23613 12023 23647
rect 12082 23613 12116 23647
rect 12357 23613 12391 23647
rect 12633 23613 12667 23647
rect 12725 23613 12759 23647
rect 13645 23613 13679 23647
rect 13921 23613 13955 23647
rect 14841 23613 14875 23647
rect 16405 23613 16439 23647
rect 19073 23613 19107 23647
rect 19625 23613 19659 23647
rect 19901 23613 19935 23647
rect 19993 23613 20027 23647
rect 21005 23613 21039 23647
rect 21925 23613 21959 23647
rect 26617 23613 26651 23647
rect 27445 23613 27479 23647
rect 27767 23613 27801 23647
rect 27905 23613 27939 23647
rect 28089 23613 28123 23647
rect 28549 23613 28583 23647
rect 29653 23613 29687 23647
rect 29837 23613 29871 23647
rect 30297 23613 30331 23647
rect 7573 23545 7607 23579
rect 12909 23545 12943 23579
rect 13737 23545 13771 23579
rect 17877 23545 17911 23579
rect 19809 23545 19843 23579
rect 24317 23545 24351 23579
rect 26065 23545 26099 23579
rect 27997 23545 28031 23579
rect 28457 23545 28491 23579
rect 30113 23545 30147 23579
rect 5917 23477 5951 23511
rect 7021 23477 7055 23511
rect 7481 23477 7515 23511
rect 9229 23477 9263 23511
rect 9413 23477 9447 23511
rect 10885 23477 10919 23511
rect 14197 23477 14231 23511
rect 14933 23477 14967 23511
rect 15761 23477 15795 23511
rect 17325 23477 17359 23511
rect 17969 23477 18003 23511
rect 18981 23477 19015 23511
rect 19441 23477 19475 23511
rect 20177 23477 20211 23511
rect 21097 23477 21131 23511
rect 27261 23477 27295 23511
rect 7757 23273 7791 23307
rect 10701 23273 10735 23307
rect 14473 23273 14507 23307
rect 19809 23273 19843 23307
rect 22201 23273 22235 23307
rect 25053 23273 25087 23307
rect 26157 23273 26191 23307
rect 27813 23273 27847 23307
rect 4169 23205 4203 23239
rect 10149 23205 10183 23239
rect 14381 23205 14415 23239
rect 18613 23205 18647 23239
rect 20269 23205 20303 23239
rect 26525 23205 26559 23239
rect 27261 23205 27295 23239
rect 6009 23137 6043 23171
rect 8033 23137 8067 23171
rect 8217 23137 8251 23171
rect 8493 23137 8527 23171
rect 8677 23137 8711 23171
rect 8769 23137 8803 23171
rect 9965 23137 9999 23171
rect 10609 23137 10643 23171
rect 10769 23137 10803 23171
rect 10891 23137 10925 23171
rect 11069 23137 11103 23171
rect 11805 23137 11839 23171
rect 11897 23137 11931 23171
rect 12081 23137 12115 23171
rect 12357 23137 12391 23171
rect 12541 23137 12575 23171
rect 12725 23137 12759 23171
rect 14933 23137 14967 23171
rect 18521 23137 18555 23171
rect 18705 23137 18739 23171
rect 18889 23137 18923 23171
rect 19993 23137 20027 23171
rect 22569 23137 22603 23171
rect 22661 23137 22695 23171
rect 23489 23137 23523 23171
rect 24041 23137 24075 23171
rect 24961 23137 24995 23171
rect 26341 23137 26375 23171
rect 26433 23137 26467 23171
rect 26643 23137 26677 23171
rect 26801 23137 26835 23171
rect 27077 23137 27111 23171
rect 27353 23137 27387 23171
rect 27537 23137 27571 23171
rect 27997 23137 28031 23171
rect 28089 23137 28123 23171
rect 28273 23137 28307 23171
rect 29285 23137 29319 23171
rect 29653 23137 29687 23171
rect 30205 23137 30239 23171
rect 31125 23137 31159 23171
rect 31769 23137 31803 23171
rect 3433 23069 3467 23103
rect 6285 23069 6319 23103
rect 8309 23069 8343 23103
rect 8861 23069 8895 23103
rect 9689 23069 9723 23103
rect 12265 23069 12299 23103
rect 13737 23069 13771 23103
rect 14197 23069 14231 23103
rect 15209 23069 15243 23103
rect 17141 23069 17175 23103
rect 22753 23069 22787 23103
rect 25881 23069 25915 23103
rect 28181 23069 28215 23103
rect 31217 23069 31251 23103
rect 9781 23001 9815 23035
rect 11069 23001 11103 23035
rect 12173 23001 12207 23035
rect 21741 23001 21775 23035
rect 27445 23001 27479 23035
rect 4077 22933 4111 22967
rect 5457 22933 5491 22967
rect 8033 22933 8067 22967
rect 9505 22933 9539 22967
rect 11621 22933 11655 22967
rect 12633 22933 12667 22967
rect 13185 22933 13219 22967
rect 14841 22933 14875 22967
rect 16681 22933 16715 22967
rect 17785 22933 17819 22967
rect 18337 22933 18371 22967
rect 19257 22933 19291 22967
rect 22109 22933 22143 22967
rect 25237 22933 25271 22967
rect 26893 22933 26927 22967
rect 29653 22933 29687 22967
rect 29837 22933 29871 22967
rect 30297 22933 30331 22967
rect 30941 22933 30975 22967
rect 3065 22729 3099 22763
rect 6101 22729 6135 22763
rect 9229 22729 9263 22763
rect 10425 22729 10459 22763
rect 12541 22729 12575 22763
rect 14473 22729 14507 22763
rect 15761 22729 15795 22763
rect 16589 22729 16623 22763
rect 17785 22729 17819 22763
rect 24304 22729 24338 22763
rect 26157 22729 26191 22763
rect 31033 22729 31067 22763
rect 31309 22729 31343 22763
rect 10977 22661 11011 22695
rect 20729 22661 20763 22695
rect 27905 22661 27939 22695
rect 4537 22593 4571 22627
rect 6745 22593 6779 22627
rect 7021 22593 7055 22627
rect 8861 22593 8895 22627
rect 11989 22593 12023 22627
rect 12357 22593 12391 22627
rect 13001 22593 13035 22627
rect 16313 22593 16347 22627
rect 19809 22593 19843 22627
rect 20085 22593 20119 22627
rect 22477 22593 22511 22627
rect 24041 22593 24075 22627
rect 25789 22593 25823 22627
rect 26801 22593 26835 22627
rect 26893 22593 26927 22627
rect 27169 22593 27203 22627
rect 29285 22593 29319 22627
rect 33057 22593 33091 22627
rect 4813 22525 4847 22559
rect 5089 22525 5123 22559
rect 5457 22525 5491 22559
rect 9045 22525 9079 22559
rect 9321 22525 9355 22559
rect 9781 22525 9815 22559
rect 10793 22525 10827 22559
rect 11161 22525 11195 22559
rect 11897 22525 11931 22559
rect 12265 22525 12299 22559
rect 12725 22525 12759 22559
rect 15485 22525 15519 22559
rect 16681 22525 16715 22559
rect 17233 22525 17267 22559
rect 20177 22525 20211 22559
rect 20361 22525 20395 22559
rect 20545 22525 20579 22559
rect 21097 22525 21131 22559
rect 21189 22525 21223 22559
rect 23765 22525 23799 22559
rect 26341 22525 26375 22559
rect 26663 22525 26697 22559
rect 28089 22525 28123 22559
rect 28273 22525 28307 22559
rect 33333 22525 33367 22559
rect 33977 22525 34011 22559
rect 4997 22457 5031 22491
rect 10609 22457 10643 22491
rect 20453 22457 20487 22491
rect 21833 22457 21867 22491
rect 26433 22457 26467 22491
rect 26525 22457 26559 22491
rect 29561 22457 29595 22491
rect 32781 22457 32815 22491
rect 33241 22457 33275 22491
rect 6561 22389 6595 22423
rect 8493 22389 8527 22423
rect 11345 22389 11379 22423
rect 12081 22389 12115 22423
rect 14933 22389 14967 22423
rect 18061 22389 18095 22423
rect 18337 22389 18371 22423
rect 21005 22389 21039 22423
rect 21925 22389 21959 22423
rect 22845 22389 22879 22423
rect 23857 22389 23891 22423
rect 28181 22389 28215 22423
rect 28457 22389 28491 22423
rect 33793 22389 33827 22423
rect 3433 22185 3467 22219
rect 3893 22185 3927 22219
rect 6009 22185 6043 22219
rect 7757 22185 7791 22219
rect 8033 22185 8067 22219
rect 8401 22185 8435 22219
rect 9689 22185 9723 22219
rect 16221 22185 16255 22219
rect 19993 22185 20027 22219
rect 25237 22185 25271 22219
rect 25513 22185 25547 22219
rect 26525 22185 26559 22219
rect 27261 22185 27295 22219
rect 31861 22185 31895 22219
rect 32229 22185 32263 22219
rect 3801 22117 3835 22151
rect 9873 22117 9907 22151
rect 10057 22117 10091 22151
rect 11713 22117 11747 22151
rect 13185 22117 13219 22151
rect 14749 22117 14783 22151
rect 17969 22117 18003 22151
rect 18429 22117 18463 22151
rect 21465 22117 21499 22151
rect 23213 22117 23247 22151
rect 26893 22117 26927 22151
rect 30389 22117 30423 22151
rect 32381 22117 32415 22151
rect 32597 22117 32631 22151
rect 3341 22049 3375 22083
rect 4250 22049 4284 22083
rect 6193 22049 6227 22083
rect 6285 22049 6319 22083
rect 7665 22049 7699 22083
rect 8217 22049 8251 22083
rect 8493 22049 8527 22083
rect 10149 22049 10183 22083
rect 10333 22049 10367 22083
rect 12081 22049 12115 22083
rect 12357 22049 12391 22083
rect 14105 22049 14139 22083
rect 16957 22049 16991 22083
rect 17325 22049 17359 22083
rect 18889 22049 18923 22083
rect 19257 22049 19291 22083
rect 21925 22049 21959 22083
rect 22937 22049 22971 22083
rect 23489 22049 23523 22083
rect 25605 22049 25639 22083
rect 26525 22049 26559 22083
rect 26617 22049 26651 22083
rect 26801 22049 26835 22083
rect 27077 22049 27111 22083
rect 27353 22049 27387 22083
rect 27813 22049 27847 22083
rect 28181 22049 28215 22083
rect 28641 22049 28675 22083
rect 28917 22049 28951 22083
rect 29469 22049 29503 22083
rect 29561 22049 29595 22083
rect 4077 21981 4111 22015
rect 4537 21981 4571 22015
rect 9045 21981 9079 22015
rect 12173 21981 12207 22015
rect 12265 21981 12299 22015
rect 13829 21981 13863 22015
rect 14013 21981 14047 22015
rect 14473 21981 14507 22015
rect 16865 21981 16899 22015
rect 17233 21981 17267 22015
rect 19073 21981 19107 22015
rect 21741 21981 21775 22015
rect 22845 21981 22879 22015
rect 23305 21981 23339 22015
rect 23765 21981 23799 22015
rect 28273 21981 28307 22015
rect 28733 21981 28767 22015
rect 30113 21981 30147 22015
rect 6653 21913 6687 21947
rect 16589 21913 16623 21947
rect 17601 21913 17635 21947
rect 18153 21913 18187 21947
rect 19441 21913 19475 21947
rect 22661 21913 22695 21947
rect 3249 21845 3283 21879
rect 6929 21845 6963 21879
rect 9597 21845 9631 21879
rect 10333 21845 10367 21879
rect 11621 21845 11655 21879
rect 11897 21845 11931 21879
rect 16681 21845 16715 21879
rect 17969 21845 18003 21879
rect 18521 21845 18555 21879
rect 18797 21845 18831 21879
rect 19809 21845 19843 21879
rect 22017 21845 22051 21879
rect 22385 21845 22419 21879
rect 27629 21845 27663 21879
rect 27905 21845 27939 21879
rect 28917 21845 28951 21879
rect 29101 21845 29135 21879
rect 32413 21845 32447 21879
rect 5457 21641 5491 21675
rect 7849 21641 7883 21675
rect 9873 21641 9907 21675
rect 14013 21641 14047 21675
rect 15117 21641 15151 21675
rect 15853 21641 15887 21675
rect 18153 21641 18187 21675
rect 23489 21641 23523 21675
rect 29469 21641 29503 21675
rect 31585 21641 31619 21675
rect 5273 21573 5307 21607
rect 19441 21573 19475 21607
rect 24869 21573 24903 21607
rect 5641 21505 5675 21539
rect 6101 21505 6135 21539
rect 6745 21505 6779 21539
rect 11345 21505 11379 21539
rect 14473 21505 14507 21539
rect 14657 21505 14691 21539
rect 16405 21505 16439 21539
rect 16681 21505 16715 21539
rect 22753 21505 22787 21539
rect 26065 21505 26099 21539
rect 29653 21505 29687 21539
rect 29929 21505 29963 21539
rect 30205 21505 30239 21539
rect 4813 21437 4847 21471
rect 5733 21437 5767 21471
rect 6193 21437 6227 21471
rect 6377 21437 6411 21471
rect 9597 21437 9631 21471
rect 11437 21437 11471 21471
rect 11529 21437 11563 21471
rect 11621 21437 11655 21471
rect 12265 21437 12299 21471
rect 15945 21437 15979 21471
rect 19165 21437 19199 21471
rect 19441 21437 19475 21471
rect 21005 21437 21039 21471
rect 23581 21437 23615 21471
rect 25697 21437 25731 21471
rect 25881 21437 25915 21471
rect 26617 21437 26651 21471
rect 29745 21437 29779 21471
rect 29837 21437 29871 21471
rect 30113 21437 30147 21471
rect 30297 21437 30331 21471
rect 31033 21437 31067 21471
rect 31677 21437 31711 21471
rect 31861 21437 31895 21471
rect 32597 21437 32631 21471
rect 4537 21369 4571 21403
rect 6009 21369 6043 21403
rect 6285 21369 6319 21403
rect 9137 21369 9171 21403
rect 9781 21369 9815 21403
rect 12541 21369 12575 21403
rect 21281 21369 21315 21403
rect 31217 21369 31251 21403
rect 31401 21369 31435 21403
rect 33793 21369 33827 21403
rect 3065 21301 3099 21335
rect 7113 21301 7147 21335
rect 9505 21301 9539 21335
rect 11805 21301 11839 21335
rect 14749 21301 14783 21335
rect 15393 21301 15427 21335
rect 18889 21301 18923 21335
rect 19901 21301 19935 21335
rect 23029 21301 23063 21335
rect 25697 21301 25731 21335
rect 30389 21301 30423 21335
rect 31861 21301 31895 21335
rect 4629 21097 4663 21131
rect 10977 21097 11011 21131
rect 13553 21097 13587 21131
rect 17785 21097 17819 21131
rect 21373 21097 21407 21131
rect 23765 21097 23799 21131
rect 27813 21097 27847 21131
rect 30313 21097 30347 21131
rect 30481 21097 30515 21131
rect 30865 21097 30899 21131
rect 3249 21029 3283 21063
rect 5641 21029 5675 21063
rect 5733 21029 5767 21063
rect 9505 21029 9539 21063
rect 11621 21029 11655 21063
rect 15025 21029 15059 21063
rect 22385 21029 22419 21063
rect 23949 21029 23983 21063
rect 28181 21029 28215 21063
rect 30113 21029 30147 21063
rect 30665 21029 30699 21063
rect 4445 20961 4479 20995
rect 5549 20961 5583 20995
rect 5917 20961 5951 20995
rect 6101 20961 6135 20995
rect 8953 20961 8987 20995
rect 10517 20961 10551 20995
rect 10885 20961 10919 20995
rect 11069 20961 11103 20995
rect 11437 20961 11471 20995
rect 14473 20961 14507 20995
rect 16865 20961 16899 20995
rect 18337 20961 18371 20995
rect 21005 20961 21039 20995
rect 21189 20961 21223 20995
rect 21649 20961 21683 20995
rect 22661 20961 22695 20995
rect 23857 20961 23891 20995
rect 24041 20961 24075 20995
rect 25605 20961 25639 20995
rect 25789 20961 25823 20995
rect 26985 20961 27019 20995
rect 27077 20961 27111 20995
rect 27445 20961 27479 20995
rect 27721 20961 27755 20995
rect 27997 20961 28031 20995
rect 33793 20961 33827 20995
rect 5273 20893 5307 20927
rect 6377 20893 6411 20927
rect 7849 20893 7883 20927
rect 8217 20893 8251 20927
rect 9045 20893 9079 20927
rect 9321 20893 9355 20927
rect 10241 20893 10275 20927
rect 10333 20893 10367 20927
rect 10426 20893 10460 20927
rect 11161 20893 11195 20927
rect 11805 20893 11839 20927
rect 13645 20893 13679 20927
rect 18613 20893 18647 20927
rect 20085 20893 20119 20927
rect 20821 20893 20855 20927
rect 21557 20893 21591 20927
rect 21925 20893 21959 20927
rect 22017 20893 22051 20927
rect 25329 20893 25363 20927
rect 25421 20893 25455 20927
rect 26525 20893 26559 20927
rect 31125 20893 31159 20927
rect 31769 20893 31803 20927
rect 32597 20893 32631 20927
rect 33333 20893 33367 20927
rect 5365 20825 5399 20859
rect 10057 20825 10091 20859
rect 8861 20757 8895 20791
rect 11253 20757 11287 20791
rect 12357 20757 12391 20791
rect 14289 20757 14323 20791
rect 16313 20757 16347 20791
rect 18153 20757 18187 20791
rect 20269 20757 20303 20791
rect 21189 20757 21223 20791
rect 24317 20757 24351 20791
rect 24685 20757 24719 20791
rect 25881 20757 25915 20791
rect 27353 20757 27387 20791
rect 27629 20757 27663 20791
rect 30297 20757 30331 20791
rect 30849 20757 30883 20791
rect 31033 20757 31067 20791
rect 32045 20757 32079 20791
rect 32781 20757 32815 20791
rect 33885 20757 33919 20791
rect 5181 20553 5215 20587
rect 9045 20553 9079 20587
rect 9873 20553 9907 20587
rect 9965 20553 9999 20587
rect 13829 20553 13863 20587
rect 18613 20553 18647 20587
rect 21005 20553 21039 20587
rect 21373 20553 21407 20587
rect 22385 20553 22419 20587
rect 26065 20553 26099 20587
rect 26433 20553 26467 20587
rect 26985 20553 27019 20587
rect 27629 20553 27663 20587
rect 27905 20553 27939 20587
rect 29469 20553 29503 20587
rect 29929 20553 29963 20587
rect 31953 20553 31987 20587
rect 9505 20485 9539 20519
rect 9597 20485 9631 20519
rect 10149 20485 10183 20519
rect 19625 20485 19659 20519
rect 25881 20485 25915 20519
rect 29009 20485 29043 20519
rect 30665 20485 30699 20519
rect 3617 20417 3651 20451
rect 4261 20417 4295 20451
rect 4537 20417 4571 20451
rect 7481 20417 7515 20451
rect 8493 20417 8527 20451
rect 8677 20417 8711 20451
rect 10425 20417 10459 20451
rect 11069 20417 11103 20451
rect 11345 20417 11379 20451
rect 11713 20417 11747 20451
rect 15577 20417 15611 20451
rect 15761 20417 15795 20451
rect 17509 20417 17543 20451
rect 17601 20417 17635 20451
rect 19165 20417 19199 20451
rect 24133 20417 24167 20451
rect 24409 20417 24443 20451
rect 27997 20417 28031 20451
rect 29285 20417 29319 20451
rect 31309 20417 31343 20451
rect 32229 20417 32263 20451
rect 32505 20417 32539 20451
rect 4077 20349 4111 20383
rect 7849 20349 7883 20383
rect 9413 20349 9447 20383
rect 9689 20349 9723 20383
rect 10977 20349 11011 20383
rect 11437 20349 11471 20383
rect 18521 20349 18555 20383
rect 19073 20349 19107 20383
rect 19441 20349 19475 20383
rect 20177 20349 20211 20383
rect 21097 20349 21131 20383
rect 21557 20349 21591 20383
rect 21649 20349 21683 20383
rect 21925 20349 21959 20383
rect 23673 20349 23707 20383
rect 26249 20349 26283 20383
rect 26525 20349 26559 20383
rect 27169 20349 27203 20383
rect 27353 20349 27387 20383
rect 27629 20349 27663 20383
rect 27721 20349 27755 20383
rect 29193 20349 29227 20383
rect 29653 20349 29687 20383
rect 30573 20349 30607 20383
rect 30757 20349 30791 20383
rect 31033 20349 31067 20383
rect 7205 20281 7239 20315
rect 8401 20281 8435 20315
rect 11621 20281 11655 20315
rect 11989 20281 12023 20315
rect 15301 20281 15335 20315
rect 16037 20281 16071 20315
rect 18429 20281 18463 20315
rect 20453 20281 20487 20315
rect 22017 20281 22051 20315
rect 27445 20281 27479 20315
rect 29745 20281 29779 20315
rect 29961 20281 29995 20315
rect 31585 20281 31619 20315
rect 3709 20213 3743 20247
rect 4169 20213 4203 20247
rect 5733 20213 5767 20247
rect 8033 20213 8067 20247
rect 11161 20213 11195 20247
rect 13461 20213 13495 20247
rect 18245 20213 18279 20247
rect 18981 20213 19015 20247
rect 20085 20213 20119 20247
rect 23765 20213 23799 20247
rect 28641 20213 28675 20247
rect 30113 20213 30147 20247
rect 30941 20213 30975 20247
rect 31493 20213 31527 20247
rect 33977 20213 34011 20247
rect 5273 20009 5307 20043
rect 6193 20009 6227 20043
rect 7757 20009 7791 20043
rect 9137 20009 9171 20043
rect 10609 20009 10643 20043
rect 11621 20009 11655 20043
rect 12909 20009 12943 20043
rect 13369 20009 13403 20043
rect 13737 20009 13771 20043
rect 15485 20009 15519 20043
rect 16313 20009 16347 20043
rect 16773 20009 16807 20043
rect 18889 20009 18923 20043
rect 19349 20009 19383 20043
rect 22845 20009 22879 20043
rect 27077 20009 27111 20043
rect 28917 20009 28951 20043
rect 32321 20009 32355 20043
rect 33057 20009 33091 20043
rect 33149 20009 33183 20043
rect 9597 19941 9631 19975
rect 11805 19941 11839 19975
rect 12081 19941 12115 19975
rect 13829 19941 13863 19975
rect 14197 19941 14231 19975
rect 16681 19941 16715 19975
rect 19993 19941 20027 19975
rect 20453 19941 20487 19975
rect 25329 19941 25363 19975
rect 27997 19941 28031 19975
rect 29561 19941 29595 19975
rect 30849 19941 30883 19975
rect 32505 19941 32539 19975
rect 5365 19873 5399 19907
rect 5733 19873 5767 19907
rect 6009 19873 6043 19907
rect 6745 19873 6779 19907
rect 8585 19873 8619 19907
rect 10425 19873 10459 19907
rect 10885 19873 10919 19907
rect 10977 19873 11011 19907
rect 11345 19873 11379 19907
rect 11713 19873 11747 19907
rect 12265 19873 12299 19907
rect 12357 19873 12391 19907
rect 13001 19873 13035 19907
rect 17417 19873 17451 19907
rect 18337 19873 18371 19907
rect 18981 19873 19015 19907
rect 19625 19873 19659 19907
rect 19717 19873 19751 19907
rect 20177 19873 20211 19907
rect 20913 19873 20947 19907
rect 23121 19873 23155 19907
rect 23305 19873 23339 19907
rect 25237 19873 25271 19907
rect 26065 19873 26099 19907
rect 27261 19873 27295 19907
rect 27721 19873 27755 19907
rect 28273 19873 28307 19907
rect 29101 19873 29135 19907
rect 30573 19873 30607 19907
rect 32597 19873 32631 19907
rect 4537 19805 4571 19839
rect 4813 19805 4847 19839
rect 5641 19805 5675 19839
rect 6101 19805 6135 19839
rect 7113 19805 7147 19839
rect 8033 19805 8067 19839
rect 9045 19805 9079 19839
rect 13921 19805 13955 19839
rect 16957 19805 16991 19839
rect 18613 19805 18647 19839
rect 19073 19805 19107 19839
rect 20085 19805 20119 19839
rect 21097 19805 21131 19839
rect 21373 19805 21407 19839
rect 23213 19805 23247 19839
rect 25973 19805 26007 19839
rect 27445 19805 27479 19839
rect 28181 19805 28215 19839
rect 29285 19805 29319 19839
rect 33241 19805 33275 19839
rect 9597 19737 9631 19771
rect 11069 19737 11103 19771
rect 11989 19737 12023 19771
rect 19441 19737 19475 19771
rect 32689 19737 32723 19771
rect 3065 19669 3099 19703
rect 5457 19669 5491 19703
rect 8861 19669 8895 19703
rect 9781 19669 9815 19703
rect 11161 19669 11195 19703
rect 11437 19669 11471 19703
rect 12081 19669 12115 19703
rect 12541 19669 12575 19703
rect 17509 19669 17543 19703
rect 18061 19669 18095 19703
rect 18429 19669 18463 19703
rect 19165 19669 19199 19703
rect 23489 19669 23523 19703
rect 24973 19669 25007 19703
rect 26157 19669 26191 19703
rect 27261 19669 27295 19703
rect 27997 19669 28031 19703
rect 28457 19669 28491 19703
rect 29469 19669 29503 19703
rect 5089 19465 5123 19499
rect 5273 19465 5307 19499
rect 7008 19465 7042 19499
rect 8585 19465 8619 19499
rect 10241 19465 10275 19499
rect 11345 19465 11379 19499
rect 13277 19465 13311 19499
rect 14289 19465 14323 19499
rect 15853 19465 15887 19499
rect 16313 19465 16347 19499
rect 16681 19465 16715 19499
rect 17049 19465 17083 19499
rect 22109 19465 22143 19499
rect 25053 19465 25087 19499
rect 27537 19465 27571 19499
rect 28089 19397 28123 19431
rect 28917 19397 28951 19431
rect 29653 19397 29687 19431
rect 6009 19329 6043 19363
rect 9873 19329 9907 19363
rect 11345 19329 11379 19363
rect 11713 19329 11747 19363
rect 13001 19329 13035 19363
rect 13645 19329 13679 19363
rect 18889 19329 18923 19363
rect 19257 19329 19291 19363
rect 23765 19329 23799 19363
rect 27445 19329 27479 19363
rect 33793 19329 33827 19363
rect 3249 19261 3283 19295
rect 4445 19261 4479 19295
rect 4721 19261 4755 19295
rect 5089 19261 5123 19295
rect 5641 19261 5675 19295
rect 6745 19261 6779 19295
rect 9137 19261 9171 19295
rect 9965 19261 9999 19295
rect 10609 19261 10643 19295
rect 10701 19261 10735 19295
rect 11253 19261 11287 19295
rect 11805 19261 11839 19295
rect 13185 19261 13219 19295
rect 15117 19261 15151 19295
rect 15301 19261 15335 19295
rect 15945 19261 15979 19295
rect 17141 19261 17175 19295
rect 18981 19261 19015 19295
rect 21097 19261 21131 19295
rect 22017 19261 22051 19295
rect 23857 19261 23891 19295
rect 24409 19261 24443 19295
rect 25237 19261 25271 19295
rect 25329 19261 25363 19295
rect 26709 19261 26743 19295
rect 26801 19261 26835 19295
rect 26985 19261 27019 19295
rect 27169 19261 27203 19295
rect 28273 19261 28307 19295
rect 30113 19261 30147 19295
rect 31769 19261 31803 19295
rect 32781 19261 32815 19295
rect 9505 19193 9539 19227
rect 11529 19193 11563 19227
rect 21005 19193 21039 19227
rect 23949 19193 23983 19227
rect 27077 19193 27111 19227
rect 27287 19193 27321 19227
rect 29745 19193 29779 19227
rect 29929 19193 29963 19227
rect 5549 19125 5583 19159
rect 6653 19125 6687 19159
rect 8493 19125 8527 19159
rect 11069 19125 11103 19159
rect 12265 19125 12299 19159
rect 12449 19125 12483 19159
rect 14565 19125 14599 19159
rect 15393 19125 15427 19159
rect 20729 19125 20763 19159
rect 24317 19125 24351 19159
rect 26065 19125 26099 19159
rect 27721 19125 27755 19159
rect 27813 19125 27847 19159
rect 27905 19125 27939 19159
rect 29101 19125 29135 19159
rect 29285 19125 29319 19159
rect 29377 19125 29411 19159
rect 29469 19125 29503 19159
rect 31217 19125 31251 19159
rect 32505 19125 32539 19159
rect 4169 18921 4203 18955
rect 6929 18921 6963 18955
rect 7389 18921 7423 18955
rect 7757 18921 7791 18955
rect 8953 18921 8987 18955
rect 12265 18921 12299 18955
rect 19441 18921 19475 18955
rect 19625 18921 19659 18955
rect 28089 18921 28123 18955
rect 29377 18921 29411 18955
rect 30205 18921 30239 18955
rect 30297 18921 30331 18955
rect 31861 18921 31895 18955
rect 9965 18853 9999 18887
rect 11069 18853 11103 18887
rect 24593 18853 24627 18887
rect 3065 18785 3099 18819
rect 3617 18785 3651 18819
rect 4261 18785 4295 18819
rect 7021 18785 7055 18819
rect 7665 18785 7699 18819
rect 8585 18785 8619 18819
rect 9045 18785 9079 18819
rect 9597 18785 9631 18819
rect 13185 18785 13219 18819
rect 13921 18785 13955 18819
rect 14289 18785 14323 18819
rect 19073 18785 19107 18819
rect 19809 18785 19843 18819
rect 19901 18785 19935 18819
rect 21189 18785 21223 18819
rect 24317 18785 24351 18819
rect 26249 18785 26283 18819
rect 26433 18785 26467 18819
rect 26801 18785 26835 18819
rect 27445 18785 27479 18819
rect 29193 18785 29227 18819
rect 29561 18785 29595 18819
rect 30021 18785 30055 18819
rect 30113 18785 30147 18819
rect 30573 18785 30607 18819
rect 31953 18785 31987 18819
rect 33517 18785 33551 18819
rect 4537 18717 4571 18751
rect 6009 18717 6043 18751
rect 6101 18717 6135 18751
rect 8401 18717 8435 18751
rect 8493 18717 8527 18751
rect 11253 18717 11287 18751
rect 12357 18717 12391 18751
rect 12449 18717 12483 18751
rect 13461 18717 13495 18751
rect 14565 18717 14599 18751
rect 16405 18717 16439 18751
rect 16681 18717 16715 18751
rect 18153 18717 18187 18751
rect 18889 18717 18923 18751
rect 21005 18717 21039 18751
rect 23489 18717 23523 18751
rect 26065 18717 26099 18751
rect 26525 18717 26559 18751
rect 29653 18717 29687 18751
rect 30481 18717 30515 18751
rect 30757 18717 30791 18751
rect 31401 18717 31435 18751
rect 33057 18717 33091 18751
rect 10793 18649 10827 18683
rect 11897 18649 11931 18683
rect 20361 18649 20395 18683
rect 3249 18581 3283 18615
rect 6745 18581 6779 18615
rect 10609 18581 10643 18615
rect 11805 18581 11839 18615
rect 12909 18581 12943 18615
rect 13829 18581 13863 18615
rect 16037 18581 16071 18615
rect 18337 18581 18371 18615
rect 19441 18581 19475 18615
rect 20085 18581 20119 18615
rect 21373 18581 21407 18615
rect 23213 18581 23247 18615
rect 24133 18581 24167 18615
rect 26341 18581 26375 18615
rect 28641 18581 28675 18615
rect 29561 18581 29595 18615
rect 30849 18581 30883 18615
rect 32045 18581 32079 18615
rect 12062 18377 12096 18411
rect 14473 18377 14507 18411
rect 14565 18377 14599 18411
rect 16773 18377 16807 18411
rect 19073 18377 19107 18411
rect 23029 18377 23063 18411
rect 25789 18377 25823 18411
rect 29469 18377 29503 18411
rect 30665 18377 30699 18411
rect 9045 18309 9079 18343
rect 9965 18309 9999 18343
rect 17601 18309 17635 18343
rect 19533 18309 19567 18343
rect 24133 18309 24167 18343
rect 27997 18309 28031 18343
rect 28549 18309 28583 18343
rect 29561 18309 29595 18343
rect 30849 18309 30883 18343
rect 5273 18241 5307 18275
rect 5733 18241 5767 18275
rect 6193 18241 6227 18275
rect 6469 18241 6503 18275
rect 6586 18241 6620 18275
rect 6745 18241 6779 18275
rect 8493 18241 8527 18275
rect 8585 18241 8619 18275
rect 9689 18241 9723 18275
rect 11437 18241 11471 18275
rect 11805 18241 11839 18275
rect 13553 18241 13587 18275
rect 13829 18241 13863 18275
rect 15025 18241 15059 18275
rect 15117 18241 15151 18275
rect 17325 18241 17359 18275
rect 17760 18241 17794 18275
rect 17877 18241 17911 18275
rect 18705 18241 18739 18275
rect 21281 18241 21315 18275
rect 23581 18241 23615 18275
rect 24777 18241 24811 18275
rect 33517 18241 33551 18275
rect 33701 18241 33735 18275
rect 3341 18173 3375 18207
rect 3801 18173 3835 18207
rect 4629 18173 4663 18207
rect 5549 18173 5583 18207
rect 10149 18173 10183 18207
rect 10425 18173 10459 18207
rect 16405 18173 16439 18207
rect 17233 18173 17267 18207
rect 18245 18173 18279 18207
rect 18521 18173 18555 18207
rect 18613 18173 18647 18207
rect 18797 18173 18831 18207
rect 18981 18173 19015 18207
rect 23305 18173 23339 18207
rect 25513 18173 25547 18207
rect 25697 18173 25731 18207
rect 26617 18173 26651 18207
rect 26801 18173 26835 18207
rect 26985 18173 27019 18207
rect 27169 18173 27203 18207
rect 27905 18173 27939 18207
rect 28424 18173 28458 18207
rect 28825 18173 28859 18207
rect 29101 18173 29135 18207
rect 29929 18173 29963 18207
rect 32965 18173 32999 18207
rect 33425 18173 33459 18207
rect 7849 18105 7883 18139
rect 8677 18105 8711 18139
rect 14933 18105 14967 18139
rect 15761 18105 15795 18139
rect 21557 18105 21591 18139
rect 23213 18105 23247 18139
rect 23765 18105 23799 18139
rect 26065 18105 26099 18139
rect 27721 18105 27755 18139
rect 28300 18105 28334 18139
rect 28917 18105 28951 18139
rect 29285 18105 29319 18139
rect 29837 18105 29871 18139
rect 30481 18105 30515 18139
rect 30697 18105 30731 18139
rect 32689 18105 32723 18139
rect 3433 18037 3467 18071
rect 7389 18037 7423 18071
rect 9137 18037 9171 18071
rect 10333 18037 10367 18071
rect 10885 18037 10919 18071
rect 17141 18037 17175 18071
rect 17969 18037 18003 18071
rect 18337 18037 18371 18071
rect 19993 18037 20027 18071
rect 20545 18037 20579 18071
rect 23673 18037 23707 18071
rect 24225 18037 24259 18071
rect 24961 18037 24995 18071
rect 26893 18037 26927 18071
rect 28733 18037 28767 18071
rect 29193 18037 29227 18071
rect 29745 18037 29779 18071
rect 30113 18037 30147 18071
rect 31217 18037 31251 18071
rect 33057 18037 33091 18071
rect 4997 17833 5031 17867
rect 22661 17833 22695 17867
rect 27721 17833 27755 17867
rect 31769 17833 31803 17867
rect 33609 17833 33643 17867
rect 6929 17765 6963 17799
rect 8309 17765 8343 17799
rect 12173 17765 12207 17799
rect 12909 17765 12943 17799
rect 13461 17765 13495 17799
rect 15853 17765 15887 17799
rect 16037 17765 16071 17799
rect 16865 17765 16899 17799
rect 17785 17765 17819 17799
rect 18981 17765 19015 17799
rect 26249 17765 26283 17799
rect 33885 17765 33919 17799
rect 13185 17697 13219 17731
rect 15761 17697 15795 17731
rect 17325 17697 17359 17731
rect 18521 17697 18555 17731
rect 19533 17697 19567 17731
rect 19717 17697 19751 17731
rect 20177 17697 20211 17731
rect 20637 17697 20671 17731
rect 20913 17697 20947 17731
rect 21373 17697 21407 17731
rect 23489 17697 23523 17731
rect 28181 17697 28215 17731
rect 28457 17697 28491 17731
rect 29377 17697 29411 17731
rect 29561 17697 29595 17731
rect 30113 17697 30147 17731
rect 30297 17697 30331 17731
rect 31217 17697 31251 17731
rect 33793 17697 33827 17731
rect 4537 17629 4571 17663
rect 4813 17629 4847 17663
rect 6469 17629 6503 17663
rect 6745 17629 6779 17663
rect 8033 17629 8067 17663
rect 12265 17629 12299 17663
rect 14933 17629 14967 17663
rect 15025 17629 15059 17663
rect 17233 17629 17267 17663
rect 18705 17629 18739 17663
rect 19349 17629 19383 17663
rect 20269 17629 20303 17663
rect 20453 17629 20487 17663
rect 23765 17629 23799 17663
rect 25973 17629 26007 17663
rect 28365 17629 28399 17663
rect 29193 17629 29227 17663
rect 30481 17629 30515 17663
rect 31861 17629 31895 17663
rect 32137 17629 32171 17663
rect 7113 17561 7147 17595
rect 17785 17561 17819 17595
rect 27997 17561 28031 17595
rect 3065 17493 3099 17527
rect 7757 17493 7791 17527
rect 9781 17493 9815 17527
rect 10885 17493 10919 17527
rect 15669 17493 15703 17527
rect 17049 17493 17083 17527
rect 18337 17493 18371 17527
rect 18521 17493 18555 17527
rect 19809 17493 19843 17527
rect 25237 17493 25271 17527
rect 28457 17493 28491 17527
rect 28641 17493 28675 17527
rect 29561 17493 29595 17527
rect 30205 17493 30239 17527
rect 31033 17493 31067 17527
rect 5549 17289 5583 17323
rect 6285 17289 6319 17323
rect 9597 17289 9631 17323
rect 12357 17289 12391 17323
rect 13829 17289 13863 17323
rect 18613 17289 18647 17323
rect 21465 17289 21499 17323
rect 23029 17289 23063 17323
rect 29745 17289 29779 17323
rect 33057 17289 33091 17323
rect 18521 17221 18555 17255
rect 26985 17221 27019 17255
rect 5089 17153 5123 17187
rect 6193 17153 6227 17187
rect 6929 17153 6963 17187
rect 7205 17153 7239 17187
rect 8769 17153 8803 17187
rect 10885 17153 10919 17187
rect 12633 17153 12667 17187
rect 12725 17153 12759 17187
rect 13645 17153 13679 17187
rect 14289 17153 14323 17187
rect 14381 17153 14415 17187
rect 18178 17153 18212 17187
rect 18705 17153 18739 17187
rect 19257 17153 19291 17187
rect 20729 17153 20763 17187
rect 22017 17153 22051 17187
rect 23581 17153 23615 17187
rect 26065 17153 26099 17187
rect 27997 17153 28031 17187
rect 29469 17153 29503 17187
rect 32689 17153 32723 17187
rect 32965 17153 32999 17187
rect 33609 17153 33643 17187
rect 4261 17085 4295 17119
rect 4997 17085 5031 17119
rect 6469 17085 6503 17119
rect 6561 17085 6595 17119
rect 6837 17085 6871 17119
rect 9321 17085 9355 17119
rect 9689 17085 9723 17119
rect 10241 17085 10275 17119
rect 10609 17085 10643 17119
rect 14841 17085 14875 17119
rect 15577 17085 15611 17119
rect 15761 17085 15795 17119
rect 17693 17085 17727 17119
rect 18061 17085 18095 17119
rect 18429 17085 18463 17119
rect 18981 17085 19015 17119
rect 21097 17085 21131 17119
rect 21833 17085 21867 17119
rect 21925 17085 21959 17119
rect 22385 17085 22419 17119
rect 22937 17085 22971 17119
rect 24317 17085 24351 17119
rect 25145 17085 25179 17119
rect 25881 17085 25915 17119
rect 27721 17085 27755 17119
rect 29561 17085 29595 17119
rect 30389 17085 30423 17119
rect 3249 17017 3283 17051
rect 4905 17017 4939 17051
rect 6653 17017 6687 17051
rect 12817 17017 12851 17051
rect 15301 17017 15335 17051
rect 16037 17017 16071 17051
rect 21005 17017 21039 17051
rect 4537 16949 4571 16983
rect 8677 16949 8711 16983
rect 9965 16949 9999 16983
rect 10333 16949 10367 16983
rect 13185 16949 13219 16983
rect 14197 16949 14231 16983
rect 14933 16949 14967 16983
rect 17509 16949 17543 16983
rect 17969 16949 18003 16983
rect 18337 16949 18371 16983
rect 23765 16949 23799 16983
rect 24501 16949 24535 16983
rect 25237 16949 25271 16983
rect 26709 16949 26743 16983
rect 30573 16949 30607 16983
rect 31217 16949 31251 16983
rect 3893 16745 3927 16779
rect 4721 16745 4755 16779
rect 5549 16745 5583 16779
rect 7021 16745 7055 16779
rect 7757 16745 7791 16779
rect 8953 16745 8987 16779
rect 10885 16745 10919 16779
rect 15945 16745 15979 16779
rect 16313 16745 16347 16779
rect 22385 16745 22419 16779
rect 22845 16745 22879 16779
rect 22937 16745 22971 16779
rect 23949 16745 23983 16779
rect 26065 16745 26099 16779
rect 28825 16745 28859 16779
rect 29745 16745 29779 16779
rect 29837 16745 29871 16779
rect 29929 16745 29963 16779
rect 30363 16745 30397 16779
rect 30763 16745 30797 16779
rect 9965 16677 9999 16711
rect 15485 16677 15519 16711
rect 18153 16677 18187 16711
rect 20177 16677 20211 16711
rect 30573 16677 30607 16711
rect 31861 16677 31895 16711
rect 3801 16609 3835 16643
rect 4261 16609 4295 16643
rect 5273 16609 5307 16643
rect 5457 16609 5491 16643
rect 5733 16609 5767 16643
rect 7665 16609 7699 16643
rect 8493 16609 8527 16643
rect 8585 16609 8619 16643
rect 9045 16609 9079 16643
rect 9689 16609 9723 16643
rect 10333 16609 10367 16643
rect 12725 16609 12759 16643
rect 13185 16609 13219 16643
rect 15853 16609 15887 16643
rect 16957 16609 16991 16643
rect 17601 16609 17635 16643
rect 20453 16609 20487 16643
rect 20637 16609 20671 16643
rect 23857 16609 23891 16643
rect 24179 16609 24213 16643
rect 25605 16609 25639 16643
rect 25973 16609 26007 16643
rect 26249 16609 26283 16643
rect 26341 16609 26375 16643
rect 26433 16609 26467 16643
rect 26617 16609 26651 16643
rect 27077 16609 27111 16643
rect 27169 16609 27203 16643
rect 27537 16609 27571 16643
rect 27813 16609 27847 16643
rect 28181 16609 28215 16643
rect 28365 16609 28399 16643
rect 28733 16609 28767 16643
rect 30113 16609 30147 16643
rect 30665 16609 30699 16643
rect 30849 16609 30883 16643
rect 30941 16609 30975 16643
rect 31033 16609 31067 16643
rect 31677 16609 31711 16643
rect 31769 16609 31803 16643
rect 31953 16609 31987 16643
rect 32229 16609 32263 16643
rect 4353 16541 4387 16575
rect 4537 16541 4571 16575
rect 8309 16541 8343 16575
rect 10977 16541 11011 16575
rect 12449 16541 12483 16575
rect 13461 16541 13495 16575
rect 15669 16541 15703 16575
rect 20913 16541 20947 16575
rect 22753 16541 22787 16575
rect 28457 16541 28491 16575
rect 29561 16541 29595 16575
rect 33057 16541 33091 16575
rect 23305 16473 23339 16507
rect 27813 16473 27847 16507
rect 27997 16473 28031 16507
rect 30205 16473 30239 16507
rect 3157 16405 3191 16439
rect 14933 16405 14967 16439
rect 16773 16405 16807 16439
rect 18705 16405 18739 16439
rect 20361 16405 20395 16439
rect 30389 16405 30423 16439
rect 4813 16201 4847 16235
rect 8217 16201 8251 16235
rect 13185 16201 13219 16235
rect 14013 16201 14047 16235
rect 16037 16201 16071 16235
rect 16773 16201 16807 16235
rect 25145 16201 25179 16235
rect 28825 16201 28859 16235
rect 29469 16201 29503 16235
rect 32045 16201 32079 16235
rect 14565 16133 14599 16167
rect 20729 16133 20763 16167
rect 26433 16133 26467 16167
rect 29745 16133 29779 16167
rect 7205 16065 7239 16099
rect 13093 16065 13127 16099
rect 13829 16065 13863 16099
rect 15025 16065 15059 16099
rect 16589 16065 16623 16099
rect 17417 16065 17451 16099
rect 17693 16065 17727 16099
rect 22753 16065 22787 16099
rect 23029 16065 23063 16099
rect 26525 16065 26559 16099
rect 29653 16065 29687 16099
rect 30205 16065 30239 16099
rect 3065 15997 3099 16031
rect 5089 15997 5123 16031
rect 7941 15997 7975 16031
rect 10425 15997 10459 16031
rect 11161 15997 11195 16031
rect 11345 15997 11379 16031
rect 13921 15997 13955 16031
rect 15117 15997 15151 16031
rect 19625 15997 19659 16031
rect 19901 15997 19935 16031
rect 20545 15997 20579 16031
rect 20729 15997 20763 16031
rect 20913 15997 20947 16031
rect 25237 15997 25271 16031
rect 26709 15997 26743 16031
rect 27261 15997 27295 16031
rect 27353 15997 27387 16031
rect 29377 15997 29411 16031
rect 30021 15997 30055 16031
rect 31861 15997 31895 16031
rect 32137 15997 32171 16031
rect 32781 15997 32815 16031
rect 3341 15929 3375 15963
rect 4997 15929 5031 15963
rect 6929 15929 6963 15963
rect 10149 15929 10183 15963
rect 17969 15929 18003 15963
rect 26065 15929 26099 15963
rect 26249 15929 26283 15963
rect 29653 15929 29687 15963
rect 29745 15929 29779 15963
rect 29929 15929 29963 15963
rect 33793 15929 33827 15963
rect 5457 15861 5491 15895
rect 7297 15861 7331 15895
rect 8677 15861 8711 15895
rect 10609 15861 10643 15895
rect 15209 15861 15243 15895
rect 19441 15861 19475 15895
rect 22201 15861 22235 15895
rect 24501 15861 24535 15895
rect 30849 15861 30883 15895
rect 31677 15861 31711 15895
rect 32413 15861 32447 15895
rect 4905 15657 4939 15691
rect 7021 15657 7055 15691
rect 8033 15657 8067 15691
rect 9045 15657 9079 15691
rect 10241 15657 10275 15691
rect 11529 15657 11563 15691
rect 11989 15657 12023 15691
rect 14105 15657 14139 15691
rect 17325 15657 17359 15691
rect 18705 15657 18739 15691
rect 20913 15657 20947 15691
rect 23581 15657 23615 15691
rect 23857 15657 23891 15691
rect 27169 15657 27203 15691
rect 33149 15657 33183 15691
rect 3249 15589 3283 15623
rect 4721 15589 4755 15623
rect 5825 15589 5859 15623
rect 7481 15589 7515 15623
rect 10701 15589 10735 15623
rect 16589 15589 16623 15623
rect 28733 15589 28767 15623
rect 30297 15589 30331 15623
rect 31861 15589 31895 15623
rect 4353 15521 4387 15555
rect 5457 15521 5491 15555
rect 5641 15521 5675 15555
rect 5917 15521 5951 15555
rect 6009 15521 6043 15555
rect 8217 15521 8251 15555
rect 8401 15521 8435 15555
rect 9137 15521 9171 15555
rect 10609 15521 10643 15555
rect 11069 15521 11103 15555
rect 12081 15521 12115 15555
rect 13345 15521 13379 15555
rect 16313 15521 16347 15555
rect 16497 15521 16531 15555
rect 16681 15521 16715 15555
rect 17601 15521 17635 15555
rect 18889 15521 18923 15555
rect 20545 15521 20579 15555
rect 22385 15521 22419 15555
rect 23213 15521 23247 15555
rect 23673 15521 23707 15555
rect 23765 15521 23799 15555
rect 27445 15521 27479 15555
rect 27537 15521 27571 15555
rect 28089 15521 28123 15555
rect 28641 15521 28675 15555
rect 29193 15521 29227 15555
rect 33793 15521 33827 15555
rect 6377 15453 6411 15487
rect 8861 15453 8895 15487
rect 9597 15453 9631 15487
rect 14197 15453 14231 15487
rect 14473 15453 14507 15487
rect 16957 15453 16991 15487
rect 17141 15453 17175 15487
rect 17233 15453 17267 15487
rect 17509 15453 17543 15487
rect 19349 15453 19383 15487
rect 21465 15453 21499 15487
rect 28917 15453 28951 15487
rect 30021 15453 30055 15487
rect 6193 15385 6227 15419
rect 7113 15385 7147 15419
rect 7665 15385 7699 15419
rect 9505 15385 9539 15419
rect 12449 15385 12483 15419
rect 31769 15385 31803 15419
rect 7481 15317 7515 15351
rect 11161 15317 11195 15351
rect 13277 15317 13311 15351
rect 15945 15317 15979 15351
rect 16865 15317 16899 15351
rect 18061 15317 18095 15351
rect 19993 15317 20027 15351
rect 21833 15317 21867 15351
rect 23029 15317 23063 15351
rect 27721 15317 27755 15351
rect 28181 15317 28215 15351
rect 33885 15317 33919 15351
rect 4905 15113 4939 15147
rect 6009 15113 6043 15147
rect 6377 15113 6411 15147
rect 6837 15113 6871 15147
rect 7849 15113 7883 15147
rect 11069 15113 11103 15147
rect 14841 15113 14875 15147
rect 19625 15113 19659 15147
rect 23811 15113 23845 15147
rect 31309 15113 31343 15147
rect 33609 15113 33643 15147
rect 3801 15045 3835 15079
rect 5181 15045 5215 15079
rect 5733 15045 5767 15079
rect 17509 15045 17543 15079
rect 18613 15045 18647 15079
rect 19809 15045 19843 15079
rect 20177 15045 20211 15079
rect 23213 15045 23247 15079
rect 3709 14977 3743 15011
rect 4353 14977 4387 15011
rect 10609 14977 10643 15011
rect 11897 14977 11931 15011
rect 13921 14977 13955 15011
rect 15301 14977 15335 15011
rect 16865 14977 16899 15011
rect 17877 14977 17911 15011
rect 18521 14977 18555 15011
rect 20085 14977 20119 15011
rect 21097 14977 21131 15011
rect 21189 14977 21223 15011
rect 21925 14977 21959 15011
rect 25605 14977 25639 15011
rect 27077 14977 27111 15011
rect 31861 14977 31895 15011
rect 4261 14909 4295 14943
rect 5917 14909 5951 14943
rect 7067 14909 7101 14943
rect 7205 14909 7239 14943
rect 7481 14909 7515 14943
rect 8677 14909 8711 14943
rect 10333 14909 10367 14943
rect 10977 14909 11011 14943
rect 11621 14909 11655 14943
rect 14749 14909 14783 14943
rect 14841 14909 14875 14943
rect 15393 14909 15427 14943
rect 15853 14909 15887 14943
rect 17601 14909 17635 14943
rect 17785 14909 17819 14943
rect 18613 14909 18647 14943
rect 18705 14909 18739 14943
rect 19441 14909 19475 14943
rect 19993 14909 20027 14943
rect 20913 14909 20947 14943
rect 22293 14909 22327 14943
rect 22477 14909 22511 14943
rect 23121 14909 23155 14943
rect 23305 14909 23339 14943
rect 25237 14909 25271 14943
rect 26065 14909 26099 14943
rect 26709 14909 26743 14943
rect 29101 14909 29135 14943
rect 29837 14909 29871 14943
rect 30021 14909 30055 14943
rect 31401 14909 31435 14943
rect 31677 14909 31711 14943
rect 7297 14841 7331 14875
rect 8033 14841 8067 14875
rect 9689 14841 9723 14875
rect 13645 14841 13679 14875
rect 14933 14841 14967 14875
rect 16589 14841 16623 14875
rect 18889 14841 18923 14875
rect 20545 14841 20579 14875
rect 21808 14841 21842 14875
rect 23029 14841 23063 14875
rect 27353 14841 27387 14875
rect 32137 14841 32171 14875
rect 3065 14773 3099 14807
rect 4169 14773 4203 14807
rect 6929 14773 6963 14807
rect 9045 14773 9079 14807
rect 9781 14773 9815 14807
rect 10793 14773 10827 14807
rect 11529 14773 11563 14807
rect 14197 14773 14231 14807
rect 14473 14773 14507 14807
rect 15577 14773 15611 14807
rect 17693 14773 17727 14807
rect 19349 14773 19383 14807
rect 21557 14773 21591 14807
rect 21649 14773 21683 14807
rect 22017 14773 22051 14807
rect 29285 14773 29319 14807
rect 30665 14773 30699 14807
rect 31585 14773 31619 14807
rect 4905 14569 4939 14603
rect 6653 14569 6687 14603
rect 7757 14569 7791 14603
rect 13921 14569 13955 14603
rect 15577 14569 15611 14603
rect 22661 14569 22695 14603
rect 24041 14569 24075 14603
rect 24777 14569 24811 14603
rect 25605 14569 25639 14603
rect 26709 14569 26743 14603
rect 27721 14569 27755 14603
rect 29745 14569 29779 14603
rect 29837 14569 29871 14603
rect 3341 14501 3375 14535
rect 5917 14501 5951 14535
rect 6009 14501 6043 14535
rect 22845 14501 22879 14535
rect 26203 14501 26237 14535
rect 28457 14501 28491 14535
rect 29377 14501 29411 14535
rect 31309 14501 31343 14535
rect 3065 14433 3099 14467
rect 5825 14433 5859 14467
rect 6193 14433 6227 14467
rect 7481 14433 7515 14467
rect 8217 14433 8251 14467
rect 13277 14433 13311 14467
rect 13829 14433 13863 14467
rect 14197 14433 14231 14467
rect 15025 14433 15059 14467
rect 16313 14433 16347 14467
rect 16405 14433 16439 14467
rect 17509 14433 17543 14467
rect 17601 14433 17635 14467
rect 17785 14433 17819 14467
rect 17877 14433 17911 14467
rect 20453 14433 20487 14467
rect 20545 14433 20579 14467
rect 20821 14433 20855 14467
rect 22937 14433 22971 14467
rect 24869 14433 24903 14467
rect 25789 14433 25823 14467
rect 25973 14433 26007 14467
rect 26341 14433 26375 14467
rect 26433 14433 26467 14467
rect 26525 14433 26559 14467
rect 27813 14433 27847 14467
rect 29101 14433 29135 14467
rect 29193 14433 29227 14467
rect 29469 14433 29503 14467
rect 29561 14433 29595 14467
rect 31585 14433 31619 14467
rect 32781 14433 32815 14467
rect 5457 14365 5491 14399
rect 8309 14365 8343 14399
rect 8585 14365 8619 14399
rect 10057 14365 10091 14399
rect 10425 14365 10459 14399
rect 10701 14365 10735 14399
rect 12173 14365 12207 14399
rect 12265 14365 12299 14399
rect 14105 14365 14139 14399
rect 14565 14365 14599 14399
rect 16681 14365 16715 14399
rect 17325 14365 17359 14399
rect 20085 14365 20119 14399
rect 20361 14365 20395 14399
rect 20913 14365 20947 14399
rect 21189 14365 21223 14399
rect 26065 14365 26099 14399
rect 27077 14365 27111 14399
rect 32873 14365 32907 14399
rect 33057 14365 33091 14399
rect 4813 14297 4847 14331
rect 6285 14297 6319 14331
rect 6837 14297 6871 14331
rect 5641 14229 5675 14263
rect 6653 14229 6687 14263
rect 8125 14229 8159 14263
rect 12909 14229 12943 14263
rect 14841 14229 14875 14263
rect 15669 14229 15703 14263
rect 18613 14229 18647 14263
rect 23213 14229 23247 14263
rect 23673 14229 23707 14263
rect 29009 14229 29043 14263
rect 32413 14229 32447 14263
rect 33517 14229 33551 14263
rect 4721 14025 4755 14059
rect 4997 14025 5031 14059
rect 6837 14025 6871 14059
rect 8677 14025 8711 14059
rect 9137 14025 9171 14059
rect 10057 14025 10091 14059
rect 11069 14025 11103 14059
rect 13645 14025 13679 14059
rect 14749 14025 14783 14059
rect 16865 14025 16899 14059
rect 17141 14025 17175 14059
rect 18797 14025 18831 14059
rect 19901 14025 19935 14059
rect 22293 14025 22327 14059
rect 25881 14025 25915 14059
rect 26065 14025 26099 14059
rect 27077 14025 27111 14059
rect 32321 14025 32355 14059
rect 33241 14025 33275 14059
rect 8953 13957 8987 13991
rect 12909 13957 12943 13991
rect 14197 13957 14231 13991
rect 15761 13957 15795 13991
rect 17509 13957 17543 13991
rect 25697 13957 25731 13991
rect 3249 13889 3283 13923
rect 5825 13889 5859 13923
rect 7205 13889 7239 13923
rect 9597 13889 9631 13923
rect 9689 13889 9723 13923
rect 10793 13889 10827 13923
rect 11529 13889 11563 13923
rect 11713 13889 11747 13923
rect 13461 13889 13495 13923
rect 15393 13889 15427 13923
rect 16405 13889 16439 13923
rect 22937 13889 22971 13923
rect 23096 13889 23130 13923
rect 23489 13889 23523 13923
rect 24593 13889 24627 13923
rect 25421 13889 25455 13923
rect 26893 13889 26927 13923
rect 27169 13889 27203 13923
rect 30021 13889 30055 13923
rect 32873 13889 32907 13923
rect 33793 13889 33827 13923
rect 4445 13821 4479 13855
rect 5089 13821 5123 13855
rect 5641 13821 5675 13855
rect 6929 13821 6963 13855
rect 10149 13821 10183 13855
rect 11897 13821 11931 13855
rect 12541 13821 12575 13855
rect 14381 13821 14415 13855
rect 14473 13821 14507 13855
rect 14657 13821 14691 13855
rect 14933 13821 14967 13855
rect 15255 13821 15289 13855
rect 15761 13821 15795 13855
rect 15945 13821 15979 13855
rect 16037 13821 16071 13855
rect 16496 13821 16530 13855
rect 16589 13821 16623 13855
rect 16681 13821 16715 13855
rect 17785 13821 17819 13855
rect 17969 13821 18003 13855
rect 18705 13821 18739 13855
rect 20729 13821 20763 13855
rect 20913 13821 20947 13855
rect 21188 13821 21222 13855
rect 21281 13821 21315 13855
rect 21557 13821 21591 13855
rect 21649 13821 21683 13855
rect 21833 13821 21867 13855
rect 21925 13821 21959 13855
rect 22109 13821 22143 13855
rect 23213 13821 23247 13855
rect 23949 13821 23983 13855
rect 24133 13821 24167 13855
rect 24409 13821 24443 13855
rect 26249 13821 26283 13855
rect 26341 13821 26375 13855
rect 26433 13821 26467 13855
rect 26617 13821 26651 13855
rect 26709 13821 26743 13855
rect 26801 13821 26835 13855
rect 27077 13821 27111 13855
rect 29101 13821 29135 13855
rect 29377 13821 29411 13855
rect 29561 13821 29595 13855
rect 29837 13821 29871 13855
rect 30389 13821 30423 13855
rect 30665 13821 30699 13855
rect 30757 13821 30791 13855
rect 31217 13821 31251 13855
rect 31401 13821 31435 13855
rect 31493 13821 31527 13855
rect 9505 13753 9539 13787
rect 11437 13753 11471 13787
rect 12909 13753 12943 13787
rect 15025 13753 15059 13787
rect 15117 13753 15151 13787
rect 18245 13753 18279 13787
rect 27445 13753 27479 13787
rect 30205 13753 30239 13787
rect 30573 13753 30607 13787
rect 5549 13685 5583 13719
rect 6469 13685 6503 13719
rect 13369 13685 13403 13719
rect 14013 13685 14047 13719
rect 14565 13685 14599 13719
rect 16957 13685 16991 13719
rect 17141 13685 17175 13719
rect 18153 13685 18187 13719
rect 20085 13685 20119 13719
rect 24225 13685 24259 13719
rect 28917 13685 28951 13719
rect 29193 13685 29227 13719
rect 30941 13685 30975 13719
rect 4629 13481 4663 13515
rect 6653 13481 6687 13515
rect 7849 13481 7883 13515
rect 9321 13481 9355 13515
rect 9597 13481 9631 13515
rect 10425 13481 10459 13515
rect 11253 13481 11287 13515
rect 11621 13481 11655 13515
rect 13461 13481 13495 13515
rect 14473 13481 14507 13515
rect 15761 13481 15795 13515
rect 16865 13481 16899 13515
rect 17601 13481 17635 13515
rect 20637 13481 20671 13515
rect 21649 13481 21683 13515
rect 23857 13481 23891 13515
rect 25881 13481 25915 13515
rect 27445 13481 27479 13515
rect 29469 13481 29503 13515
rect 30849 13481 30883 13515
rect 6101 13413 6135 13447
rect 9965 13413 9999 13447
rect 10517 13413 10551 13447
rect 13670 13413 13704 13447
rect 26157 13413 26191 13447
rect 26867 13413 26901 13447
rect 26985 13413 27019 13447
rect 28273 13413 28307 13447
rect 28733 13413 28767 13447
rect 30481 13413 30515 13447
rect 32781 13413 32815 13447
rect 4261 13345 4295 13379
rect 6377 13345 6411 13379
rect 6837 13345 6871 13379
rect 8217 13345 8251 13379
rect 10149 13345 10183 13379
rect 13185 13345 13219 13379
rect 13553 13345 13587 13379
rect 15025 13345 15059 13379
rect 15577 13345 15611 13379
rect 16037 13345 16071 13379
rect 16313 13345 16347 13379
rect 16497 13345 16531 13379
rect 16957 13345 16991 13379
rect 17233 13345 17267 13379
rect 17785 13345 17819 13379
rect 17969 13345 18003 13379
rect 19073 13345 19107 13379
rect 19166 13345 19200 13379
rect 20453 13345 20487 13379
rect 20729 13345 20763 13379
rect 21741 13345 21775 13379
rect 22201 13345 22235 13379
rect 23949 13345 23983 13379
rect 24593 13345 24627 13379
rect 24685 13345 24719 13379
rect 26065 13345 26099 13379
rect 26249 13345 26283 13379
rect 26367 13345 26401 13379
rect 27077 13345 27111 13379
rect 27169 13345 27203 13379
rect 28181 13345 28215 13379
rect 28365 13345 28399 13379
rect 28641 13345 28675 13379
rect 28825 13345 28859 13379
rect 29009 13345 29043 13379
rect 30205 13345 30239 13379
rect 30389 13345 30423 13379
rect 30573 13345 30607 13379
rect 32597 13345 32631 13379
rect 32873 13345 32907 13379
rect 33977 13345 34011 13379
rect 3249 13277 3283 13311
rect 7481 13277 7515 13311
rect 8401 13277 8435 13311
rect 11805 13277 11839 13311
rect 14197 13277 14231 13311
rect 14381 13277 14415 13311
rect 16589 13277 16623 13311
rect 17141 13277 17175 13311
rect 20269 13277 20303 13311
rect 21005 13277 21039 13311
rect 22017 13277 22051 13311
rect 22753 13277 22787 13311
rect 24041 13277 24075 13311
rect 24501 13277 24535 13311
rect 25145 13277 25179 13311
rect 25697 13277 25731 13311
rect 26525 13277 26559 13311
rect 26709 13277 26743 13311
rect 27353 13277 27387 13311
rect 27997 13277 28031 13311
rect 29193 13277 29227 13311
rect 32321 13277 32355 13311
rect 13829 13209 13863 13243
rect 14841 13209 14875 13243
rect 20177 13209 20211 13243
rect 23489 13209 23523 13243
rect 8033 13141 8067 13175
rect 8769 13141 8803 13175
rect 12357 13141 12391 13175
rect 13001 13141 13035 13175
rect 15945 13141 15979 13175
rect 16589 13141 16623 13175
rect 17049 13141 17083 13175
rect 17417 13141 17451 13175
rect 17969 13141 18003 13175
rect 19257 13141 19291 13175
rect 22201 13141 22235 13175
rect 22385 13141 22419 13175
rect 23305 13141 23339 13175
rect 25053 13141 25087 13175
rect 30113 13141 30147 13175
rect 33793 13141 33827 13175
rect 3433 12937 3467 12971
rect 3801 12937 3835 12971
rect 9965 12937 9999 12971
rect 13829 12937 13863 12971
rect 16221 12937 16255 12971
rect 16773 12937 16807 12971
rect 16865 12937 16899 12971
rect 17877 12937 17911 12971
rect 19257 12937 19291 12971
rect 20637 12937 20671 12971
rect 22845 12937 22879 12971
rect 25145 12937 25179 12971
rect 26065 12937 26099 12971
rect 27721 12937 27755 12971
rect 29009 12937 29043 12971
rect 31861 12937 31895 12971
rect 21465 12869 21499 12903
rect 33793 12869 33827 12903
rect 7573 12801 7607 12835
rect 11345 12801 11379 12835
rect 11529 12801 11563 12835
rect 13737 12801 13771 12835
rect 14381 12801 14415 12835
rect 15209 12801 15243 12835
rect 15485 12801 15519 12835
rect 16129 12801 16163 12835
rect 16405 12801 16439 12835
rect 18797 12801 18831 12835
rect 20085 12801 20119 12835
rect 23397 12801 23431 12835
rect 23673 12801 23707 12835
rect 25789 12801 25823 12835
rect 27445 12801 27479 12835
rect 31309 12801 31343 12835
rect 3893 12733 3927 12767
rect 4629 12733 4663 12767
rect 5733 12733 5767 12767
rect 7113 12733 7147 12767
rect 7389 12733 7423 12767
rect 7849 12733 7883 12767
rect 8769 12733 8803 12767
rect 8953 12733 8987 12767
rect 9137 12733 9171 12767
rect 10333 12733 10367 12767
rect 11897 12733 11931 12767
rect 11989 12733 12023 12767
rect 16037 12733 16071 12767
rect 16497 12733 16531 12767
rect 16589 12733 16623 12767
rect 16773 12733 16807 12767
rect 17049 12733 17083 12767
rect 17417 12733 17451 12767
rect 17509 12733 17543 12767
rect 17601 12733 17635 12767
rect 18981 12733 19015 12767
rect 19073 12733 19107 12767
rect 19349 12733 19383 12767
rect 19625 12733 19659 12767
rect 19717 12733 19751 12767
rect 26617 12733 26651 12767
rect 27353 12733 27387 12767
rect 27905 12733 27939 12767
rect 29193 12733 29227 12767
rect 29561 12733 29595 12767
rect 30389 12733 30423 12767
rect 33977 12733 34011 12767
rect 8861 12665 8895 12699
rect 12265 12665 12299 12699
rect 15761 12665 15795 12699
rect 17141 12665 17175 12699
rect 17233 12665 17267 12699
rect 18245 12665 18279 12699
rect 19993 12665 20027 12699
rect 21557 12665 21591 12699
rect 27261 12665 27295 12699
rect 28089 12665 28123 12699
rect 4537 12597 4571 12631
rect 5273 12597 5307 12631
rect 6377 12597 6411 12631
rect 6469 12597 6503 12631
rect 7205 12597 7239 12631
rect 8493 12597 8527 12631
rect 8585 12597 8619 12631
rect 9597 12597 9631 12631
rect 10885 12597 10919 12631
rect 11253 12597 11287 12631
rect 11805 12597 11839 12631
rect 15853 12597 15887 12631
rect 17868 12597 17902 12631
rect 19441 12597 19475 12631
rect 25237 12597 25271 12631
rect 26893 12597 26927 12631
rect 30205 12597 30239 12631
rect 31033 12597 31067 12631
rect 3617 12393 3651 12427
rect 3985 12393 4019 12427
rect 6837 12393 6871 12427
rect 11989 12393 12023 12427
rect 12357 12393 12391 12427
rect 12909 12393 12943 12427
rect 13185 12393 13219 12427
rect 13553 12393 13587 12427
rect 13645 12393 13679 12427
rect 14657 12393 14691 12427
rect 17049 12393 17083 12427
rect 18797 12393 18831 12427
rect 19266 12393 19300 12427
rect 19809 12393 19843 12427
rect 20729 12393 20763 12427
rect 23949 12393 23983 12427
rect 26249 12393 26283 12427
rect 26525 12393 26559 12427
rect 28641 12393 28675 12427
rect 29469 12393 29503 12427
rect 30297 12393 30331 12427
rect 33517 12393 33551 12427
rect 5917 12325 5951 12359
rect 6561 12325 6595 12359
rect 8677 12325 8711 12359
rect 10517 12325 10551 12359
rect 16865 12325 16899 12359
rect 18337 12325 18371 12359
rect 18889 12325 18923 12359
rect 26893 12325 26927 12359
rect 28825 12325 28859 12359
rect 29745 12325 29779 12359
rect 29837 12325 29871 12359
rect 31769 12325 31803 12359
rect 3341 12257 3375 12291
rect 6193 12257 6227 12291
rect 6331 12257 6365 12291
rect 6469 12257 6503 12291
rect 6677 12257 6711 12291
rect 8217 12257 8251 12291
rect 10241 12257 10275 12291
rect 12817 12257 12851 12291
rect 14289 12257 14323 12291
rect 14657 12257 14691 12291
rect 14841 12257 14875 12291
rect 14933 12257 14967 12291
rect 16497 12257 16531 12291
rect 19901 12257 19935 12291
rect 20913 12257 20947 12291
rect 21465 12257 21499 12291
rect 21741 12257 21775 12291
rect 23489 12257 23523 12291
rect 23857 12257 23891 12291
rect 24409 12257 24443 12291
rect 24593 12257 24627 12291
rect 26709 12257 26743 12291
rect 26985 12257 27019 12291
rect 29009 12257 29043 12291
rect 29193 12257 29227 12291
rect 29285 12257 29319 12291
rect 29561 12257 29595 12291
rect 29929 12257 29963 12291
rect 32045 12257 32079 12291
rect 4077 12189 4111 12223
rect 4169 12189 4203 12223
rect 7481 12189 7515 12223
rect 8401 12189 8435 12223
rect 13737 12189 13771 12223
rect 15301 12189 15335 12223
rect 15485 12189 15519 12223
rect 15761 12189 15795 12223
rect 16313 12189 16347 12223
rect 20269 12189 20303 12223
rect 21097 12189 21131 12223
rect 22293 12189 22327 12223
rect 22569 12189 22603 12223
rect 25329 12189 25363 12223
rect 25467 12189 25501 12223
rect 25605 12189 25639 12223
rect 32689 12189 32723 12223
rect 15098 12121 15132 12155
rect 15209 12121 15243 12155
rect 18613 12121 18647 12155
rect 25053 12121 25087 12155
rect 30113 12121 30147 12155
rect 3433 12053 3467 12087
rect 4445 12053 4479 12087
rect 6929 12053 6963 12087
rect 8125 12053 8159 12087
rect 10149 12053 10183 12087
rect 12725 12053 12759 12087
rect 14381 12053 14415 12087
rect 16865 12053 16899 12087
rect 19257 12053 19291 12087
rect 19441 12053 19475 12087
rect 23673 12053 23707 12087
rect 27077 12053 27111 12087
rect 32137 12053 32171 12087
rect 33057 12053 33091 12087
rect 3065 11849 3099 11883
rect 5273 11849 5307 11883
rect 5457 11849 5491 11883
rect 6377 11849 6411 11883
rect 6745 11849 6779 11883
rect 8769 11849 8803 11883
rect 9597 11849 9631 11883
rect 12449 11849 12483 11883
rect 13001 11849 13035 11883
rect 14105 11849 14139 11883
rect 14381 11849 14415 11883
rect 18521 11849 18555 11883
rect 18705 11849 18739 11883
rect 21373 11849 21407 11883
rect 22661 11849 22695 11883
rect 27064 11849 27098 11883
rect 28549 11849 28583 11883
rect 31309 11849 31343 11883
rect 31953 11849 31987 11883
rect 32137 11849 32171 11883
rect 12817 11781 12851 11815
rect 15761 11781 15795 11815
rect 16589 11781 16623 11815
rect 17325 11781 17359 11815
rect 25697 11781 25731 11815
rect 4537 11713 4571 11747
rect 6009 11713 6043 11747
rect 8493 11713 8527 11747
rect 13461 11713 13495 11747
rect 15209 11713 15243 11747
rect 15945 11713 15979 11747
rect 16037 11713 16071 11747
rect 16129 11713 16163 11747
rect 16957 11713 16991 11747
rect 18797 11713 18831 11747
rect 19349 11713 19383 11747
rect 22937 11713 22971 11747
rect 23213 11713 23247 11747
rect 26801 11713 26835 11747
rect 32781 11713 32815 11747
rect 33517 11713 33551 11747
rect 4813 11645 4847 11679
rect 6469 11645 6503 11679
rect 9689 11645 9723 11679
rect 11529 11645 11563 11679
rect 11989 11645 12023 11679
rect 13185 11645 13219 11679
rect 13369 11645 13403 11679
rect 14289 11645 14323 11679
rect 14473 11645 14507 11679
rect 15577 11645 15611 11679
rect 17141 11645 17175 11679
rect 18889 11645 18923 11679
rect 19441 11645 19475 11679
rect 19625 11645 19659 11679
rect 20085 11645 20119 11679
rect 21005 11645 21039 11679
rect 21649 11645 21683 11679
rect 21833 11645 21867 11679
rect 24961 11645 24995 11679
rect 25697 11645 25731 11679
rect 25881 11645 25915 11679
rect 29193 11645 29227 11679
rect 30573 11645 30607 11679
rect 31401 11645 31435 11679
rect 33057 11645 33091 11679
rect 5917 11577 5951 11611
rect 8217 11577 8251 11611
rect 24869 11577 24903 11611
rect 29929 11577 29963 11611
rect 32505 11577 32539 11611
rect 5825 11509 5859 11543
rect 11253 11509 11287 11543
rect 17693 11509 17727 11543
rect 20729 11509 20763 11543
rect 24685 11509 24719 11543
rect 29837 11509 29871 11543
rect 32597 11509 32631 11543
rect 8861 11305 8895 11339
rect 11345 11305 11379 11339
rect 13645 11305 13679 11339
rect 15577 11305 15611 11339
rect 19257 11305 19291 11339
rect 19993 11305 20027 11339
rect 26065 11305 26099 11339
rect 28181 11305 28215 11339
rect 29009 11305 29043 11339
rect 30849 11305 30883 11339
rect 3249 11237 3283 11271
rect 6101 11237 6135 11271
rect 7665 11237 7699 11271
rect 11161 11237 11195 11271
rect 13001 11237 13035 11271
rect 16313 11237 16347 11271
rect 16681 11237 16715 11271
rect 16773 11237 16807 11271
rect 19717 11237 19751 11271
rect 22385 11237 22419 11271
rect 24133 11237 24167 11271
rect 25605 11237 25639 11271
rect 29377 11237 29411 11271
rect 31033 11237 31067 11271
rect 32137 11237 32171 11271
rect 33885 11237 33919 11271
rect 4445 11169 4479 11203
rect 5457 11169 5491 11203
rect 8585 11169 8619 11203
rect 10793 11169 10827 11203
rect 12449 11169 12483 11203
rect 12541 11169 12575 11203
rect 13553 11169 13587 11203
rect 14197 11169 14231 11203
rect 14749 11169 14783 11203
rect 15209 11169 15243 11203
rect 16865 11169 16899 11203
rect 17601 11169 17635 11203
rect 17693 11169 17727 11203
rect 17877 11169 17911 11203
rect 19165 11169 19199 11203
rect 19349 11169 19383 11203
rect 19901 11169 19935 11203
rect 22477 11169 22511 11203
rect 23121 11169 23155 11203
rect 25697 11169 25731 11203
rect 27261 11169 27295 11203
rect 28273 11169 28307 11203
rect 28641 11169 28675 11203
rect 28825 11169 28859 11203
rect 29101 11169 29135 11203
rect 31125 11169 31159 11203
rect 33793 11169 33827 11203
rect 5089 11101 5123 11135
rect 8033 11101 8067 11135
rect 10333 11101 10367 11135
rect 10609 11101 10643 11135
rect 12081 11101 12115 11135
rect 13737 11101 13771 11135
rect 16129 11101 16163 11135
rect 17325 11101 17359 11135
rect 20361 11101 20395 11135
rect 21925 11101 21959 11135
rect 22569 11101 22603 11135
rect 23489 11101 23523 11135
rect 24869 11101 24903 11135
rect 25513 11101 25547 11135
rect 26433 11101 26467 11135
rect 27905 11101 27939 11135
rect 31861 11101 31895 11135
rect 33609 11101 33643 11135
rect 12265 11033 12299 11067
rect 14105 11033 14139 11067
rect 22017 11033 22051 11067
rect 23213 11033 23247 11067
rect 5917 10965 5951 10999
rect 11161 10965 11195 10999
rect 11529 10965 11563 10999
rect 13185 10965 13219 10999
rect 14565 10965 14599 10999
rect 15945 10965 15979 10999
rect 17049 10965 17083 10999
rect 17509 10965 17543 10999
rect 17693 10965 17727 10999
rect 18061 10965 18095 10999
rect 18613 10965 18647 10999
rect 21005 10965 21039 10999
rect 21281 10965 21315 10999
rect 24225 10965 24259 10999
rect 27353 10965 27387 10999
rect 4555 10761 4589 10795
rect 8861 10761 8895 10795
rect 9781 10761 9815 10795
rect 11345 10761 11379 10795
rect 11700 10761 11734 10795
rect 16957 10761 16991 10795
rect 18889 10761 18923 10795
rect 23121 10761 23155 10795
rect 24961 10761 24995 10795
rect 26065 10761 26099 10795
rect 28365 10761 28399 10795
rect 6193 10693 6227 10727
rect 9965 10693 9999 10727
rect 14565 10693 14599 10727
rect 17785 10693 17819 10727
rect 18429 10693 18463 10727
rect 5549 10625 5583 10659
rect 5733 10625 5767 10659
rect 8033 10625 8067 10659
rect 11437 10625 11471 10659
rect 19625 10625 19659 10659
rect 23213 10625 23247 10659
rect 23489 10625 23523 10659
rect 25605 10625 25639 10659
rect 28917 10625 28951 10659
rect 33793 10625 33827 10659
rect 4813 10557 4847 10591
rect 5081 10557 5115 10591
rect 8309 10557 8343 10591
rect 8493 10557 8527 10591
rect 8677 10557 8711 10591
rect 8953 10557 8987 10591
rect 9229 10557 9263 10591
rect 9413 10557 9447 10591
rect 9597 10557 9631 10591
rect 10057 10557 10091 10591
rect 10793 10557 10827 10591
rect 10977 10557 11011 10591
rect 11161 10557 11195 10591
rect 15301 10557 15335 10591
rect 15761 10557 15795 10591
rect 15945 10557 15979 10591
rect 16313 10557 16347 10591
rect 17049 10557 17083 10591
rect 19165 10557 19199 10591
rect 19257 10557 19291 10591
rect 20545 10557 20579 10591
rect 20913 10557 20947 10591
rect 21373 10557 21407 10591
rect 27813 10557 27847 10591
rect 28733 10557 28767 10591
rect 29745 10557 29779 10591
rect 29929 10557 29963 10591
rect 30757 10557 30791 10591
rect 30849 10557 30883 10591
rect 32597 10557 32631 10591
rect 7757 10489 7791 10523
rect 8401 10489 8435 10523
rect 9505 10489 9539 10523
rect 11069 10489 11103 10523
rect 13277 10489 13311 10523
rect 17325 10489 17359 10523
rect 19717 10489 19751 10523
rect 21649 10489 21683 10523
rect 27537 10489 27571 10523
rect 29193 10489 29227 10523
rect 3065 10421 3099 10455
rect 5181 10421 5215 10455
rect 5825 10421 5859 10455
rect 6285 10421 6319 10455
rect 8125 10421 8159 10455
rect 10333 10421 10367 10455
rect 13185 10421 13219 10455
rect 15393 10421 15427 10455
rect 15853 10421 15887 10455
rect 20637 10421 20671 10455
rect 21097 10421 21131 10455
rect 25053 10421 25087 10455
rect 28825 10421 28859 10455
rect 30573 10421 30607 10455
rect 3617 10217 3651 10251
rect 6285 10217 6319 10251
rect 8309 10217 8343 10251
rect 9321 10217 9355 10251
rect 14013 10217 14047 10251
rect 16037 10217 16071 10251
rect 17049 10217 17083 10251
rect 17325 10217 17359 10251
rect 17693 10217 17727 10251
rect 18153 10217 18187 10251
rect 20085 10217 20119 10251
rect 23121 10217 23155 10251
rect 23949 10217 23983 10251
rect 25973 10217 26007 10251
rect 26525 10217 26559 10251
rect 31769 10217 31803 10251
rect 3433 10149 3467 10183
rect 4077 10149 4111 10183
rect 4169 10149 4203 10183
rect 4721 10149 4755 10183
rect 8953 10149 8987 10183
rect 9873 10149 9907 10183
rect 11529 10149 11563 10183
rect 14565 10149 14599 10183
rect 16957 10149 16991 10183
rect 18613 10149 18647 10183
rect 30113 10149 30147 10183
rect 3525 10081 3559 10115
rect 3985 10081 4019 10115
rect 4353 10081 4387 10115
rect 4445 10081 4479 10115
rect 7205 10081 7239 10115
rect 11253 10081 11287 10115
rect 14289 10081 14323 10115
rect 16589 10081 16623 10115
rect 17785 10081 17819 10115
rect 18337 10081 18371 10115
rect 23213 10081 23247 10115
rect 24961 10081 24995 10115
rect 26065 10081 26099 10115
rect 27445 10081 27479 10115
rect 27537 10081 27571 10115
rect 30389 10081 30423 10115
rect 30481 10081 30515 10115
rect 33977 10081 34011 10115
rect 6193 10013 6227 10047
rect 6837 10013 6871 10047
rect 13001 10013 13035 10047
rect 13369 10013 13403 10047
rect 16313 10013 16347 10047
rect 16681 10013 16715 10047
rect 17166 10013 17200 10047
rect 17601 10013 17635 10047
rect 20453 10013 20487 10047
rect 20729 10013 20763 10047
rect 22201 10013 22235 10047
rect 22293 10013 22327 10047
rect 23673 10013 23707 10047
rect 23857 10013 23891 10047
rect 24409 10013 24443 10047
rect 25697 10013 25731 10047
rect 26249 10013 26283 10047
rect 26433 10013 26467 10047
rect 27629 10013 27663 10047
rect 7665 9945 7699 9979
rect 24317 9945 24351 9979
rect 26893 9945 26927 9979
rect 3801 9877 3835 9911
rect 8585 9877 8619 9911
rect 11161 9877 11195 9911
rect 22937 9877 22971 9911
rect 25145 9877 25179 9911
rect 27077 9877 27111 9911
rect 28641 9877 28675 9911
rect 33793 9877 33827 9911
rect 11713 9673 11747 9707
rect 13277 9673 13311 9707
rect 14841 9673 14875 9707
rect 16865 9673 16899 9707
rect 17049 9673 17083 9707
rect 29561 9673 29595 9707
rect 31401 9673 31435 9707
rect 5457 9605 5491 9639
rect 7113 9605 7147 9639
rect 14657 9605 14691 9639
rect 18797 9605 18831 9639
rect 22569 9605 22603 9639
rect 26065 9605 26099 9639
rect 3249 9537 3283 9571
rect 4629 9537 4663 9571
rect 5273 9537 5307 9571
rect 6009 9537 6043 9571
rect 6101 9537 6135 9571
rect 7021 9537 7055 9571
rect 7665 9537 7699 9571
rect 8861 9537 8895 9571
rect 15485 9537 15519 9571
rect 16589 9537 16623 9571
rect 20177 9537 20211 9571
rect 21465 9537 21499 9571
rect 22477 9537 22511 9571
rect 23121 9537 23155 9571
rect 24133 9537 24167 9571
rect 25605 9537 25639 9571
rect 26617 9537 26651 9571
rect 26985 9537 27019 9571
rect 29009 9537 29043 9571
rect 30941 9537 30975 9571
rect 4261 9469 4295 9503
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 7481 9469 7515 9503
rect 8493 9469 8527 9503
rect 13369 9469 13403 9503
rect 13829 9469 13863 9503
rect 14197 9469 14231 9503
rect 15301 9469 15335 9503
rect 17233 9469 17267 9503
rect 17509 9469 17543 9503
rect 18705 9469 18739 9503
rect 19717 9469 19751 9503
rect 20361 9469 20395 9503
rect 23029 9469 23063 9503
rect 23857 9469 23891 9503
rect 30205 9469 30239 9503
rect 18061 9401 18095 9435
rect 18245 9401 18279 9435
rect 20545 9401 20579 9435
rect 21281 9401 21315 9435
rect 27261 9401 27295 9435
rect 29193 9401 29227 9435
rect 29653 9401 29687 9435
rect 6377 9333 6411 9367
rect 7573 9333 7607 9367
rect 7941 9333 7975 9367
rect 9965 9333 9999 9367
rect 13093 9333 13127 9367
rect 15209 9333 15243 9367
rect 15945 9333 15979 9367
rect 17417 9333 17451 9367
rect 17785 9333 17819 9367
rect 18521 9333 18555 9367
rect 19165 9333 19199 9367
rect 20913 9333 20947 9367
rect 21373 9333 21407 9367
rect 21833 9333 21867 9367
rect 22937 9333 22971 9367
rect 28733 9333 28767 9367
rect 29101 9333 29135 9367
rect 30389 9333 30423 9367
rect 4629 9129 4663 9163
rect 9689 9129 9723 9163
rect 10241 9129 10275 9163
rect 10471 9129 10505 9163
rect 17764 9129 17798 9163
rect 20453 9129 20487 9163
rect 20821 9129 20855 9163
rect 24869 9129 24903 9163
rect 25237 9129 25271 9163
rect 29561 9129 29595 9163
rect 8125 9061 8159 9095
rect 17969 9061 18003 9095
rect 23489 9061 23523 9095
rect 31585 9061 31619 9095
rect 4537 8993 4571 9027
rect 5365 8993 5399 9027
rect 6101 8993 6135 9027
rect 8217 8993 8251 9027
rect 9229 8993 9263 9027
rect 9873 8993 9907 9027
rect 11897 8993 11931 9027
rect 14933 8993 14967 9027
rect 17141 8993 17175 9027
rect 18797 8993 18831 9027
rect 19650 8993 19684 9027
rect 21557 8993 21591 9027
rect 25329 8993 25363 9027
rect 25421 8993 25455 9027
rect 26755 8993 26789 9027
rect 28825 8993 28859 9027
rect 28917 8993 28951 9027
rect 29653 8993 29687 9027
rect 31677 8993 31711 9027
rect 4169 8925 4203 8959
rect 5273 8925 5307 8959
rect 6377 8925 6411 8959
rect 9505 8925 9539 8959
rect 12265 8925 12299 8959
rect 14657 8925 14691 8959
rect 16773 8925 16807 8959
rect 17509 8925 17543 8959
rect 18613 8925 18647 8959
rect 19533 8925 19567 8959
rect 19809 8925 19843 8959
rect 21373 8925 21407 8959
rect 21833 8925 21867 8959
rect 24133 8925 24167 8959
rect 24685 8925 24719 8959
rect 24777 8925 24811 8959
rect 25697 8925 25731 8959
rect 25881 8925 25915 8959
rect 26617 8925 26651 8959
rect 26893 8925 26927 8959
rect 28457 8925 28491 8959
rect 28733 8925 28767 8959
rect 29929 8925 29963 8959
rect 32597 8925 32631 8959
rect 17601 8857 17635 8891
rect 19257 8857 19291 8891
rect 23305 8857 23339 8891
rect 26341 8857 26375 8891
rect 27813 8857 27847 8891
rect 31401 8857 31435 8891
rect 3617 8789 3651 8823
rect 4445 8789 4479 8823
rect 6009 8789 6043 8823
rect 7849 8789 7883 8823
rect 8585 8789 8619 8823
rect 9505 8789 9539 8823
rect 13185 8789 13219 8823
rect 15485 8789 15519 8823
rect 17785 8789 17819 8823
rect 27537 8789 27571 8823
rect 32045 8789 32079 8823
rect 3328 8585 3362 8619
rect 5089 8585 5123 8619
rect 5457 8585 5491 8619
rect 6941 8585 6975 8619
rect 10793 8585 10827 8619
rect 14657 8585 14691 8619
rect 15393 8585 15427 8619
rect 18521 8585 18555 8619
rect 18889 8585 18923 8619
rect 19257 8585 19291 8619
rect 20545 8585 20579 8619
rect 23029 8585 23063 8619
rect 23581 8585 23615 8619
rect 25329 8585 25363 8619
rect 26249 8585 26283 8619
rect 27353 8585 27387 8619
rect 29561 8585 29595 8619
rect 33011 8585 33045 8619
rect 33425 8585 33459 8619
rect 11529 8517 11563 8551
rect 12265 8517 12299 8551
rect 13921 8517 13955 8551
rect 17417 8517 17451 8551
rect 25605 8517 25639 8551
rect 33793 8517 33827 8551
rect 3065 8449 3099 8483
rect 7205 8449 7239 8483
rect 7389 8449 7423 8483
rect 9137 8449 9171 8483
rect 9781 8449 9815 8483
rect 13093 8449 13127 8483
rect 13369 8449 13403 8483
rect 14013 8449 14047 8483
rect 14841 8449 14875 8483
rect 15945 8449 15979 8483
rect 16773 8449 16807 8483
rect 17141 8449 17175 8483
rect 19257 8449 19291 8483
rect 19467 8449 19501 8483
rect 21281 8449 21315 8483
rect 21741 8449 21775 8483
rect 22155 8449 22189 8483
rect 27997 8449 28031 8483
rect 30573 8449 30607 8483
rect 31217 8449 31251 8483
rect 11621 8381 11655 8415
rect 13553 8381 13587 8415
rect 14933 8381 14967 8415
rect 17258 8381 17292 8415
rect 17693 8381 17727 8415
rect 17877 8381 17911 8415
rect 17969 8381 18003 8415
rect 19625 8381 19659 8415
rect 19809 8381 19843 8415
rect 21097 8381 21131 8415
rect 22017 8381 22051 8415
rect 22293 8381 22327 8415
rect 22937 8381 22971 8415
rect 23213 8381 23247 8415
rect 23305 8381 23339 8415
rect 23673 8381 23707 8415
rect 24869 8381 24903 8415
rect 27077 8381 27111 8415
rect 27537 8381 27571 8415
rect 27629 8381 27663 8415
rect 28089 8381 28123 8415
rect 28733 8381 28767 8415
rect 29009 8381 29043 8415
rect 29193 8381 29227 8415
rect 29377 8381 29411 8415
rect 30205 8381 30239 8415
rect 31585 8381 31619 8415
rect 33977 8381 34011 8415
rect 7665 8313 7699 8347
rect 10241 8313 10275 8347
rect 13461 8313 13495 8347
rect 15209 8313 15243 8347
rect 16681 8313 16715 8347
rect 17049 8313 17083 8347
rect 20085 8313 20119 8347
rect 28365 8313 28399 8347
rect 28457 8313 28491 8347
rect 29285 8313 29319 8347
rect 29929 8313 29963 8347
rect 4813 8245 4847 8279
rect 9229 8245 9263 8279
rect 15409 8245 15443 8279
rect 15577 8245 15611 8279
rect 17509 8245 17543 8279
rect 24317 8245 24351 8279
rect 26709 8245 26743 8279
rect 26985 8245 27019 8279
rect 27813 8245 27847 8279
rect 3249 8041 3283 8075
rect 3801 8041 3835 8075
rect 5733 8041 5767 8075
rect 6469 8041 6503 8075
rect 8125 8041 8159 8075
rect 8493 8041 8527 8075
rect 8585 8041 8619 8075
rect 10609 8041 10643 8075
rect 12449 8041 12483 8075
rect 14289 8041 14323 8075
rect 14657 8041 14691 8075
rect 16497 8041 16531 8075
rect 17417 8041 17451 8075
rect 18153 8041 18187 8075
rect 23121 8041 23155 8075
rect 25697 8041 25731 8075
rect 27077 8041 27111 8075
rect 28089 8041 28123 8075
rect 31217 8041 31251 8075
rect 32045 8041 32079 8075
rect 7481 7973 7515 8007
rect 17785 7973 17819 8007
rect 19901 7973 19935 8007
rect 21925 7973 21959 8007
rect 24133 7973 24167 8007
rect 32413 7973 32447 8007
rect 3065 7905 3099 7939
rect 4169 7905 4203 7939
rect 4261 7905 4295 7939
rect 4629 7905 4663 7939
rect 5641 7905 5675 7939
rect 5917 7905 5951 7939
rect 6101 7905 6135 7939
rect 6285 7905 6319 7939
rect 6377 7905 6411 7939
rect 7021 7905 7055 7939
rect 9045 7905 9079 7939
rect 9229 7905 9263 7939
rect 9781 7905 9815 7939
rect 10149 7905 10183 7939
rect 10701 7905 10735 7939
rect 11621 7905 11655 7939
rect 11805 7905 11839 7939
rect 11897 7905 11931 7939
rect 11989 7905 12023 7939
rect 14473 7905 14507 7939
rect 14657 7905 14691 7939
rect 14749 7905 14783 7939
rect 16865 7905 16899 7939
rect 17141 7905 17175 7939
rect 18337 7905 18371 7939
rect 18797 7905 18831 7939
rect 19073 7905 19107 7939
rect 19165 7905 19199 7939
rect 19441 7905 19475 7939
rect 27169 7905 27203 7939
rect 32873 7905 32907 7939
rect 33425 7905 33459 7939
rect 3709 7837 3743 7871
rect 4353 7837 4387 7871
rect 5181 7837 5215 7871
rect 8769 7837 8803 7871
rect 9505 7837 9539 7871
rect 9873 7837 9907 7871
rect 10241 7837 10275 7871
rect 11437 7837 11471 7871
rect 13001 7837 13035 7871
rect 13737 7837 13771 7871
rect 15025 7837 15059 7871
rect 17417 7837 17451 7871
rect 23857 7837 23891 7871
rect 25605 7837 25639 7871
rect 26249 7837 26283 7871
rect 26433 7837 26467 7871
rect 28641 7837 28675 7871
rect 28917 7837 28951 7871
rect 31033 7837 31067 7871
rect 31769 7837 31803 7871
rect 32505 7837 32539 7871
rect 32689 7837 32723 7871
rect 18797 7769 18831 7803
rect 19717 7769 19751 7803
rect 30389 7769 30423 7803
rect 6101 7701 6135 7735
rect 10425 7701 10459 7735
rect 11069 7701 11103 7735
rect 12173 7701 12207 7735
rect 13185 7701 13219 7735
rect 16957 7701 16991 7735
rect 17233 7701 17267 7735
rect 18429 7701 18463 7735
rect 19533 7701 19567 7735
rect 21189 7701 21223 7735
rect 22385 7701 22419 7735
rect 22753 7701 22787 7735
rect 23765 7701 23799 7735
rect 27813 7701 27847 7735
rect 30481 7701 30515 7735
rect 7481 7497 7515 7531
rect 10149 7497 10183 7531
rect 12160 7497 12194 7531
rect 13645 7497 13679 7531
rect 15301 7497 15335 7531
rect 15761 7497 15795 7531
rect 16681 7497 16715 7531
rect 18797 7497 18831 7531
rect 24501 7497 24535 7531
rect 25421 7497 25455 7531
rect 26065 7497 26099 7531
rect 28181 7497 28215 7531
rect 29009 7497 29043 7531
rect 29548 7497 29582 7531
rect 31585 7497 31619 7531
rect 3525 7361 3559 7395
rect 7021 7361 7055 7395
rect 11161 7361 11195 7395
rect 11897 7361 11931 7395
rect 16221 7361 16255 7395
rect 16405 7361 16439 7395
rect 17325 7361 17359 7395
rect 19809 7361 19843 7395
rect 21465 7361 21499 7395
rect 21557 7361 21591 7395
rect 22569 7361 22603 7395
rect 24961 7361 24995 7395
rect 25053 7361 25087 7395
rect 27813 7361 27847 7395
rect 29285 7361 29319 7395
rect 31769 7361 31803 7395
rect 32045 7361 32079 7395
rect 3157 7293 3191 7327
rect 5273 7293 5307 7327
rect 6101 7293 6135 7327
rect 6193 7293 6227 7327
rect 6377 7293 6411 7327
rect 6561 7293 6595 7327
rect 8677 7293 8711 7327
rect 11345 7293 11379 7327
rect 14289 7293 14323 7327
rect 14657 7293 14691 7327
rect 14933 7293 14967 7327
rect 16129 7293 16163 7327
rect 16773 7293 16807 7327
rect 17049 7293 17083 7327
rect 19349 7293 19383 7327
rect 19717 7293 19751 7327
rect 20545 7293 20579 7327
rect 21097 7293 21131 7327
rect 21189 7293 21223 7327
rect 21833 7293 21867 7327
rect 21925 7293 21959 7327
rect 22201 7293 22235 7327
rect 25329 7293 25363 7327
rect 28089 7293 28123 7327
rect 28365 7293 28399 7327
rect 31401 7293 31435 7327
rect 31493 7293 31527 7327
rect 6469 7225 6503 7259
rect 14565 7225 14599 7259
rect 15117 7225 15151 7259
rect 22017 7225 22051 7259
rect 22845 7225 22879 7259
rect 27537 7225 27571 7259
rect 31309 7225 31343 7259
rect 4629 7157 4663 7191
rect 5457 7157 5491 7191
rect 6745 7157 6779 7191
rect 8585 7157 8619 7191
rect 10609 7157 10643 7191
rect 11437 7157 11471 7191
rect 13737 7157 13771 7191
rect 20453 7157 20487 7191
rect 20637 7157 20671 7191
rect 20913 7157 20947 7191
rect 21649 7157 21683 7191
rect 24317 7157 24351 7191
rect 24869 7157 24903 7191
rect 25789 7157 25823 7191
rect 31033 7157 31067 7191
rect 33517 7157 33551 7191
rect 3801 6953 3835 6987
rect 6101 6953 6135 6987
rect 12909 6953 12943 6987
rect 18797 6953 18831 6987
rect 25329 6953 25363 6987
rect 26525 6953 26559 6987
rect 27721 6953 27755 6987
rect 30481 6953 30515 6987
rect 32137 6953 32171 6987
rect 3709 6885 3743 6919
rect 4537 6885 4571 6919
rect 16957 6885 16991 6919
rect 18153 6885 18187 6919
rect 27813 6885 27847 6919
rect 30849 6885 30883 6919
rect 3341 6817 3375 6851
rect 4261 6817 4295 6851
rect 8309 6817 8343 6851
rect 13737 6817 13771 6851
rect 13829 6817 13863 6851
rect 16037 6817 16071 6851
rect 17417 6817 17451 6851
rect 22109 6817 22143 6851
rect 23489 6817 23523 6851
rect 25513 6817 25547 6851
rect 26617 6817 26651 6851
rect 27077 6817 27111 6851
rect 27997 6817 28031 6851
rect 28641 6817 28675 6851
rect 30941 6817 30975 6851
rect 32321 6817 32355 6851
rect 33425 6817 33459 6851
rect 3617 6749 3651 6783
rect 7573 6749 7607 6783
rect 7849 6749 7883 6783
rect 9229 6749 9263 6783
rect 9505 6749 9539 6783
rect 10977 6749 11011 6783
rect 11069 6749 11103 6783
rect 12449 6749 12483 6783
rect 16313 6749 16347 6783
rect 18981 6749 19015 6783
rect 19717 6749 19751 6783
rect 19993 6749 20027 6783
rect 21465 6749 21499 6783
rect 23029 6749 23063 6783
rect 25697 6749 25731 6783
rect 26341 6749 26375 6783
rect 28181 6749 28215 6783
rect 31125 6749 31159 6783
rect 15117 6681 15151 6715
rect 26985 6681 27019 6715
rect 3249 6613 3283 6647
rect 4169 6613 4203 6647
rect 6009 6613 6043 6647
rect 11713 6613 11747 6647
rect 11897 6613 11931 6647
rect 19625 6613 19659 6647
rect 21557 6613 21591 6647
rect 22477 6613 22511 6647
rect 24777 6613 24811 6647
rect 25973 6613 26007 6647
rect 30113 6613 30147 6647
rect 31493 6613 31527 6647
rect 3985 6409 4019 6443
rect 5733 6409 5767 6443
rect 12357 6409 12391 6443
rect 13093 6409 13127 6443
rect 15485 6409 15519 6443
rect 21452 6409 21486 6443
rect 22937 6409 22971 6443
rect 23489 6409 23523 6443
rect 25145 6409 25179 6443
rect 25513 6409 25547 6443
rect 30021 6409 30055 6443
rect 30849 6409 30883 6443
rect 33701 6409 33735 6443
rect 7481 6341 7515 6375
rect 18797 6341 18831 6375
rect 26985 6341 27019 6375
rect 29009 6341 29043 6375
rect 29101 6341 29135 6375
rect 30389 6341 30423 6375
rect 32781 6341 32815 6375
rect 6837 6273 6871 6307
rect 7573 6273 7607 6307
rect 10333 6273 10367 6307
rect 10609 6273 10643 6307
rect 13461 6273 13495 6307
rect 16589 6273 16623 6307
rect 17233 6273 17267 6307
rect 19257 6273 19291 6307
rect 19349 6273 19383 6307
rect 19809 6273 19843 6307
rect 20177 6273 20211 6307
rect 20545 6273 20579 6307
rect 21189 6273 21223 6307
rect 27077 6273 27111 6307
rect 28824 6273 28858 6307
rect 29653 6273 29687 6307
rect 31769 6273 31803 6307
rect 32137 6273 32171 6307
rect 33425 6273 33459 6307
rect 3065 6205 3099 6239
rect 5273 6205 5307 6239
rect 6469 6205 6503 6239
rect 9597 6205 9631 6239
rect 9873 6205 9907 6239
rect 12541 6205 12575 6239
rect 12909 6205 12943 6239
rect 13185 6205 13219 6239
rect 16037 6205 16071 6239
rect 16957 6205 16991 6239
rect 19165 6205 19199 6239
rect 19901 6205 19935 6239
rect 23213 6205 23247 6239
rect 23673 6205 23707 6239
rect 23765 6205 23799 6239
rect 24041 6205 24075 6239
rect 24317 6205 24351 6239
rect 25237 6205 25271 6239
rect 26433 6205 26467 6239
rect 26801 6205 26835 6239
rect 28089 6205 28123 6239
rect 28457 6205 28491 6239
rect 28732 6205 28766 6239
rect 32413 6205 32447 6239
rect 33793 6205 33827 6239
rect 7849 6137 7883 6171
rect 9505 6137 9539 6171
rect 10885 6137 10919 6171
rect 12725 6137 12759 6171
rect 12817 6137 12851 6171
rect 20269 6137 20303 6171
rect 23121 6137 23155 6171
rect 23857 6137 23891 6171
rect 26617 6137 26651 6171
rect 26709 6137 26743 6171
rect 28365 6137 28399 6171
rect 3249 6069 3283 6103
rect 5917 6069 5951 6103
rect 9321 6069 9355 6103
rect 14933 6069 14967 6103
rect 18705 6069 18739 6103
rect 19625 6069 19659 6103
rect 24961 6069 24995 6103
rect 26249 6069 26283 6103
rect 27721 6069 27755 6103
rect 31217 6069 31251 6103
rect 32321 6069 32355 6103
rect 32873 6069 32907 6103
rect 3065 5865 3099 5899
rect 7481 5865 7515 5899
rect 8033 5865 8067 5899
rect 9045 5865 9079 5899
rect 10241 5865 10275 5899
rect 10701 5865 10735 5899
rect 11437 5865 11471 5899
rect 12173 5865 12207 5899
rect 13553 5865 13587 5899
rect 14013 5865 14047 5899
rect 17969 5865 18003 5899
rect 21741 5865 21775 5899
rect 23581 5865 23615 5899
rect 27353 5865 27387 5899
rect 30389 5865 30423 5899
rect 30849 5865 30883 5899
rect 31217 5865 31251 5899
rect 7757 5797 7791 5831
rect 11805 5797 11839 5831
rect 17417 5797 17451 5831
rect 21005 5797 21039 5831
rect 23121 5797 23155 5831
rect 28365 5797 28399 5831
rect 30757 5797 30791 5831
rect 32045 5797 32079 5831
rect 33885 5797 33919 5831
rect 4813 5729 4847 5763
rect 6377 5729 6411 5763
rect 7573 5729 7607 5763
rect 7849 5729 7883 5763
rect 10333 5729 10367 5763
rect 11345 5729 11379 5763
rect 11621 5729 11655 5763
rect 11713 5729 11747 5763
rect 11989 5729 12023 5763
rect 12265 5729 12299 5763
rect 13645 5729 13679 5763
rect 14565 5729 14599 5763
rect 14749 5729 14783 5763
rect 17509 5729 17543 5763
rect 17877 5729 17911 5763
rect 21097 5729 21131 5763
rect 24225 5729 24259 5763
rect 25513 5729 25547 5763
rect 26709 5729 26743 5763
rect 27629 5729 27663 5763
rect 28641 5729 28675 5763
rect 31769 5729 31803 5763
rect 33793 5729 33827 5763
rect 4537 5661 4571 5695
rect 5641 5661 5675 5695
rect 6745 5661 6779 5695
rect 8585 5661 8619 5695
rect 9229 5661 9263 5695
rect 10425 5661 10459 5695
rect 12357 5661 12391 5695
rect 13001 5661 13035 5695
rect 13737 5661 13771 5695
rect 15025 5661 15059 5695
rect 17141 5661 17175 5695
rect 19073 5661 19107 5695
rect 19349 5661 19383 5695
rect 24363 5661 24397 5695
rect 24501 5661 24535 5695
rect 25237 5661 25271 5695
rect 25421 5661 25455 5695
rect 25697 5661 25731 5695
rect 26157 5661 26191 5695
rect 26433 5661 26467 5695
rect 26571 5661 26605 5695
rect 27813 5661 27847 5695
rect 28917 5661 28951 5695
rect 30573 5661 30607 5695
rect 31493 5661 31527 5695
rect 5825 5593 5859 5627
rect 9873 5593 9907 5627
rect 13185 5593 13219 5627
rect 22845 5593 22879 5627
rect 24777 5593 24811 5627
rect 5089 5525 5123 5559
rect 7297 5525 7331 5559
rect 9781 5525 9815 5559
rect 16497 5525 16531 5559
rect 16589 5525 16623 5559
rect 18705 5525 18739 5559
rect 20821 5525 20855 5559
rect 27537 5525 27571 5559
rect 33517 5525 33551 5559
rect 7941 5321 7975 5355
rect 14105 5321 14139 5355
rect 14289 5321 14323 5355
rect 14841 5321 14875 5355
rect 15945 5321 15979 5355
rect 19533 5321 19567 5355
rect 20453 5321 20487 5355
rect 21741 5321 21775 5355
rect 23305 5321 23339 5355
rect 24133 5321 24167 5355
rect 26709 5321 26743 5355
rect 30113 5321 30147 5355
rect 23029 5253 23063 5287
rect 25881 5253 25915 5287
rect 30481 5253 30515 5287
rect 4997 5185 5031 5219
rect 5089 5185 5123 5219
rect 7205 5185 7239 5219
rect 8125 5185 8159 5219
rect 10425 5185 10459 5219
rect 11161 5185 11195 5219
rect 11529 5185 11563 5219
rect 11805 5185 11839 5219
rect 15393 5185 15427 5219
rect 16865 5185 16899 5219
rect 20085 5185 20119 5219
rect 21097 5185 21131 5219
rect 24777 5185 24811 5219
rect 25329 5185 25363 5219
rect 26341 5185 26375 5219
rect 28181 5185 28215 5219
rect 28457 5185 28491 5219
rect 31769 5185 31803 5219
rect 33793 5185 33827 5219
rect 4445 5117 4479 5151
rect 7665 5117 7699 5151
rect 8217 5117 8251 5151
rect 13461 5117 13495 5151
rect 14197 5117 14231 5151
rect 14657 5117 14691 5151
rect 15301 5117 15335 5151
rect 16681 5117 16715 5151
rect 17969 5117 18003 5151
rect 18521 5117 18555 5151
rect 19073 5117 19107 5151
rect 23673 5117 23707 5151
rect 25513 5117 25547 5151
rect 29101 5117 29135 5151
rect 29837 5117 29871 5151
rect 30205 5117 30239 5151
rect 32137 5117 32171 5151
rect 32597 5117 32631 5151
rect 3249 5049 3283 5083
rect 4905 5049 4939 5083
rect 6929 5049 6963 5083
rect 7573 5049 7607 5083
rect 8493 5049 8527 5083
rect 8585 5049 8619 5083
rect 10149 5049 10183 5083
rect 14565 5049 14599 5083
rect 15209 5049 15243 5083
rect 4537 4981 4571 5015
rect 5457 4981 5491 5015
rect 7757 4981 7791 5015
rect 8677 4981 8711 5015
rect 10609 4981 10643 5015
rect 13277 4981 13311 5015
rect 16313 4981 16347 5015
rect 16773 4981 16807 5015
rect 17325 4981 17359 5015
rect 19165 4981 19199 5015
rect 23765 4981 23799 5015
rect 25421 4981 25455 5015
rect 28549 4981 28583 5015
rect 29285 4981 29319 5015
rect 31217 4981 31251 5015
rect 32045 4981 32079 5015
rect 3341 4777 3375 4811
rect 5457 4777 5491 4811
rect 6561 4777 6595 4811
rect 6929 4777 6963 4811
rect 10701 4777 10735 4811
rect 11897 4777 11931 4811
rect 12265 4777 12299 4811
rect 20085 4777 20119 4811
rect 27169 4777 27203 4811
rect 28181 4777 28215 4811
rect 28641 4777 28675 4811
rect 29009 4777 29043 4811
rect 29101 4777 29135 4811
rect 31861 4777 31895 4811
rect 5273 4709 5307 4743
rect 5733 4709 5767 4743
rect 16313 4709 16347 4743
rect 17969 4709 18003 4743
rect 23121 4709 23155 4743
rect 30389 4709 30423 4743
rect 3065 4641 3099 4675
rect 5365 4641 5399 4675
rect 5641 4641 5675 4675
rect 5825 4641 5859 4675
rect 6009 4641 6043 4675
rect 6469 4641 6503 4675
rect 7205 4641 7239 4675
rect 9781 4641 9815 4675
rect 10793 4641 10827 4675
rect 12909 4641 12943 4675
rect 16037 4641 16071 4675
rect 18061 4641 18095 4675
rect 18337 4641 18371 4675
rect 22201 4641 22235 4675
rect 23213 4641 23247 4675
rect 25237 4641 25271 4675
rect 25329 4641 25363 4675
rect 29653 4641 29687 4675
rect 32229 4641 32263 4675
rect 4813 4573 4847 4607
rect 5089 4573 5123 4607
rect 6377 4573 6411 4607
rect 9505 4573 9539 4607
rect 13369 4573 13403 4607
rect 13645 4573 13679 4607
rect 15117 4573 15151 4607
rect 15853 4573 15887 4607
rect 18613 4573 18647 4607
rect 21925 4573 21959 4607
rect 22293 4573 22327 4607
rect 22845 4573 22879 4607
rect 24961 4573 24995 4607
rect 25605 4573 25639 4607
rect 27721 4573 27755 4607
rect 29193 4573 29227 4607
rect 30113 4573 30147 4607
rect 33425 4573 33459 4607
rect 8033 4505 8067 4539
rect 29929 4505 29963 4539
rect 3249 4437 3283 4471
rect 7849 4437 7883 4471
rect 15209 4437 15243 4471
rect 17785 4437 17819 4471
rect 20453 4437 20487 4471
rect 23489 4437 23523 4471
rect 27077 4437 27111 4471
rect 29561 4437 29595 4471
rect 5181 4233 5215 4267
rect 5733 4233 5767 4267
rect 6101 4233 6135 4267
rect 6837 4233 6871 4267
rect 9597 4233 9631 4267
rect 13737 4233 13771 4267
rect 15301 4233 15335 4267
rect 16221 4233 16255 4267
rect 18429 4233 18463 4267
rect 24869 4233 24903 4267
rect 26065 4233 26099 4267
rect 26893 4233 26927 4267
rect 29469 4233 29503 4267
rect 6561 4165 6595 4199
rect 16497 4165 16531 4199
rect 18245 4165 18279 4199
rect 4537 4097 4571 4131
rect 8309 4097 8343 4131
rect 8401 4097 8435 4131
rect 13185 4097 13219 4131
rect 14289 4097 14323 4131
rect 14749 4097 14783 4131
rect 18981 4097 19015 4131
rect 20085 4097 20119 4131
rect 20729 4097 20763 4131
rect 21097 4097 21131 4131
rect 21189 4097 21223 4131
rect 23305 4097 23339 4131
rect 23581 4097 23615 4131
rect 25513 4097 25547 4131
rect 26617 4097 26651 4131
rect 27721 4097 27755 4131
rect 27997 4097 28031 4131
rect 4445 4029 4479 4063
rect 8493 4029 8527 4063
rect 8953 4029 8987 4063
rect 14105 4029 14139 4063
rect 14197 4029 14231 4063
rect 15393 4029 15427 4063
rect 18797 4029 18831 4063
rect 21281 4029 21315 4063
rect 23765 4029 23799 4063
rect 24225 4029 24259 4063
rect 26985 4029 27019 4063
rect 33701 4029 33735 4063
rect 33977 4029 34011 4063
rect 3249 3961 3283 3995
rect 8861 3893 8895 3927
rect 18889 3893 18923 3927
rect 19533 3893 19567 3927
rect 21649 3893 21683 3927
rect 23673 3893 23707 3927
rect 24133 3893 24167 3927
rect 33517 3893 33551 3927
rect 33793 3893 33827 3927
rect 9045 3689 9079 3723
rect 14657 3689 14691 3723
rect 25973 3689 26007 3723
rect 28917 3689 28951 3723
rect 4445 3553 4479 3587
rect 6653 3553 6687 3587
rect 16405 3553 16439 3587
rect 20729 3553 20763 3587
rect 32321 3553 32355 3587
rect 33977 3553 34011 3587
rect 3249 3485 3283 3519
rect 5457 3485 5491 3519
rect 16681 3485 16715 3519
rect 21189 3485 21223 3519
rect 33057 3485 33091 3519
rect 33793 3417 33827 3451
rect 9689 3145 9723 3179
rect 11253 3145 11287 3179
rect 23673 3145 23707 3179
rect 26065 3145 26099 3179
rect 28641 3145 28675 3179
rect 31677 3145 31711 3179
rect 3249 3077 3283 3111
rect 13829 3077 13863 3111
rect 5457 3009 5491 3043
rect 5733 3009 5767 3043
rect 8493 3009 8527 3043
rect 12265 3009 12299 3043
rect 14841 3009 14875 3043
rect 17417 3009 17451 3043
rect 19257 3009 19291 3043
rect 22385 3009 22419 3043
rect 24961 3009 24995 3043
rect 27537 3009 27571 3043
rect 30113 3009 30147 3043
rect 32873 3009 32907 3043
rect 3065 2941 3099 2975
rect 5273 2941 5307 2975
rect 7849 2941 7883 2975
rect 8033 2941 8067 2975
rect 9505 2941 9539 2975
rect 11069 2941 11103 2975
rect 13001 2941 13035 2975
rect 13645 2941 13679 2975
rect 14197 2941 14231 2975
rect 16773 2941 16807 2975
rect 18797 2941 18831 2975
rect 21925 2941 21959 2975
rect 23489 2941 23523 2975
rect 24501 2941 24535 2975
rect 26249 2941 26283 2975
rect 27077 2941 27111 2975
rect 28825 2941 28859 2975
rect 29837 2941 29871 2975
rect 31861 2941 31895 2975
rect 32229 2941 32263 2975
rect 33977 2941 34011 2975
rect 4077 2873 4111 2907
rect 6653 2873 6687 2907
rect 33793 2805 33827 2839
<< metal1 >>
rect 2760 34298 34316 34320
rect 2760 34246 7210 34298
rect 7262 34246 7274 34298
rect 7326 34246 7338 34298
rect 7390 34246 7402 34298
rect 7454 34246 7466 34298
rect 7518 34246 15099 34298
rect 15151 34246 15163 34298
rect 15215 34246 15227 34298
rect 15279 34246 15291 34298
rect 15343 34246 15355 34298
rect 15407 34246 22988 34298
rect 23040 34246 23052 34298
rect 23104 34246 23116 34298
rect 23168 34246 23180 34298
rect 23232 34246 23244 34298
rect 23296 34246 30877 34298
rect 30929 34246 30941 34298
rect 30993 34246 31005 34298
rect 31057 34246 31069 34298
rect 31121 34246 31133 34298
rect 31185 34246 34316 34298
rect 2760 34224 34316 34246
rect 7742 34144 7748 34196
rect 7800 34144 7806 34196
rect 15470 34144 15476 34196
rect 15528 34144 15534 34196
rect 22554 34144 22560 34196
rect 22612 34144 22618 34196
rect 4341 34119 4399 34125
rect 4341 34085 4353 34119
rect 4387 34116 4399 34119
rect 4522 34116 4528 34128
rect 4387 34088 4528 34116
rect 4387 34085 4399 34088
rect 4341 34079 4399 34085
rect 4522 34076 4528 34088
rect 4580 34076 4586 34128
rect 5810 34076 5816 34128
rect 5868 34076 5874 34128
rect 3050 34008 3056 34060
rect 3108 34008 3114 34060
rect 4706 34008 4712 34060
rect 4764 34048 4770 34060
rect 5077 34051 5135 34057
rect 5077 34048 5089 34051
rect 4764 34020 5089 34048
rect 4764 34008 4770 34020
rect 5077 34017 5089 34020
rect 5123 34017 5135 34051
rect 5077 34011 5135 34017
rect 5828 33980 5856 34076
rect 5994 34008 6000 34060
rect 6052 34008 6058 34060
rect 7760 34048 7788 34144
rect 12894 34076 12900 34128
rect 12952 34116 12958 34128
rect 14093 34119 14151 34125
rect 14093 34116 14105 34119
rect 12952 34088 14105 34116
rect 12952 34076 12958 34088
rect 14093 34085 14105 34088
rect 14139 34085 14151 34119
rect 15488 34116 15516 34144
rect 15488 34088 15792 34116
rect 14093 34079 14151 34085
rect 8021 34051 8079 34057
rect 8021 34048 8033 34051
rect 7760 34020 8033 34048
rect 8021 34017 8033 34020
rect 8067 34017 8079 34051
rect 8021 34011 8079 34017
rect 9033 34051 9091 34057
rect 9033 34017 9045 34051
rect 9079 34017 9091 34051
rect 9033 34011 9091 34017
rect 6365 33983 6423 33989
rect 6365 33980 6377 33983
rect 5828 33952 6377 33980
rect 6365 33949 6377 33952
rect 6411 33949 6423 33983
rect 9048 33980 9076 34011
rect 9122 34008 9128 34060
rect 9180 34048 9186 34060
rect 9180 34020 9720 34048
rect 9180 34008 9186 34020
rect 9214 33980 9220 33992
rect 9048 33952 9220 33980
rect 6365 33943 6423 33949
rect 9214 33940 9220 33952
rect 9272 33940 9278 33992
rect 9692 33989 9720 34020
rect 10318 34008 10324 34060
rect 10376 34048 10382 34060
rect 10597 34051 10655 34057
rect 10597 34048 10609 34051
rect 10376 34020 10609 34048
rect 10376 34008 10382 34020
rect 10597 34017 10609 34020
rect 10643 34017 10655 34051
rect 12529 34051 12587 34057
rect 12529 34048 12541 34051
rect 10597 34011 10655 34017
rect 12406 34020 12541 34048
rect 9677 33983 9735 33989
rect 9677 33949 9689 33983
rect 9723 33949 9735 33983
rect 9677 33943 9735 33949
rect 10870 33940 10876 33992
rect 10928 33940 10934 33992
rect 11698 33940 11704 33992
rect 11756 33940 11762 33992
rect 10594 33872 10600 33924
rect 10652 33912 10658 33924
rect 12406 33912 12434 34020
rect 12529 34017 12541 34020
rect 12575 34048 12587 34051
rect 12618 34048 12624 34060
rect 12575 34020 12624 34048
rect 12575 34017 12587 34020
rect 12529 34011 12587 34017
rect 12618 34008 12624 34020
rect 12676 34008 12682 34060
rect 13354 34008 13360 34060
rect 13412 34008 13418 34060
rect 14182 34008 14188 34060
rect 14240 34048 14246 34060
rect 15764 34057 15792 34088
rect 19978 34076 19984 34128
rect 20036 34116 20042 34128
rect 21085 34119 21143 34125
rect 21085 34116 21097 34119
rect 20036 34088 21097 34116
rect 20036 34076 20042 34088
rect 21085 34085 21097 34088
rect 21131 34085 21143 34119
rect 21085 34079 21143 34085
rect 15565 34051 15623 34057
rect 15565 34048 15577 34051
rect 14240 34020 15577 34048
rect 14240 34008 14246 34020
rect 15565 34017 15577 34020
rect 15611 34017 15623 34051
rect 15565 34011 15623 34017
rect 15749 34051 15807 34057
rect 15749 34017 15761 34051
rect 15795 34017 15807 34051
rect 15749 34011 15807 34017
rect 18414 34008 18420 34060
rect 18472 34008 18478 34060
rect 22094 34008 22100 34060
rect 22152 34008 22158 34060
rect 22572 34048 22600 34144
rect 23842 34076 23848 34128
rect 23900 34076 23906 34128
rect 28350 34076 28356 34128
rect 28408 34116 28414 34128
rect 28813 34119 28871 34125
rect 28813 34116 28825 34119
rect 28408 34088 28825 34116
rect 28408 34076 28414 34088
rect 28813 34085 28825 34088
rect 28859 34085 28871 34119
rect 28813 34079 28871 34085
rect 22649 34051 22707 34057
rect 22649 34048 22661 34051
rect 22572 34020 22661 34048
rect 22649 34017 22661 34020
rect 22695 34017 22707 34051
rect 22649 34011 22707 34017
rect 15194 33940 15200 33992
rect 15252 33940 15258 33992
rect 17402 33940 17408 33992
rect 17460 33980 17466 33992
rect 18785 33983 18843 33989
rect 18785 33980 18797 33983
rect 17460 33952 18797 33980
rect 17460 33940 17466 33952
rect 18785 33949 18797 33952
rect 18831 33949 18843 33983
rect 23860 33980 23888 34076
rect 24118 34008 24124 34060
rect 24176 34008 24182 34060
rect 26050 34008 26056 34060
rect 26108 34008 26114 34060
rect 30006 34008 30012 34060
rect 30064 34008 30070 34060
rect 31202 34008 31208 34060
rect 31260 34008 31266 34060
rect 24397 33983 24455 33989
rect 24397 33980 24409 33983
rect 23860 33952 24409 33980
rect 18785 33943 18843 33949
rect 24397 33949 24409 33952
rect 24443 33949 24455 33983
rect 24397 33943 24455 33949
rect 25130 33940 25136 33992
rect 25188 33980 25194 33992
rect 26513 33983 26571 33989
rect 26513 33980 26525 33983
rect 25188 33952 26525 33980
rect 25188 33940 25194 33952
rect 26513 33949 26525 33952
rect 26559 33949 26571 33983
rect 26513 33943 26571 33949
rect 29638 33940 29644 33992
rect 29696 33980 29702 33992
rect 31757 33983 31815 33989
rect 31757 33980 31769 33983
rect 29696 33952 31769 33980
rect 29696 33940 29702 33952
rect 31757 33949 31769 33952
rect 31803 33949 31815 33983
rect 31757 33943 31815 33949
rect 10652 33884 12434 33912
rect 10652 33872 10658 33884
rect 3237 33847 3295 33853
rect 3237 33813 3249 33847
rect 3283 33844 3295 33847
rect 5534 33844 5540 33856
rect 3283 33816 5540 33844
rect 3283 33813 3295 33816
rect 3237 33807 3295 33813
rect 5534 33804 5540 33816
rect 5592 33804 5598 33856
rect 8202 33804 8208 33856
rect 8260 33804 8266 33856
rect 12250 33804 12256 33856
rect 12308 33804 12314 33856
rect 12434 33804 12440 33856
rect 12492 33804 12498 33856
rect 14182 33804 14188 33856
rect 14240 33844 14246 33856
rect 14645 33847 14703 33853
rect 14645 33844 14657 33847
rect 14240 33816 14657 33844
rect 14240 33804 14246 33816
rect 14645 33813 14657 33816
rect 14691 33813 14703 33847
rect 14645 33807 14703 33813
rect 15381 33847 15439 33853
rect 15381 33813 15393 33847
rect 15427 33844 15439 33847
rect 15746 33844 15752 33856
rect 15427 33816 15752 33844
rect 15427 33813 15439 33816
rect 15381 33807 15439 33813
rect 15746 33804 15752 33816
rect 15804 33804 15810 33856
rect 15933 33847 15991 33853
rect 15933 33813 15945 33847
rect 15979 33844 15991 33847
rect 16942 33844 16948 33856
rect 15979 33816 16948 33844
rect 15979 33813 15991 33816
rect 15933 33807 15991 33813
rect 16942 33804 16948 33816
rect 17000 33804 17006 33856
rect 22830 33804 22836 33856
rect 22888 33804 22894 33856
rect 2760 33754 34316 33776
rect 2760 33702 6550 33754
rect 6602 33702 6614 33754
rect 6666 33702 6678 33754
rect 6730 33702 6742 33754
rect 6794 33702 6806 33754
rect 6858 33702 14439 33754
rect 14491 33702 14503 33754
rect 14555 33702 14567 33754
rect 14619 33702 14631 33754
rect 14683 33702 14695 33754
rect 14747 33702 22328 33754
rect 22380 33702 22392 33754
rect 22444 33702 22456 33754
rect 22508 33702 22520 33754
rect 22572 33702 22584 33754
rect 22636 33702 30217 33754
rect 30269 33702 30281 33754
rect 30333 33702 30345 33754
rect 30397 33702 30409 33754
rect 30461 33702 30473 33754
rect 30525 33702 34316 33754
rect 2760 33680 34316 33702
rect 12618 33600 12624 33652
rect 12676 33640 12682 33652
rect 33042 33640 33048 33652
rect 12676 33612 15608 33640
rect 12676 33600 12682 33612
rect 3234 33464 3240 33516
rect 3292 33504 3298 33516
rect 3513 33507 3571 33513
rect 3513 33504 3525 33507
rect 3292 33476 3525 33504
rect 3292 33464 3298 33476
rect 3513 33473 3525 33476
rect 3559 33473 3571 33507
rect 3513 33467 3571 33473
rect 5902 33464 5908 33516
rect 5960 33464 5966 33516
rect 12250 33464 12256 33516
rect 12308 33504 12314 33516
rect 12713 33507 12771 33513
rect 12713 33504 12725 33507
rect 12308 33476 12725 33504
rect 12308 33464 12314 33476
rect 12713 33473 12725 33476
rect 12759 33473 12771 33507
rect 12713 33467 12771 33473
rect 13817 33507 13875 33513
rect 13817 33473 13829 33507
rect 13863 33504 13875 33507
rect 14182 33504 14188 33516
rect 13863 33476 14188 33504
rect 13863 33473 13875 33476
rect 13817 33467 13875 33473
rect 14182 33464 14188 33476
rect 14240 33464 14246 33516
rect 4709 33439 4767 33445
rect 4709 33405 4721 33439
rect 4755 33436 4767 33439
rect 4755 33408 5120 33436
rect 4755 33405 4767 33408
rect 4709 33399 4767 33405
rect 5092 33309 5120 33408
rect 5442 33396 5448 33448
rect 5500 33396 5506 33448
rect 7926 33396 7932 33448
rect 7984 33436 7990 33448
rect 8665 33439 8723 33445
rect 8665 33436 8677 33439
rect 7984 33408 8677 33436
rect 7984 33396 7990 33408
rect 8665 33405 8677 33408
rect 8711 33405 8723 33439
rect 8665 33399 8723 33405
rect 10778 33396 10784 33448
rect 10836 33396 10842 33448
rect 15580 33445 15608 33612
rect 30392 33612 33048 33640
rect 19702 33504 19708 33516
rect 18800 33476 19708 33504
rect 12989 33439 13047 33445
rect 12989 33405 13001 33439
rect 13035 33436 13047 33439
rect 13541 33439 13599 33445
rect 13541 33436 13553 33439
rect 13035 33408 13553 33436
rect 13035 33405 13047 33408
rect 12989 33399 13047 33405
rect 13541 33405 13553 33408
rect 13587 33405 13599 33439
rect 13541 33399 13599 33405
rect 15565 33439 15623 33445
rect 15565 33405 15577 33439
rect 15611 33405 15623 33439
rect 15565 33399 15623 33405
rect 8938 33328 8944 33380
rect 8996 33328 9002 33380
rect 10689 33371 10747 33377
rect 10689 33368 10701 33371
rect 10166 33340 10701 33368
rect 10689 33337 10701 33340
rect 10735 33337 10747 33371
rect 12434 33368 12440 33380
rect 12282 33340 12440 33368
rect 10689 33331 10747 33337
rect 12434 33328 12440 33340
rect 12492 33328 12498 33380
rect 13078 33328 13084 33380
rect 13136 33328 13142 33380
rect 13265 33371 13323 33377
rect 13265 33337 13277 33371
rect 13311 33368 13323 33371
rect 13354 33368 13360 33380
rect 13311 33340 13360 33368
rect 13311 33337 13323 33340
rect 13265 33331 13323 33337
rect 13354 33328 13360 33340
rect 13412 33328 13418 33380
rect 13556 33368 13584 33399
rect 18690 33396 18696 33448
rect 18748 33396 18754 33448
rect 18800 33445 18828 33476
rect 19702 33464 19708 33476
rect 19760 33464 19766 33516
rect 26418 33464 26424 33516
rect 26476 33504 26482 33516
rect 26973 33507 27031 33513
rect 26973 33504 26985 33507
rect 26476 33476 26985 33504
rect 26476 33464 26482 33476
rect 26973 33473 26985 33476
rect 27019 33473 27031 33507
rect 26973 33467 27031 33473
rect 30285 33507 30343 33513
rect 30285 33473 30297 33507
rect 30331 33504 30343 33507
rect 30392 33504 30420 33612
rect 33042 33600 33048 33612
rect 33100 33600 33106 33652
rect 30331 33476 30420 33504
rect 30331 33473 30343 33476
rect 30285 33467 30343 33473
rect 31294 33464 31300 33516
rect 31352 33504 31358 33516
rect 31757 33507 31815 33513
rect 31757 33504 31769 33507
rect 31352 33476 31769 33504
rect 31352 33464 31358 33476
rect 31757 33473 31769 33476
rect 31803 33473 31815 33507
rect 31757 33467 31815 33473
rect 18785 33439 18843 33445
rect 18785 33405 18797 33439
rect 18831 33405 18843 33439
rect 18785 33399 18843 33405
rect 18877 33439 18935 33445
rect 18877 33405 18889 33439
rect 18923 33405 18935 33439
rect 18877 33399 18935 33405
rect 14090 33368 14096 33380
rect 13556 33340 14096 33368
rect 14090 33328 14096 33340
rect 14148 33328 14154 33380
rect 15473 33371 15531 33377
rect 15473 33368 15485 33371
rect 15042 33340 15485 33368
rect 15473 33337 15485 33340
rect 15519 33337 15531 33371
rect 18708 33368 18736 33396
rect 18892 33368 18920 33399
rect 21266 33396 21272 33448
rect 21324 33436 21330 33448
rect 21361 33439 21419 33445
rect 21361 33436 21373 33439
rect 21324 33408 21373 33436
rect 21324 33396 21330 33408
rect 21361 33405 21373 33408
rect 21407 33405 21419 33439
rect 21361 33399 21419 33405
rect 26510 33396 26516 33448
rect 26568 33396 26574 33448
rect 31021 33439 31079 33445
rect 31021 33405 31033 33439
rect 31067 33405 31079 33439
rect 31021 33399 31079 33405
rect 18708 33340 18920 33368
rect 31036 33368 31064 33399
rect 31386 33396 31392 33448
rect 31444 33396 31450 33448
rect 32674 33368 32680 33380
rect 31036 33340 32680 33368
rect 15473 33331 15531 33337
rect 32674 33328 32680 33340
rect 32732 33328 32738 33380
rect 5077 33303 5135 33309
rect 5077 33269 5089 33303
rect 5123 33300 5135 33303
rect 5166 33300 5172 33312
rect 5123 33272 5172 33300
rect 5123 33269 5135 33272
rect 5077 33263 5135 33269
rect 5166 33260 5172 33272
rect 5224 33260 5230 33312
rect 10413 33303 10471 33309
rect 10413 33269 10425 33303
rect 10459 33300 10471 33303
rect 11054 33300 11060 33312
rect 10459 33272 11060 33300
rect 10459 33269 10471 33272
rect 10413 33263 10471 33269
rect 11054 33260 11060 33272
rect 11112 33260 11118 33312
rect 11241 33303 11299 33309
rect 11241 33269 11253 33303
rect 11287 33300 11299 33303
rect 12526 33300 12532 33312
rect 11287 33272 12532 33300
rect 11287 33269 11299 33272
rect 11241 33263 11299 33269
rect 12526 33260 12532 33272
rect 12584 33260 12590 33312
rect 15289 33303 15347 33309
rect 15289 33269 15301 33303
rect 15335 33300 15347 33303
rect 15378 33300 15384 33312
rect 15335 33272 15384 33300
rect 15335 33269 15347 33272
rect 15289 33263 15347 33269
rect 15378 33260 15384 33272
rect 15436 33260 15442 33312
rect 18598 33260 18604 33312
rect 18656 33300 18662 33312
rect 18693 33303 18751 33309
rect 18693 33300 18705 33303
rect 18656 33272 18705 33300
rect 18656 33260 18662 33272
rect 18693 33269 18705 33272
rect 18739 33269 18751 33303
rect 18693 33263 18751 33269
rect 19058 33260 19064 33312
rect 19116 33260 19122 33312
rect 21542 33260 21548 33312
rect 21600 33260 21606 33312
rect 2760 33210 34316 33232
rect 2760 33158 7210 33210
rect 7262 33158 7274 33210
rect 7326 33158 7338 33210
rect 7390 33158 7402 33210
rect 7454 33158 7466 33210
rect 7518 33158 15099 33210
rect 15151 33158 15163 33210
rect 15215 33158 15227 33210
rect 15279 33158 15291 33210
rect 15343 33158 15355 33210
rect 15407 33158 22988 33210
rect 23040 33158 23052 33210
rect 23104 33158 23116 33210
rect 23168 33158 23180 33210
rect 23232 33158 23244 33210
rect 23296 33158 30877 33210
rect 30929 33158 30941 33210
rect 30993 33158 31005 33210
rect 31057 33158 31069 33210
rect 31121 33158 31133 33210
rect 31185 33158 34316 33210
rect 2760 33136 34316 33158
rect 1946 33056 1952 33108
rect 2004 33096 2010 33108
rect 5902 33096 5908 33108
rect 2004 33068 5908 33096
rect 2004 33056 2010 33068
rect 5902 33056 5908 33068
rect 5960 33056 5966 33108
rect 8938 33056 8944 33108
rect 8996 33096 9002 33108
rect 9033 33099 9091 33105
rect 9033 33096 9045 33099
rect 8996 33068 9045 33096
rect 8996 33056 9002 33068
rect 9033 33065 9045 33068
rect 9079 33065 9091 33099
rect 11422 33096 11428 33108
rect 9033 33059 9091 33065
rect 9140 33068 11428 33096
rect 3234 32988 3240 33040
rect 3292 32988 3298 33040
rect 3786 32988 3792 33040
rect 3844 33028 3850 33040
rect 4709 33031 4767 33037
rect 4709 33028 4721 33031
rect 3844 33000 4721 33028
rect 3844 32988 3850 33000
rect 4709 32997 4721 33000
rect 4755 32997 4767 33031
rect 9140 33028 9168 33068
rect 11422 33056 11428 33068
rect 11480 33056 11486 33108
rect 11609 33099 11667 33105
rect 11609 33065 11621 33099
rect 11655 33096 11667 33099
rect 11698 33096 11704 33108
rect 11655 33068 11704 33096
rect 11655 33065 11667 33068
rect 11609 33059 11667 33065
rect 11698 33056 11704 33068
rect 11756 33056 11762 33108
rect 12526 33096 12532 33108
rect 12452 33068 12532 33096
rect 4709 32991 4767 32997
rect 5644 33000 9168 33028
rect 10137 33031 10195 33037
rect 4433 32963 4491 32969
rect 4433 32929 4445 32963
rect 4479 32960 4491 32963
rect 5644 32960 5672 33000
rect 10137 32997 10149 33031
rect 10183 33028 10195 33031
rect 11333 33031 11391 33037
rect 11333 33028 11345 33031
rect 10183 33000 11345 33028
rect 10183 32997 10195 33000
rect 10137 32991 10195 32997
rect 11333 32997 11345 33000
rect 11379 32997 11391 33031
rect 11333 32991 11391 32997
rect 11882 32988 11888 33040
rect 11940 32988 11946 33040
rect 4479 32932 5672 32960
rect 4479 32929 4491 32932
rect 4433 32923 4491 32929
rect 5718 32920 5724 32972
rect 5776 32920 5782 32972
rect 6917 32963 6975 32969
rect 6917 32929 6929 32963
rect 6963 32960 6975 32963
rect 7282 32960 7288 32972
rect 6963 32932 7288 32960
rect 6963 32929 6975 32932
rect 6917 32923 6975 32929
rect 7282 32920 7288 32932
rect 7340 32920 7346 32972
rect 9953 32963 10011 32969
rect 9953 32929 9965 32963
rect 9999 32929 10011 32963
rect 9953 32923 10011 32929
rect 6181 32895 6239 32901
rect 6181 32861 6193 32895
rect 6227 32861 6239 32895
rect 6181 32855 6239 32861
rect 9677 32895 9735 32901
rect 9677 32861 9689 32895
rect 9723 32892 9735 32895
rect 9769 32895 9827 32901
rect 9769 32892 9781 32895
rect 9723 32864 9781 32892
rect 9723 32861 9735 32864
rect 9677 32855 9735 32861
rect 9769 32861 9781 32864
rect 9815 32861 9827 32895
rect 9968 32892 9996 32923
rect 10042 32920 10048 32972
rect 10100 32920 10106 32972
rect 10275 32963 10333 32969
rect 10275 32929 10287 32963
rect 10321 32960 10333 32963
rect 10962 32960 10968 32972
rect 10321 32932 10968 32960
rect 10321 32929 10333 32932
rect 10275 32923 10333 32929
rect 10962 32920 10968 32932
rect 11020 32920 11026 32972
rect 11054 32920 11060 32972
rect 11112 32960 11118 32972
rect 11149 32963 11207 32969
rect 11149 32960 11161 32963
rect 11112 32932 11161 32960
rect 11112 32920 11118 32932
rect 11149 32929 11161 32932
rect 11195 32929 11207 32963
rect 11149 32923 11207 32929
rect 11241 32963 11299 32969
rect 11241 32929 11253 32963
rect 11287 32929 11299 32963
rect 11241 32923 11299 32929
rect 11425 32963 11483 32969
rect 11425 32929 11437 32963
rect 11471 32960 11483 32963
rect 11471 32932 11744 32960
rect 11810 32953 11868 32959
rect 11810 32950 11822 32953
rect 11471 32929 11483 32932
rect 11425 32923 11483 32929
rect 10134 32892 10140 32904
rect 9968 32864 10140 32892
rect 9769 32855 9827 32861
rect 5350 32784 5356 32836
rect 5408 32824 5414 32836
rect 6196 32824 6224 32855
rect 10134 32852 10140 32864
rect 10192 32852 10198 32904
rect 10413 32895 10471 32901
rect 10413 32861 10425 32895
rect 10459 32892 10471 32895
rect 11256 32892 11284 32923
rect 10459 32864 11284 32892
rect 10459 32861 10471 32864
rect 10413 32855 10471 32861
rect 10594 32824 10600 32836
rect 5408 32796 10600 32824
rect 5408 32784 5414 32796
rect 10594 32784 10600 32796
rect 10652 32784 10658 32836
rect 11072 32768 11100 32864
rect 11716 32836 11744 32932
rect 11808 32919 11822 32950
rect 11856 32919 11868 32953
rect 11974 32920 11980 32972
rect 12032 32920 12038 32972
rect 12158 32969 12164 32972
rect 12115 32963 12164 32969
rect 12115 32929 12127 32963
rect 12161 32929 12164 32963
rect 12115 32923 12164 32929
rect 12158 32920 12164 32923
rect 12216 32920 12222 32972
rect 12452 32969 12480 33068
rect 12526 33056 12532 33068
rect 12584 33056 12590 33108
rect 13814 33096 13820 33108
rect 13648 33068 13820 33096
rect 13648 32969 13676 33068
rect 13814 33056 13820 33068
rect 13872 33096 13878 33108
rect 14001 33099 14059 33105
rect 14001 33096 14013 33099
rect 13872 33068 14013 33096
rect 13872 33056 13878 33068
rect 14001 33065 14013 33068
rect 14047 33065 14059 33099
rect 15010 33096 15016 33108
rect 14001 33059 14059 33065
rect 14200 33068 15016 33096
rect 14200 33028 14228 33068
rect 15010 33056 15016 33068
rect 15068 33056 15074 33108
rect 30300 33068 36124 33096
rect 30300 33037 30328 33068
rect 36096 33040 36124 33068
rect 15749 33031 15807 33037
rect 15749 33028 15761 33031
rect 13832 33000 14228 33028
rect 15120 33000 15761 33028
rect 12437 32963 12495 32969
rect 12437 32929 12449 32963
rect 12483 32929 12495 32963
rect 13357 32963 13415 32969
rect 13357 32960 13369 32963
rect 12437 32923 12495 32929
rect 13004 32932 13369 32960
rect 11808 32913 11868 32919
rect 11698 32784 11704 32836
rect 11756 32784 11762 32836
rect 11808 32824 11836 32913
rect 12250 32852 12256 32904
rect 12308 32892 12314 32904
rect 13004 32901 13032 32932
rect 13357 32929 13369 32932
rect 13403 32929 13415 32963
rect 13357 32923 13415 32929
rect 13541 32963 13599 32969
rect 13541 32929 13553 32963
rect 13587 32929 13599 32963
rect 13541 32923 13599 32929
rect 13633 32963 13691 32969
rect 13633 32929 13645 32963
rect 13679 32929 13691 32963
rect 13633 32923 13691 32929
rect 12989 32895 13047 32901
rect 12989 32892 13001 32895
rect 12308 32864 13001 32892
rect 12308 32852 12314 32864
rect 12989 32861 13001 32864
rect 13035 32861 13047 32895
rect 12989 32855 13047 32861
rect 13173 32827 13231 32833
rect 13173 32824 13185 32827
rect 11808 32796 13185 32824
rect 13173 32793 13185 32796
rect 13219 32793 13231 32827
rect 13173 32787 13231 32793
rect 7282 32716 7288 32768
rect 7340 32716 7346 32768
rect 10965 32759 11023 32765
rect 10965 32725 10977 32759
rect 11011 32756 11023 32759
rect 11054 32756 11060 32768
rect 11011 32728 11060 32756
rect 11011 32725 11023 32728
rect 10965 32719 11023 32725
rect 11054 32716 11060 32728
rect 11112 32716 11118 32768
rect 11146 32716 11152 32768
rect 11204 32756 11210 32768
rect 13556 32756 13584 32923
rect 13832 32833 13860 33000
rect 15120 32972 15148 33000
rect 15749 32997 15761 33000
rect 15795 32997 15807 33031
rect 15749 32991 15807 32997
rect 30285 33031 30343 33037
rect 30285 32997 30297 33031
rect 30331 32997 30343 33031
rect 34790 33028 34796 33040
rect 30285 32991 30343 32997
rect 31680 33000 34796 33028
rect 13998 32960 14004 32972
rect 13959 32932 14004 32960
rect 13998 32920 14004 32932
rect 14056 32920 14062 32972
rect 14090 32920 14096 32972
rect 14148 32958 14154 32972
rect 14553 32963 14611 32969
rect 14553 32960 14565 32963
rect 14200 32958 14565 32960
rect 14148 32932 14565 32958
rect 14148 32930 14228 32932
rect 14148 32920 14154 32930
rect 14553 32929 14565 32932
rect 14599 32929 14611 32963
rect 14553 32923 14611 32929
rect 14737 32963 14795 32969
rect 14737 32929 14749 32963
rect 14783 32960 14795 32963
rect 14826 32960 14832 32972
rect 14783 32932 14832 32960
rect 14783 32929 14795 32932
rect 14737 32923 14795 32929
rect 14826 32920 14832 32932
rect 14884 32920 14890 32972
rect 15102 32920 15108 32972
rect 15160 32920 15166 32972
rect 15470 32920 15476 32972
rect 15528 32920 15534 32972
rect 15562 32920 15568 32972
rect 15620 32920 15626 32972
rect 15841 32963 15899 32969
rect 15841 32929 15853 32963
rect 15887 32929 15899 32963
rect 15841 32923 15899 32929
rect 19061 32963 19119 32969
rect 19061 32929 19073 32963
rect 19107 32929 19119 32963
rect 19061 32923 19119 32929
rect 14461 32895 14519 32901
rect 14461 32861 14473 32895
rect 14507 32861 14519 32895
rect 14461 32855 14519 32861
rect 14645 32895 14703 32901
rect 14645 32861 14657 32895
rect 14691 32892 14703 32895
rect 15856 32892 15884 32923
rect 14691 32864 15884 32892
rect 14691 32861 14703 32864
rect 14645 32855 14703 32861
rect 13817 32827 13875 32833
rect 13817 32793 13829 32827
rect 13863 32793 13875 32827
rect 14476 32824 14504 32855
rect 16114 32852 16120 32904
rect 16172 32852 16178 32904
rect 18874 32852 18880 32904
rect 18932 32852 18938 32904
rect 14918 32824 14924 32836
rect 14476 32796 14924 32824
rect 13817 32787 13875 32793
rect 14918 32784 14924 32796
rect 14976 32824 14982 32836
rect 15565 32827 15623 32833
rect 15565 32824 15577 32827
rect 14976 32796 15577 32824
rect 14976 32784 14982 32796
rect 15565 32793 15577 32796
rect 15611 32793 15623 32827
rect 18049 32827 18107 32833
rect 18049 32824 18061 32827
rect 15565 32787 15623 32793
rect 16500 32796 18061 32824
rect 11204 32728 13584 32756
rect 11204 32716 11210 32728
rect 13722 32716 13728 32768
rect 13780 32756 13786 32768
rect 14274 32756 14280 32768
rect 13780 32728 14280 32756
rect 13780 32716 13786 32728
rect 14274 32716 14280 32728
rect 14332 32756 14338 32768
rect 14369 32759 14427 32765
rect 14369 32756 14381 32759
rect 14332 32728 14381 32756
rect 14332 32716 14338 32728
rect 14369 32725 14381 32728
rect 14415 32756 14427 32759
rect 14829 32759 14887 32765
rect 14829 32756 14841 32759
rect 14415 32728 14841 32756
rect 14415 32725 14427 32728
rect 14369 32719 14427 32725
rect 14829 32725 14841 32728
rect 14875 32725 14887 32759
rect 14829 32719 14887 32725
rect 15010 32716 15016 32768
rect 15068 32756 15074 32768
rect 16500 32756 16528 32796
rect 18049 32793 18061 32796
rect 18095 32824 18107 32827
rect 19076 32824 19104 32923
rect 29270 32920 29276 32972
rect 29328 32920 29334 32972
rect 31680 32901 31708 33000
rect 34790 32988 34796 33000
rect 34848 32988 34854 33040
rect 36078 32988 36084 33040
rect 36136 32988 36142 33040
rect 32125 32963 32183 32969
rect 32125 32929 32137 32963
rect 32171 32929 32183 32963
rect 32125 32923 32183 32929
rect 19337 32895 19395 32901
rect 19337 32861 19349 32895
rect 19383 32861 19395 32895
rect 19337 32855 19395 32861
rect 31665 32895 31723 32901
rect 31665 32861 31677 32895
rect 31711 32861 31723 32895
rect 32140 32892 32168 32923
rect 32306 32920 32312 32972
rect 32364 32920 32370 32972
rect 32398 32892 32404 32904
rect 32140 32864 32404 32892
rect 31665 32855 31723 32861
rect 18095 32796 19104 32824
rect 18095 32793 18107 32796
rect 18049 32787 18107 32793
rect 15068 32728 16528 32756
rect 15068 32716 15074 32728
rect 16758 32716 16764 32768
rect 16816 32716 16822 32768
rect 18322 32716 18328 32768
rect 18380 32716 18386 32768
rect 19352 32756 19380 32855
rect 32398 32852 32404 32864
rect 32456 32852 32462 32904
rect 32769 32895 32827 32901
rect 32769 32861 32781 32895
rect 32815 32861 32827 32895
rect 32769 32855 32827 32861
rect 32214 32784 32220 32836
rect 32272 32824 32278 32836
rect 32784 32824 32812 32855
rect 32272 32796 32812 32824
rect 32272 32784 32278 32796
rect 19610 32756 19616 32768
rect 19352 32728 19616 32756
rect 19610 32716 19616 32728
rect 19668 32716 19674 32768
rect 2760 32666 34316 32688
rect 2760 32614 6550 32666
rect 6602 32614 6614 32666
rect 6666 32614 6678 32666
rect 6730 32614 6742 32666
rect 6794 32614 6806 32666
rect 6858 32614 14439 32666
rect 14491 32614 14503 32666
rect 14555 32614 14567 32666
rect 14619 32614 14631 32666
rect 14683 32614 14695 32666
rect 14747 32614 22328 32666
rect 22380 32614 22392 32666
rect 22444 32614 22456 32666
rect 22508 32614 22520 32666
rect 22572 32614 22584 32666
rect 22636 32614 30217 32666
rect 30269 32614 30281 32666
rect 30333 32614 30345 32666
rect 30397 32614 30409 32666
rect 30461 32614 30473 32666
rect 30525 32614 34316 32666
rect 2760 32592 34316 32614
rect 10042 32512 10048 32564
rect 10100 32552 10106 32564
rect 10597 32555 10655 32561
rect 10597 32552 10609 32555
rect 10100 32524 10609 32552
rect 10100 32512 10106 32524
rect 10597 32521 10609 32524
rect 10643 32521 10655 32555
rect 10597 32515 10655 32521
rect 11882 32512 11888 32564
rect 11940 32552 11946 32564
rect 12437 32555 12495 32561
rect 12437 32552 12449 32555
rect 11940 32524 12449 32552
rect 11940 32512 11946 32524
rect 12437 32521 12449 32524
rect 12483 32521 12495 32555
rect 13262 32552 13268 32564
rect 12437 32515 12495 32521
rect 12544 32524 13268 32552
rect 5537 32487 5595 32493
rect 5537 32453 5549 32487
rect 5583 32453 5595 32487
rect 5537 32447 5595 32453
rect 658 32376 664 32428
rect 716 32416 722 32428
rect 3237 32419 3295 32425
rect 3237 32416 3249 32419
rect 716 32388 3249 32416
rect 716 32376 722 32388
rect 3237 32385 3249 32388
rect 3283 32385 3295 32419
rect 3237 32379 3295 32385
rect 5261 32419 5319 32425
rect 5261 32385 5273 32419
rect 5307 32416 5319 32419
rect 5552 32416 5580 32447
rect 7282 32444 7288 32496
rect 7340 32484 7346 32496
rect 12544 32484 12572 32524
rect 13262 32512 13268 32524
rect 13320 32512 13326 32564
rect 13357 32555 13415 32561
rect 13357 32521 13369 32555
rect 13403 32552 13415 32555
rect 13722 32552 13728 32564
rect 13403 32524 13728 32552
rect 13403 32521 13415 32524
rect 13357 32515 13415 32521
rect 13722 32512 13728 32524
rect 13780 32512 13786 32564
rect 14093 32555 14151 32561
rect 14093 32552 14105 32555
rect 14016 32524 14105 32552
rect 7340 32456 12572 32484
rect 7340 32444 7346 32456
rect 12802 32444 12808 32496
rect 12860 32484 12866 32496
rect 13814 32484 13820 32496
rect 12860 32456 13820 32484
rect 12860 32444 12866 32456
rect 13814 32444 13820 32456
rect 13872 32484 13878 32496
rect 13909 32487 13967 32493
rect 13909 32484 13921 32487
rect 13872 32456 13921 32484
rect 13872 32444 13878 32456
rect 13909 32453 13921 32456
rect 13955 32453 13967 32487
rect 13909 32447 13967 32453
rect 14016 32484 14044 32524
rect 14093 32521 14105 32524
rect 14139 32521 14151 32555
rect 14093 32515 14151 32521
rect 14645 32555 14703 32561
rect 14645 32521 14657 32555
rect 14691 32552 14703 32555
rect 16114 32552 16120 32564
rect 14691 32524 16120 32552
rect 14691 32521 14703 32524
rect 14645 32515 14703 32521
rect 16114 32512 16120 32524
rect 16172 32512 16178 32564
rect 16758 32512 16764 32564
rect 16816 32552 16822 32564
rect 17233 32555 17291 32561
rect 17233 32552 17245 32555
rect 16816 32524 17245 32552
rect 16816 32512 16822 32524
rect 17233 32521 17245 32524
rect 17279 32521 17291 32555
rect 26786 32552 26792 32564
rect 17233 32515 17291 32521
rect 22066 32524 26792 32552
rect 14826 32484 14832 32496
rect 14016 32456 14832 32484
rect 5307 32388 5580 32416
rect 5307 32385 5319 32388
rect 5261 32379 5319 32385
rect 5994 32376 6000 32428
rect 6052 32376 6058 32428
rect 6181 32419 6239 32425
rect 6181 32385 6193 32419
rect 6227 32416 6239 32419
rect 6454 32416 6460 32428
rect 6227 32388 6460 32416
rect 6227 32385 6239 32388
rect 6181 32379 6239 32385
rect 6454 32376 6460 32388
rect 6512 32416 6518 32428
rect 6549 32419 6607 32425
rect 6549 32416 6561 32419
rect 6512 32388 6561 32416
rect 6512 32376 6518 32388
rect 6549 32385 6561 32388
rect 6595 32385 6607 32419
rect 10778 32416 10784 32428
rect 6549 32379 6607 32385
rect 9646 32388 10784 32416
rect 4430 32308 4436 32360
rect 4488 32308 4494 32360
rect 8938 32308 8944 32360
rect 8996 32308 9002 32360
rect 9309 32351 9367 32357
rect 9309 32317 9321 32351
rect 9355 32348 9367 32351
rect 9646 32348 9674 32388
rect 10778 32376 10784 32388
rect 10836 32376 10842 32428
rect 12250 32376 12256 32428
rect 12308 32416 12314 32428
rect 12308 32388 13400 32416
rect 12308 32376 12314 32388
rect 9355 32320 9674 32348
rect 10965 32351 11023 32357
rect 9355 32317 9367 32320
rect 9309 32311 9367 32317
rect 10965 32317 10977 32351
rect 11011 32348 11023 32351
rect 11698 32348 11704 32360
rect 11011 32320 11704 32348
rect 11011 32317 11023 32320
rect 10965 32311 11023 32317
rect 11698 32308 11704 32320
rect 11756 32308 11762 32360
rect 12069 32351 12127 32357
rect 12069 32317 12081 32351
rect 12115 32317 12127 32351
rect 12069 32311 12127 32317
rect 10781 32283 10839 32289
rect 10781 32249 10793 32283
rect 10827 32280 10839 32283
rect 11054 32280 11060 32292
rect 10827 32252 11060 32280
rect 10827 32249 10839 32252
rect 10781 32243 10839 32249
rect 11054 32240 11060 32252
rect 11112 32280 11118 32292
rect 12084 32280 12112 32311
rect 12342 32308 12348 32360
rect 12400 32308 12406 32360
rect 12526 32308 12532 32360
rect 12584 32348 12590 32360
rect 12802 32348 12808 32360
rect 12584 32320 12808 32348
rect 12584 32308 12590 32320
rect 12802 32308 12808 32320
rect 12860 32308 12866 32360
rect 13372 32357 13400 32388
rect 13265 32351 13323 32357
rect 13265 32317 13277 32351
rect 13311 32317 13323 32351
rect 13265 32311 13323 32317
rect 13357 32351 13415 32357
rect 13357 32317 13369 32351
rect 13403 32317 13415 32351
rect 13357 32311 13415 32317
rect 11112 32252 12112 32280
rect 11112 32240 11118 32252
rect 4617 32215 4675 32221
rect 4617 32181 4629 32215
rect 4663 32212 4675 32215
rect 5074 32212 5080 32224
rect 4663 32184 5080 32212
rect 4663 32181 4675 32184
rect 4617 32175 4675 32181
rect 5074 32172 5080 32184
rect 5132 32172 5138 32224
rect 5902 32172 5908 32224
rect 5960 32172 5966 32224
rect 8386 32172 8392 32224
rect 8444 32172 8450 32224
rect 9217 32215 9275 32221
rect 9217 32181 9229 32215
rect 9263 32212 9275 32215
rect 9306 32212 9312 32224
rect 9263 32184 9312 32212
rect 9263 32181 9275 32184
rect 9217 32175 9275 32181
rect 9306 32172 9312 32184
rect 9364 32172 9370 32224
rect 11882 32172 11888 32224
rect 11940 32172 11946 32224
rect 12084 32212 12112 32252
rect 12897 32283 12955 32289
rect 12897 32249 12909 32283
rect 12943 32249 12955 32283
rect 13280 32280 13308 32311
rect 14016 32280 14044 32456
rect 14826 32444 14832 32456
rect 14884 32484 14890 32496
rect 15381 32487 15439 32493
rect 15381 32484 15393 32487
rect 14884 32456 15393 32484
rect 14884 32444 14890 32456
rect 15381 32453 15393 32456
rect 15427 32484 15439 32487
rect 15562 32484 15568 32496
rect 15427 32456 15568 32484
rect 15427 32453 15439 32456
rect 15381 32447 15439 32453
rect 15562 32444 15568 32456
rect 15620 32444 15626 32496
rect 19610 32444 19616 32496
rect 19668 32484 19674 32496
rect 22066 32484 22094 32524
rect 26786 32512 26792 32524
rect 26844 32512 26850 32564
rect 19668 32456 22094 32484
rect 23937 32487 23995 32493
rect 19668 32444 19674 32456
rect 23937 32453 23949 32487
rect 23983 32484 23995 32487
rect 23983 32456 24624 32484
rect 23983 32453 23995 32456
rect 23937 32447 23995 32453
rect 16574 32376 16580 32428
rect 16632 32416 16638 32428
rect 17497 32419 17555 32425
rect 17497 32416 17509 32419
rect 16632 32388 17509 32416
rect 16632 32376 16638 32388
rect 17497 32385 17509 32388
rect 17543 32416 17555 32419
rect 17589 32419 17647 32425
rect 17589 32416 17601 32419
rect 17543 32388 17601 32416
rect 17543 32385 17555 32388
rect 17497 32379 17555 32385
rect 17589 32385 17601 32388
rect 17635 32385 17647 32419
rect 17589 32379 17647 32385
rect 17865 32419 17923 32425
rect 17865 32385 17877 32419
rect 17911 32416 17923 32419
rect 18322 32416 18328 32428
rect 17911 32388 18328 32416
rect 17911 32385 17923 32388
rect 17865 32379 17923 32385
rect 18322 32376 18328 32388
rect 18380 32376 18386 32428
rect 14366 32308 14372 32360
rect 14424 32308 14430 32360
rect 14645 32351 14703 32357
rect 14645 32317 14657 32351
rect 14691 32317 14703 32351
rect 14645 32311 14703 32317
rect 13280 32252 14044 32280
rect 12897 32243 12955 32249
rect 12912 32212 12940 32243
rect 14274 32240 14280 32292
rect 14332 32240 14338 32292
rect 14660 32280 14688 32311
rect 14826 32308 14832 32360
rect 14884 32308 14890 32360
rect 14918 32308 14924 32360
rect 14976 32308 14982 32360
rect 19628 32357 19656 32444
rect 19702 32376 19708 32428
rect 19760 32376 19766 32428
rect 19794 32376 19800 32428
rect 19852 32416 19858 32428
rect 23109 32419 23167 32425
rect 23109 32416 23121 32419
rect 19852 32388 23121 32416
rect 19852 32376 19858 32388
rect 23109 32385 23121 32388
rect 23155 32416 23167 32419
rect 23293 32419 23351 32425
rect 23293 32416 23305 32419
rect 23155 32388 23305 32416
rect 23155 32385 23167 32388
rect 23109 32379 23167 32385
rect 23293 32385 23305 32388
rect 23339 32416 23351 32419
rect 24486 32416 24492 32428
rect 23339 32388 24492 32416
rect 23339 32385 23351 32388
rect 23293 32379 23351 32385
rect 24486 32376 24492 32388
rect 24544 32376 24550 32428
rect 24596 32425 24624 32456
rect 24581 32419 24639 32425
rect 24581 32385 24593 32419
rect 24627 32385 24639 32419
rect 28537 32419 28595 32425
rect 28537 32416 28549 32419
rect 24581 32379 24639 32385
rect 28276 32388 28549 32416
rect 15565 32351 15623 32357
rect 15565 32317 15577 32351
rect 15611 32348 15623 32351
rect 19613 32351 19671 32357
rect 15611 32320 15792 32348
rect 15611 32317 15623 32320
rect 15565 32311 15623 32317
rect 14936 32280 14964 32308
rect 14660 32252 14964 32280
rect 12084 32184 12940 32212
rect 13078 32172 13084 32224
rect 13136 32212 13142 32224
rect 13541 32215 13599 32221
rect 13541 32212 13553 32215
rect 13136 32184 13553 32212
rect 13136 32172 13142 32184
rect 13541 32181 13553 32184
rect 13587 32181 13599 32215
rect 13541 32175 13599 32181
rect 14090 32172 14096 32224
rect 14148 32172 14154 32224
rect 14182 32172 14188 32224
rect 14240 32212 14246 32224
rect 15654 32212 15660 32224
rect 14240 32184 15660 32212
rect 14240 32172 14246 32184
rect 15654 32172 15660 32184
rect 15712 32172 15718 32224
rect 15764 32221 15792 32320
rect 19613 32317 19625 32351
rect 19659 32317 19671 32351
rect 19720 32348 19748 32376
rect 19981 32351 20039 32357
rect 19981 32348 19993 32351
rect 19720 32320 19993 32348
rect 19613 32311 19671 32317
rect 19981 32317 19993 32320
rect 20027 32348 20039 32351
rect 24949 32351 25007 32357
rect 24949 32348 24961 32351
rect 20027 32320 24961 32348
rect 20027 32317 20039 32320
rect 19981 32311 20039 32317
rect 24949 32317 24961 32320
rect 24995 32317 25007 32351
rect 24949 32311 25007 32317
rect 15930 32240 15936 32292
rect 15988 32280 15994 32292
rect 15988 32252 16054 32280
rect 15988 32240 15994 32252
rect 18598 32240 18604 32292
rect 18656 32240 18662 32292
rect 23477 32283 23535 32289
rect 23477 32249 23489 32283
rect 23523 32280 23535 32283
rect 23523 32252 25268 32280
rect 23523 32249 23535 32252
rect 23477 32243 23535 32249
rect 25240 32224 25268 32252
rect 28276 32224 28304 32388
rect 28537 32385 28549 32388
rect 28583 32385 28595 32419
rect 28537 32379 28595 32385
rect 30285 32419 30343 32425
rect 30285 32385 30297 32419
rect 30331 32416 30343 32419
rect 30374 32416 30380 32428
rect 30331 32388 30380 32416
rect 30331 32385 30343 32388
rect 30285 32379 30343 32385
rect 30374 32376 30380 32388
rect 30432 32416 30438 32428
rect 31202 32416 31208 32428
rect 30432 32388 31208 32416
rect 30432 32376 30438 32388
rect 31202 32376 31208 32388
rect 31260 32376 31266 32428
rect 33781 32419 33839 32425
rect 33781 32385 33793 32419
rect 33827 32416 33839 32419
rect 34882 32416 34888 32428
rect 33827 32388 34888 32416
rect 33827 32385 33839 32388
rect 33781 32379 33839 32385
rect 34882 32376 34888 32388
rect 34940 32376 34946 32428
rect 32769 32351 32827 32357
rect 32769 32317 32781 32351
rect 32815 32348 32827 32351
rect 33042 32348 33048 32360
rect 32815 32320 33048 32348
rect 32815 32317 32827 32320
rect 32769 32311 32827 32317
rect 33042 32308 33048 32320
rect 33100 32308 33106 32360
rect 28721 32283 28779 32289
rect 28721 32249 28733 32283
rect 28767 32280 28779 32283
rect 29641 32283 29699 32289
rect 29641 32280 29653 32283
rect 28767 32252 29653 32280
rect 28767 32249 28779 32252
rect 28721 32243 28779 32249
rect 29641 32249 29653 32252
rect 29687 32249 29699 32283
rect 29641 32243 29699 32249
rect 15749 32215 15807 32221
rect 15749 32181 15761 32215
rect 15795 32181 15807 32215
rect 15749 32175 15807 32181
rect 18782 32172 18788 32224
rect 18840 32212 18846 32224
rect 19337 32215 19395 32221
rect 19337 32212 19349 32215
rect 18840 32184 19349 32212
rect 18840 32172 18846 32184
rect 19337 32181 19349 32184
rect 19383 32181 19395 32215
rect 19337 32175 19395 32181
rect 23569 32215 23627 32221
rect 23569 32181 23581 32215
rect 23615 32212 23627 32215
rect 23842 32212 23848 32224
rect 23615 32184 23848 32212
rect 23615 32181 23627 32184
rect 23569 32175 23627 32181
rect 23842 32172 23848 32184
rect 23900 32172 23906 32224
rect 24026 32172 24032 32224
rect 24084 32172 24090 32224
rect 24854 32172 24860 32224
rect 24912 32172 24918 32224
rect 25222 32172 25228 32224
rect 25280 32172 25286 32224
rect 28258 32172 28264 32224
rect 28316 32172 28322 32224
rect 28810 32172 28816 32224
rect 28868 32172 28874 32224
rect 29178 32172 29184 32224
rect 29236 32172 29242 32224
rect 2760 32122 34316 32144
rect 2760 32070 7210 32122
rect 7262 32070 7274 32122
rect 7326 32070 7338 32122
rect 7390 32070 7402 32122
rect 7454 32070 7466 32122
rect 7518 32070 15099 32122
rect 15151 32070 15163 32122
rect 15215 32070 15227 32122
rect 15279 32070 15291 32122
rect 15343 32070 15355 32122
rect 15407 32070 22988 32122
rect 23040 32070 23052 32122
rect 23104 32070 23116 32122
rect 23168 32070 23180 32122
rect 23232 32070 23244 32122
rect 23296 32070 30877 32122
rect 30929 32070 30941 32122
rect 30993 32070 31005 32122
rect 31057 32070 31069 32122
rect 31121 32070 31133 32122
rect 31185 32070 34316 32122
rect 2760 32048 34316 32070
rect 4908 31980 7972 32008
rect 4908 31884 4936 31980
rect 5074 31900 5080 31952
rect 5132 31940 5138 31952
rect 5169 31943 5227 31949
rect 5169 31940 5181 31943
rect 5132 31912 5181 31940
rect 5132 31900 5138 31912
rect 5169 31909 5181 31912
rect 5215 31909 5227 31943
rect 6825 31943 6883 31949
rect 6825 31940 6837 31943
rect 6394 31912 6837 31940
rect 5169 31903 5227 31909
rect 6825 31909 6837 31912
rect 6871 31909 6883 31943
rect 6825 31903 6883 31909
rect 7944 31884 7972 31980
rect 9214 31968 9220 32020
rect 9272 32008 9278 32020
rect 9769 32011 9827 32017
rect 9769 32008 9781 32011
rect 9272 31980 9781 32008
rect 9272 31968 9278 31980
rect 9769 31977 9781 31980
rect 9815 31977 9827 32011
rect 9769 31971 9827 31977
rect 10134 31968 10140 32020
rect 10192 32008 10198 32020
rect 10192 31980 15424 32008
rect 10192 31968 10198 31980
rect 15396 31952 15424 31980
rect 15470 31968 15476 32020
rect 15528 32008 15534 32020
rect 15930 32008 15936 32020
rect 15528 31980 15936 32008
rect 15528 31968 15534 31980
rect 15930 31968 15936 31980
rect 15988 31968 15994 32020
rect 18325 32011 18383 32017
rect 18325 31977 18337 32011
rect 18371 32008 18383 32011
rect 18874 32008 18880 32020
rect 18371 31980 18880 32008
rect 18371 31977 18383 31980
rect 18325 31971 18383 31977
rect 18874 31968 18880 31980
rect 18932 31968 18938 32020
rect 19429 32011 19487 32017
rect 19429 31977 19441 32011
rect 19475 32008 19487 32011
rect 19794 32008 19800 32020
rect 19475 31980 19800 32008
rect 19475 31977 19487 31980
rect 19429 31971 19487 31977
rect 8297 31943 8355 31949
rect 8297 31909 8309 31943
rect 8343 31940 8355 31943
rect 8386 31940 8392 31952
rect 8343 31912 8392 31940
rect 8343 31909 8355 31912
rect 8297 31903 8355 31909
rect 8386 31900 8392 31912
rect 8444 31900 8450 31952
rect 9306 31900 9312 31952
rect 9364 31900 9370 31952
rect 11054 31900 11060 31952
rect 11112 31949 11118 31952
rect 11112 31943 11141 31949
rect 11129 31909 11141 31943
rect 11112 31903 11141 31909
rect 11609 31943 11667 31949
rect 11609 31909 11621 31943
rect 11655 31940 11667 31943
rect 11882 31940 11888 31952
rect 11655 31912 11888 31940
rect 11655 31909 11667 31912
rect 11609 31903 11667 31909
rect 11112 31900 11118 31903
rect 11882 31900 11888 31912
rect 11940 31940 11946 31952
rect 12250 31940 12256 31952
rect 11940 31912 12256 31940
rect 11940 31900 11946 31912
rect 12250 31900 12256 31912
rect 12308 31900 12314 31952
rect 12526 31900 12532 31952
rect 12584 31900 12590 31952
rect 14090 31900 14096 31952
rect 14148 31940 14154 31952
rect 14705 31943 14763 31949
rect 14705 31940 14717 31943
rect 14148 31912 14717 31940
rect 14148 31900 14154 31912
rect 4433 31875 4491 31881
rect 4433 31841 4445 31875
rect 4479 31872 4491 31875
rect 4614 31872 4620 31884
rect 4479 31844 4620 31872
rect 4479 31841 4491 31844
rect 4433 31835 4491 31841
rect 4614 31832 4620 31844
rect 4672 31832 4678 31884
rect 4890 31832 4896 31884
rect 4948 31832 4954 31884
rect 6914 31832 6920 31884
rect 6972 31832 6978 31884
rect 7926 31832 7932 31884
rect 7984 31872 7990 31884
rect 8021 31875 8079 31881
rect 8021 31872 8033 31875
rect 7984 31844 8033 31872
rect 7984 31832 7990 31844
rect 8021 31841 8033 31844
rect 8067 31841 8079 31875
rect 8021 31835 8079 31841
rect 10686 31832 10692 31884
rect 10744 31872 10750 31884
rect 10781 31875 10839 31881
rect 10781 31872 10793 31875
rect 10744 31844 10793 31872
rect 10744 31832 10750 31844
rect 10781 31841 10793 31844
rect 10827 31841 10839 31875
rect 10781 31835 10839 31841
rect 10870 31832 10876 31884
rect 10928 31832 10934 31884
rect 10962 31832 10968 31884
rect 11020 31832 11026 31884
rect 11333 31875 11391 31881
rect 11333 31841 11345 31875
rect 11379 31841 11391 31875
rect 11333 31835 11391 31841
rect 11425 31875 11483 31881
rect 11425 31841 11437 31875
rect 11471 31872 11483 31875
rect 11698 31872 11704 31884
rect 11471 31844 11704 31872
rect 11471 31841 11483 31844
rect 11425 31835 11483 31841
rect 3234 31764 3240 31816
rect 3292 31764 3298 31816
rect 6178 31764 6184 31816
rect 6236 31804 6242 31816
rect 6641 31807 6699 31813
rect 6641 31804 6653 31807
rect 6236 31776 6653 31804
rect 6236 31764 6242 31776
rect 6641 31773 6653 31776
rect 6687 31773 6699 31807
rect 6641 31767 6699 31773
rect 11241 31807 11299 31813
rect 11241 31773 11253 31807
rect 11287 31804 11299 31807
rect 11348 31804 11376 31835
rect 11698 31832 11704 31844
rect 11756 31872 11762 31884
rect 12158 31872 12164 31884
rect 11756 31844 12164 31872
rect 11756 31832 11762 31844
rect 12158 31832 12164 31844
rect 12216 31872 12222 31884
rect 12544 31872 12572 31900
rect 14292 31884 14320 31912
rect 14705 31909 14717 31912
rect 14751 31909 14763 31943
rect 14705 31903 14763 31909
rect 14826 31900 14832 31952
rect 14884 31940 14890 31952
rect 14921 31943 14979 31949
rect 14921 31940 14933 31943
rect 14884 31912 14933 31940
rect 14884 31900 14890 31912
rect 14921 31909 14933 31912
rect 14967 31940 14979 31943
rect 15197 31943 15255 31949
rect 15197 31940 15209 31943
rect 14967 31912 15209 31940
rect 14967 31909 14979 31912
rect 14921 31903 14979 31909
rect 15197 31909 15209 31912
rect 15243 31909 15255 31943
rect 15197 31903 15255 31909
rect 15378 31900 15384 31952
rect 15436 31900 15442 31952
rect 15562 31900 15568 31952
rect 15620 31900 15626 31952
rect 18782 31900 18788 31952
rect 18840 31900 18846 31952
rect 12216 31844 12572 31872
rect 12216 31832 12222 31844
rect 14274 31832 14280 31884
rect 14332 31832 14338 31884
rect 15289 31875 15347 31881
rect 15289 31841 15301 31875
rect 15335 31872 15347 31875
rect 15580 31872 15608 31900
rect 15335 31844 15608 31872
rect 18693 31875 18751 31881
rect 15335 31841 15347 31844
rect 15289 31835 15347 31841
rect 18693 31841 18705 31875
rect 18739 31872 18751 31875
rect 19150 31872 19156 31884
rect 18739 31844 19156 31872
rect 18739 31841 18751 31844
rect 18693 31835 18751 31841
rect 19150 31832 19156 31844
rect 19208 31832 19214 31884
rect 11287 31776 11376 31804
rect 11287 31773 11299 31776
rect 11241 31767 11299 31773
rect 11348 31748 11376 31776
rect 15746 31764 15752 31816
rect 15804 31804 15810 31816
rect 16574 31804 16580 31816
rect 15804 31776 16580 31804
rect 15804 31764 15810 31776
rect 16574 31764 16580 31776
rect 16632 31804 16638 31816
rect 16945 31807 17003 31813
rect 16945 31804 16957 31807
rect 16632 31776 16957 31804
rect 16632 31764 16638 31776
rect 16945 31773 16957 31776
rect 16991 31773 17003 31807
rect 16945 31767 17003 31773
rect 17770 31764 17776 31816
rect 17828 31764 17834 31816
rect 18969 31807 19027 31813
rect 18969 31804 18981 31807
rect 18927 31776 18981 31804
rect 18969 31773 18981 31776
rect 19015 31804 19027 31807
rect 19444 31804 19472 31971
rect 19794 31968 19800 31980
rect 19852 31968 19858 32020
rect 25222 31968 25228 32020
rect 25280 32008 25286 32020
rect 26050 32008 26056 32020
rect 25280 31980 26056 32008
rect 25280 31968 25286 31980
rect 26050 31968 26056 31980
rect 26108 31968 26114 32020
rect 30374 31968 30380 32020
rect 30432 31968 30438 32020
rect 23753 31943 23811 31949
rect 23753 31909 23765 31943
rect 23799 31940 23811 31943
rect 24026 31940 24032 31952
rect 23799 31912 24032 31940
rect 23799 31909 23811 31912
rect 23753 31903 23811 31909
rect 24026 31900 24032 31912
rect 24084 31900 24090 31952
rect 28905 31943 28963 31949
rect 28905 31909 28917 31943
rect 28951 31940 28963 31943
rect 29178 31940 29184 31952
rect 28951 31912 29184 31940
rect 28951 31909 28963 31912
rect 28905 31903 28963 31909
rect 29178 31900 29184 31912
rect 29236 31900 29242 31952
rect 31294 31940 31300 31952
rect 30130 31912 31300 31940
rect 31294 31900 31300 31912
rect 31352 31900 31358 31952
rect 33413 31943 33471 31949
rect 33413 31909 33425 31943
rect 33459 31940 33471 31943
rect 33502 31940 33508 31952
rect 33459 31912 33508 31940
rect 33459 31909 33471 31912
rect 33413 31903 33471 31909
rect 33502 31900 33508 31912
rect 33560 31900 33566 31952
rect 24854 31832 24860 31884
rect 24912 31832 24918 31884
rect 27614 31832 27620 31884
rect 27672 31832 27678 31884
rect 27893 31875 27951 31881
rect 27893 31841 27905 31875
rect 27939 31872 27951 31875
rect 28534 31872 28540 31884
rect 27939 31844 28540 31872
rect 27939 31841 27951 31844
rect 27893 31835 27951 31841
rect 28534 31832 28540 31844
rect 28592 31832 28598 31884
rect 32214 31832 32220 31884
rect 32272 31832 32278 31884
rect 19015 31776 19472 31804
rect 23477 31807 23535 31813
rect 19015 31773 19027 31776
rect 18969 31767 19027 31773
rect 23477 31773 23489 31807
rect 23523 31773 23535 31807
rect 28629 31807 28687 31813
rect 28629 31804 28641 31807
rect 23477 31767 23535 31773
rect 27632 31776 28641 31804
rect 11330 31696 11336 31748
rect 11388 31696 11394 31748
rect 14366 31696 14372 31748
rect 14424 31736 14430 31748
rect 14553 31739 14611 31745
rect 14553 31736 14565 31739
rect 14424 31708 14565 31736
rect 14424 31696 14430 31708
rect 14553 31705 14565 31708
rect 14599 31705 14611 31739
rect 14553 31699 14611 31705
rect 10594 31628 10600 31680
rect 10652 31628 10658 31680
rect 10870 31628 10876 31680
rect 10928 31668 10934 31680
rect 11517 31671 11575 31677
rect 11517 31668 11529 31671
rect 10928 31640 11529 31668
rect 10928 31628 10934 31640
rect 11517 31637 11529 31640
rect 11563 31637 11575 31671
rect 11517 31631 11575 31637
rect 11974 31628 11980 31680
rect 12032 31668 12038 31680
rect 14737 31671 14795 31677
rect 14737 31668 14749 31671
rect 12032 31640 14749 31668
rect 12032 31628 12038 31640
rect 14737 31637 14749 31640
rect 14783 31668 14795 31671
rect 14918 31668 14924 31680
rect 14783 31640 14924 31668
rect 14783 31637 14795 31640
rect 14737 31631 14795 31637
rect 14918 31628 14924 31640
rect 14976 31628 14982 31680
rect 17218 31628 17224 31680
rect 17276 31628 17282 31680
rect 17862 31628 17868 31680
rect 17920 31668 17926 31680
rect 18984 31668 19012 31767
rect 23492 31736 23520 31767
rect 27522 31736 27528 31748
rect 23308 31708 23520 31736
rect 26528 31708 27528 31736
rect 23308 31680 23336 31708
rect 26528 31680 26556 31708
rect 27522 31696 27528 31708
rect 27580 31736 27586 31748
rect 27632 31736 27660 31776
rect 28629 31773 28641 31776
rect 28675 31773 28687 31807
rect 28629 31767 28687 31773
rect 30558 31764 30564 31816
rect 30616 31804 30622 31816
rect 30653 31807 30711 31813
rect 30653 31804 30665 31807
rect 30616 31776 30665 31804
rect 30616 31764 30622 31776
rect 30653 31773 30665 31776
rect 30699 31773 30711 31807
rect 30653 31767 30711 31773
rect 31846 31764 31852 31816
rect 31904 31764 31910 31816
rect 32122 31764 32128 31816
rect 32180 31764 32186 31816
rect 27580 31708 27660 31736
rect 27580 31696 27586 31708
rect 17920 31640 19012 31668
rect 17920 31628 17926 31640
rect 23290 31628 23296 31680
rect 23348 31628 23354 31680
rect 26510 31628 26516 31680
rect 26568 31628 26574 31680
rect 26878 31628 26884 31680
rect 26936 31668 26942 31680
rect 26973 31671 27031 31677
rect 26973 31668 26985 31671
rect 26936 31640 26985 31668
rect 26936 31628 26942 31640
rect 26973 31637 26985 31640
rect 27019 31637 27031 31671
rect 26973 31631 27031 31637
rect 27798 31628 27804 31680
rect 27856 31628 27862 31680
rect 2760 31578 34316 31600
rect 2760 31526 6550 31578
rect 6602 31526 6614 31578
rect 6666 31526 6678 31578
rect 6730 31526 6742 31578
rect 6794 31526 6806 31578
rect 6858 31526 14439 31578
rect 14491 31526 14503 31578
rect 14555 31526 14567 31578
rect 14619 31526 14631 31578
rect 14683 31526 14695 31578
rect 14747 31526 22328 31578
rect 22380 31526 22392 31578
rect 22444 31526 22456 31578
rect 22508 31526 22520 31578
rect 22572 31526 22584 31578
rect 22636 31526 30217 31578
rect 30269 31526 30281 31578
rect 30333 31526 30345 31578
rect 30397 31526 30409 31578
rect 30461 31526 30473 31578
rect 30525 31526 34316 31578
rect 2760 31504 34316 31526
rect 4801 31467 4859 31473
rect 4801 31433 4813 31467
rect 4847 31464 4859 31467
rect 5442 31464 5448 31476
rect 4847 31436 5448 31464
rect 4847 31433 4859 31436
rect 4801 31427 4859 31433
rect 5442 31424 5448 31436
rect 5500 31424 5506 31476
rect 15289 31467 15347 31473
rect 15289 31433 15301 31467
rect 15335 31464 15347 31467
rect 15378 31464 15384 31476
rect 15335 31436 15384 31464
rect 15335 31433 15347 31436
rect 15289 31427 15347 31433
rect 15378 31424 15384 31436
rect 15436 31424 15442 31476
rect 15470 31424 15476 31476
rect 15528 31424 15534 31476
rect 18325 31467 18383 31473
rect 18325 31433 18337 31467
rect 18371 31464 18383 31467
rect 18414 31464 18420 31476
rect 18371 31436 18420 31464
rect 18371 31433 18383 31436
rect 18325 31427 18383 31433
rect 18414 31424 18420 31436
rect 18472 31424 18478 31476
rect 26786 31424 26792 31476
rect 26844 31464 26850 31476
rect 26844 31436 28212 31464
rect 26844 31424 26850 31436
rect 5074 31356 5080 31408
rect 5132 31396 5138 31408
rect 7006 31396 7012 31408
rect 5132 31368 7012 31396
rect 5132 31356 5138 31368
rect 3053 31331 3111 31337
rect 3053 31297 3065 31331
rect 3099 31328 3111 31331
rect 4890 31328 4896 31340
rect 3099 31300 4896 31328
rect 3099 31297 3111 31300
rect 3053 31291 3111 31297
rect 4890 31288 4896 31300
rect 4948 31288 4954 31340
rect 5920 31337 5948 31368
rect 7006 31356 7012 31368
rect 7064 31356 7070 31408
rect 5905 31331 5963 31337
rect 5905 31297 5917 31331
rect 5951 31297 5963 31331
rect 5905 31291 5963 31297
rect 10413 31331 10471 31337
rect 10413 31297 10425 31331
rect 10459 31328 10471 31331
rect 10594 31328 10600 31340
rect 10459 31300 10600 31328
rect 10459 31297 10471 31300
rect 10413 31291 10471 31297
rect 10594 31288 10600 31300
rect 10652 31288 10658 31340
rect 11974 31328 11980 31340
rect 10980 31300 11980 31328
rect 10980 31272 11008 31300
rect 11974 31288 11980 31300
rect 12032 31288 12038 31340
rect 16574 31288 16580 31340
rect 16632 31288 16638 31340
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31328 16911 31331
rect 17218 31328 17224 31340
rect 16899 31300 17224 31328
rect 16899 31297 16911 31300
rect 16853 31291 16911 31297
rect 17218 31288 17224 31300
rect 17276 31288 17282 31340
rect 18782 31288 18788 31340
rect 18840 31288 18846 31340
rect 22281 31331 22339 31337
rect 22281 31297 22293 31331
rect 22327 31328 22339 31331
rect 23290 31328 23296 31340
rect 22327 31300 23296 31328
rect 22327 31297 22339 31300
rect 22281 31291 22339 31297
rect 23290 31288 23296 31300
rect 23348 31288 23354 31340
rect 26510 31288 26516 31340
rect 26568 31288 26574 31340
rect 26789 31331 26847 31337
rect 26789 31297 26801 31331
rect 26835 31328 26847 31331
rect 26878 31328 26884 31340
rect 26835 31300 26884 31328
rect 26835 31297 26847 31300
rect 26789 31291 26847 31297
rect 26878 31288 26884 31300
rect 26936 31288 26942 31340
rect 5077 31263 5135 31269
rect 5077 31229 5089 31263
rect 5123 31229 5135 31263
rect 5077 31223 5135 31229
rect 3326 31152 3332 31204
rect 3384 31152 3390 31204
rect 4985 31195 5043 31201
rect 4985 31192 4997 31195
rect 4554 31164 4997 31192
rect 4985 31161 4997 31164
rect 5031 31161 5043 31195
rect 4985 31155 5043 31161
rect 5092 31192 5120 31223
rect 5534 31220 5540 31272
rect 5592 31220 5598 31272
rect 6914 31260 6920 31272
rect 5644 31232 6920 31260
rect 5644 31192 5672 31232
rect 6914 31220 6920 31232
rect 6972 31220 6978 31272
rect 7745 31263 7803 31269
rect 7745 31229 7757 31263
rect 7791 31260 7803 31263
rect 7834 31260 7840 31272
rect 7791 31232 7840 31260
rect 7791 31229 7803 31232
rect 7745 31223 7803 31229
rect 7834 31220 7840 31232
rect 7892 31260 7898 31272
rect 10134 31260 10140 31272
rect 7892 31232 10140 31260
rect 7892 31220 7898 31232
rect 10134 31220 10140 31232
rect 10192 31220 10198 31272
rect 10962 31220 10968 31272
rect 11020 31220 11026 31272
rect 11149 31263 11207 31269
rect 11149 31229 11161 31263
rect 11195 31229 11207 31263
rect 11149 31223 11207 31229
rect 5092 31164 5672 31192
rect 4890 31084 4896 31136
rect 4948 31124 4954 31136
rect 5092 31124 5120 31164
rect 6362 31152 6368 31204
rect 6420 31192 6426 31204
rect 6420 31164 10364 31192
rect 6420 31152 6426 31164
rect 10336 31136 10364 31164
rect 11164 31136 11192 31223
rect 11882 31152 11888 31204
rect 11940 31152 11946 31204
rect 4948 31096 5120 31124
rect 4948 31084 4954 31096
rect 7926 31084 7932 31136
rect 7984 31124 7990 31136
rect 9033 31127 9091 31133
rect 9033 31124 9045 31127
rect 7984 31096 9045 31124
rect 7984 31084 7990 31096
rect 9033 31093 9045 31096
rect 9079 31093 9091 31127
rect 9033 31087 9091 31093
rect 9766 31084 9772 31136
rect 9824 31084 9830 31136
rect 10318 31084 10324 31136
rect 10376 31084 10382 31136
rect 11146 31084 11152 31136
rect 11204 31084 11210 31136
rect 11330 31084 11336 31136
rect 11388 31124 11394 31136
rect 11900 31124 11928 31152
rect 11388 31096 11928 31124
rect 11992 31124 12020 31288
rect 12158 31220 12164 31272
rect 12216 31220 12222 31272
rect 15381 31263 15439 31269
rect 15381 31229 15393 31263
rect 15427 31229 15439 31263
rect 15381 31223 15439 31229
rect 15396 31192 15424 31223
rect 16482 31220 16488 31272
rect 16540 31220 16546 31272
rect 18417 31263 18475 31269
rect 18417 31229 18429 31263
rect 18463 31229 18475 31263
rect 18417 31223 18475 31229
rect 16574 31192 16580 31204
rect 15396 31164 16580 31192
rect 12069 31127 12127 31133
rect 12069 31124 12081 31127
rect 11992 31096 12081 31124
rect 11388 31084 11394 31096
rect 12069 31093 12081 31096
rect 12115 31093 12127 31127
rect 12069 31087 12127 31093
rect 12250 31084 12256 31136
rect 12308 31084 12314 31136
rect 12434 31084 12440 31136
rect 12492 31084 12498 31136
rect 13354 31084 13360 31136
rect 13412 31124 13418 31136
rect 15396 31124 15424 31164
rect 16574 31152 16580 31164
rect 16632 31152 16638 31204
rect 18138 31192 18144 31204
rect 18078 31164 18144 31192
rect 18138 31152 18144 31164
rect 18196 31152 18202 31204
rect 13412 31096 15424 31124
rect 13412 31084 13418 31096
rect 16298 31084 16304 31136
rect 16356 31084 16362 31136
rect 16592 31124 16620 31152
rect 18432 31124 18460 31223
rect 23658 31220 23664 31272
rect 23716 31220 23722 31272
rect 28184 31260 28212 31436
rect 31294 31424 31300 31476
rect 31352 31424 31358 31476
rect 28261 31331 28319 31337
rect 28261 31297 28273 31331
rect 28307 31328 28319 31331
rect 30006 31328 30012 31340
rect 28307 31300 30012 31328
rect 28307 31297 28319 31300
rect 28261 31291 28319 31297
rect 30006 31288 30012 31300
rect 30064 31288 30070 31340
rect 33778 31288 33784 31340
rect 33836 31288 33842 31340
rect 28353 31263 28411 31269
rect 28353 31260 28365 31263
rect 28184 31232 28365 31260
rect 28353 31229 28365 31232
rect 28399 31229 28411 31263
rect 28353 31223 28411 31229
rect 30742 31220 30748 31272
rect 30800 31220 30806 31272
rect 31389 31263 31447 31269
rect 31389 31229 31401 31263
rect 31435 31260 31447 31263
rect 31435 31232 31616 31260
rect 31435 31229 31447 31232
rect 31389 31223 31447 31229
rect 31588 31204 31616 31232
rect 32490 31220 32496 31272
rect 32548 31220 32554 31272
rect 32766 31220 32772 31272
rect 32824 31220 32830 31272
rect 22554 31152 22560 31204
rect 22612 31152 22618 31204
rect 27798 31152 27804 31204
rect 27856 31152 27862 31204
rect 28718 31152 28724 31204
rect 28776 31192 28782 31204
rect 29181 31195 29239 31201
rect 29181 31192 29193 31195
rect 28776 31164 29193 31192
rect 28776 31152 28782 31164
rect 29181 31161 29193 31164
rect 29227 31192 29239 31195
rect 31570 31192 31576 31204
rect 29227 31164 31576 31192
rect 29227 31161 29239 31164
rect 29181 31155 29239 31161
rect 31570 31152 31576 31164
rect 31628 31152 31634 31204
rect 31757 31195 31815 31201
rect 31757 31161 31769 31195
rect 31803 31192 31815 31195
rect 32030 31192 32036 31204
rect 31803 31164 32036 31192
rect 31803 31161 31815 31164
rect 31757 31155 31815 31161
rect 32030 31152 32036 31164
rect 32088 31152 32094 31204
rect 16592 31096 18460 31124
rect 24029 31127 24087 31133
rect 24029 31093 24041 31127
rect 24075 31124 24087 31127
rect 24118 31124 24124 31136
rect 24075 31096 24124 31124
rect 24075 31093 24087 31096
rect 24029 31087 24087 31093
rect 24118 31084 24124 31096
rect 24176 31124 24182 31136
rect 24762 31124 24768 31136
rect 24176 31096 24768 31124
rect 24176 31084 24182 31096
rect 24762 31084 24768 31096
rect 24820 31084 24826 31136
rect 28534 31084 28540 31136
rect 28592 31124 28598 31136
rect 29457 31127 29515 31133
rect 29457 31124 29469 31127
rect 28592 31096 29469 31124
rect 28592 31084 28598 31096
rect 29457 31093 29469 31096
rect 29503 31093 29515 31127
rect 29457 31087 29515 31093
rect 30190 31084 30196 31136
rect 30248 31084 30254 31136
rect 31846 31084 31852 31136
rect 31904 31084 31910 31136
rect 2760 31034 34316 31056
rect 2760 30982 7210 31034
rect 7262 30982 7274 31034
rect 7326 30982 7338 31034
rect 7390 30982 7402 31034
rect 7454 30982 7466 31034
rect 7518 30982 15099 31034
rect 15151 30982 15163 31034
rect 15215 30982 15227 31034
rect 15279 30982 15291 31034
rect 15343 30982 15355 31034
rect 15407 30982 22988 31034
rect 23040 30982 23052 31034
rect 23104 30982 23116 31034
rect 23168 30982 23180 31034
rect 23232 30982 23244 31034
rect 23296 30982 30877 31034
rect 30929 30982 30941 31034
rect 30993 30982 31005 31034
rect 31057 30982 31069 31034
rect 31121 30982 31133 31034
rect 31185 30982 34316 31034
rect 2760 30960 34316 30982
rect 4890 30920 4896 30932
rect 4632 30892 4896 30920
rect 3973 30855 4031 30861
rect 3973 30821 3985 30855
rect 4019 30852 4031 30855
rect 4632 30852 4660 30892
rect 4890 30880 4896 30892
rect 4948 30880 4954 30932
rect 6362 30880 6368 30932
rect 6420 30880 6426 30932
rect 8389 30923 8447 30929
rect 8389 30889 8401 30923
rect 8435 30920 8447 30923
rect 8938 30920 8944 30932
rect 8435 30892 8944 30920
rect 8435 30889 8447 30892
rect 8389 30883 8447 30889
rect 8938 30880 8944 30892
rect 8996 30880 9002 30932
rect 9214 30920 9220 30932
rect 9048 30892 9220 30920
rect 4019 30824 4660 30852
rect 4019 30821 4031 30824
rect 3973 30815 4031 30821
rect 4706 30812 4712 30864
rect 4764 30852 4770 30864
rect 5350 30852 5356 30864
rect 4764 30824 5356 30852
rect 4764 30812 4770 30824
rect 5350 30812 5356 30824
rect 5408 30812 5414 30864
rect 8849 30855 8907 30861
rect 8849 30821 8861 30855
rect 8895 30852 8907 30855
rect 9048 30852 9076 30892
rect 9214 30880 9220 30892
rect 9272 30880 9278 30932
rect 9766 30920 9772 30932
rect 9508 30892 9772 30920
rect 9508 30861 9536 30892
rect 9766 30880 9772 30892
rect 9824 30880 9830 30932
rect 11698 30880 11704 30932
rect 11756 30880 11762 30932
rect 12434 30880 12440 30932
rect 12492 30880 12498 30932
rect 12618 30880 12624 30932
rect 12676 30920 12682 30932
rect 13354 30920 13360 30932
rect 12676 30892 13360 30920
rect 12676 30880 12682 30892
rect 13354 30880 13360 30892
rect 13412 30880 13418 30932
rect 16482 30880 16488 30932
rect 16540 30920 16546 30932
rect 16577 30923 16635 30929
rect 16577 30920 16589 30923
rect 16540 30892 16589 30920
rect 16540 30880 16546 30892
rect 16577 30889 16589 30892
rect 16623 30889 16635 30923
rect 16577 30883 16635 30889
rect 17313 30923 17371 30929
rect 17313 30889 17325 30923
rect 17359 30920 17371 30923
rect 17770 30920 17776 30932
rect 17359 30892 17776 30920
rect 17359 30889 17371 30892
rect 17313 30883 17371 30889
rect 17770 30880 17776 30892
rect 17828 30880 17834 30932
rect 18414 30880 18420 30932
rect 18472 30880 18478 30932
rect 18782 30880 18788 30932
rect 18840 30880 18846 30932
rect 22554 30880 22560 30932
rect 22612 30920 22618 30932
rect 23477 30923 23535 30929
rect 23477 30920 23489 30923
rect 22612 30892 23489 30920
rect 22612 30880 22618 30892
rect 23477 30889 23489 30892
rect 23523 30889 23535 30923
rect 23477 30883 23535 30889
rect 27522 30880 27528 30932
rect 27580 30880 27586 30932
rect 27617 30923 27675 30929
rect 27617 30889 27629 30923
rect 27663 30920 27675 30923
rect 28534 30920 28540 30932
rect 27663 30892 28540 30920
rect 27663 30889 27675 30892
rect 27617 30883 27675 30889
rect 28534 30880 28540 30892
rect 28592 30880 28598 30932
rect 30190 30920 30196 30932
rect 29288 30892 30196 30920
rect 8895 30824 9076 30852
rect 9493 30855 9551 30861
rect 8895 30821 8907 30824
rect 8849 30815 8907 30821
rect 9493 30821 9505 30855
rect 9539 30821 9551 30855
rect 11149 30855 11207 30861
rect 11149 30852 11161 30855
rect 10718 30824 11161 30852
rect 9493 30815 9551 30821
rect 11149 30821 11161 30824
rect 11195 30821 11207 30855
rect 11882 30852 11888 30864
rect 11149 30815 11207 30821
rect 11532 30824 11888 30852
rect 8294 30744 8300 30796
rect 8352 30744 8358 30796
rect 8757 30787 8815 30793
rect 8757 30753 8769 30787
rect 8803 30784 8815 30787
rect 8803 30756 9168 30784
rect 8803 30753 8815 30756
rect 8757 30747 8815 30753
rect 5258 30676 5264 30728
rect 5316 30676 5322 30728
rect 9033 30719 9091 30725
rect 9033 30685 9045 30719
rect 9079 30685 9091 30719
rect 9140 30716 9168 30756
rect 9214 30744 9220 30796
rect 9272 30744 9278 30796
rect 10778 30744 10784 30796
rect 10836 30784 10842 30796
rect 11532 30793 11560 30824
rect 11882 30812 11888 30824
rect 11940 30852 11946 30864
rect 12452 30852 12480 30880
rect 11940 30824 12388 30852
rect 12452 30824 12848 30852
rect 11940 30812 11946 30824
rect 11057 30787 11115 30793
rect 11057 30784 11069 30787
rect 10836 30756 11069 30784
rect 10836 30744 10842 30756
rect 11057 30753 11069 30756
rect 11103 30753 11115 30787
rect 11057 30747 11115 30753
rect 11517 30787 11575 30793
rect 11517 30753 11529 30787
rect 11563 30753 11575 30787
rect 11517 30747 11575 30753
rect 11793 30787 11851 30793
rect 11793 30753 11805 30787
rect 11839 30784 11851 30787
rect 12250 30784 12256 30796
rect 11839 30756 12256 30784
rect 11839 30753 11851 30756
rect 11793 30747 11851 30753
rect 12250 30744 12256 30756
rect 12308 30744 12314 30796
rect 12360 30784 12388 30824
rect 12434 30784 12440 30796
rect 12360 30756 12440 30784
rect 12434 30744 12440 30756
rect 12492 30744 12498 30796
rect 12618 30744 12624 30796
rect 12676 30744 12682 30796
rect 9140 30688 12434 30716
rect 9033 30679 9091 30685
rect 4154 30540 4160 30592
rect 4212 30580 4218 30592
rect 4985 30583 5043 30589
rect 4985 30580 4997 30583
rect 4212 30552 4997 30580
rect 4212 30540 4218 30552
rect 4985 30549 4997 30552
rect 5031 30549 5043 30583
rect 4985 30543 5043 30549
rect 5810 30540 5816 30592
rect 5868 30540 5874 30592
rect 8202 30540 8208 30592
rect 8260 30540 8266 30592
rect 9048 30580 9076 30679
rect 10686 30608 10692 30660
rect 10744 30648 10750 30660
rect 11333 30651 11391 30657
rect 11333 30648 11345 30651
rect 10744 30620 11345 30648
rect 10744 30608 10750 30620
rect 11333 30617 11345 30620
rect 11379 30617 11391 30651
rect 12406 30648 12434 30688
rect 12710 30676 12716 30728
rect 12768 30676 12774 30728
rect 12820 30725 12848 30824
rect 13372 30793 13400 30880
rect 16761 30855 16819 30861
rect 16761 30852 16773 30855
rect 16330 30824 16773 30852
rect 16761 30821 16773 30824
rect 16807 30821 16819 30855
rect 16761 30815 16819 30821
rect 13357 30787 13415 30793
rect 13357 30753 13369 30787
rect 13403 30753 13415 30787
rect 13357 30747 13415 30753
rect 14182 30744 14188 30796
rect 14240 30784 14246 30796
rect 14829 30787 14887 30793
rect 14829 30784 14841 30787
rect 14240 30756 14841 30784
rect 14240 30744 14246 30756
rect 14829 30753 14841 30756
rect 14875 30753 14887 30787
rect 14829 30747 14887 30753
rect 16574 30744 16580 30796
rect 16632 30784 16638 30796
rect 16853 30787 16911 30793
rect 16853 30784 16865 30787
rect 16632 30756 16865 30784
rect 16632 30744 16638 30756
rect 16853 30753 16865 30756
rect 16899 30753 16911 30787
rect 16853 30747 16911 30753
rect 17678 30744 17684 30796
rect 17736 30744 17742 30796
rect 17773 30787 17831 30793
rect 17773 30753 17785 30787
rect 17819 30784 17831 30787
rect 18432 30784 18460 30880
rect 17819 30756 18460 30784
rect 18509 30787 18567 30793
rect 17819 30753 17831 30756
rect 17773 30747 17831 30753
rect 18509 30753 18521 30787
rect 18555 30784 18567 30787
rect 18800 30784 18828 30880
rect 27540 30852 27568 30880
rect 29288 30861 29316 30892
rect 30190 30880 30196 30892
rect 30248 30880 30254 30932
rect 31570 30880 31576 30932
rect 31628 30920 31634 30932
rect 31628 30892 31800 30920
rect 31628 30880 31634 30892
rect 29273 30855 29331 30861
rect 27540 30824 29040 30852
rect 18555 30756 18828 30784
rect 18555 30753 18567 30756
rect 18509 30747 18567 30753
rect 12805 30719 12863 30725
rect 12805 30685 12817 30719
rect 12851 30685 12863 30719
rect 12805 30679 12863 30685
rect 15102 30676 15108 30728
rect 15160 30676 15166 30728
rect 17862 30716 17868 30728
rect 17144 30688 17868 30716
rect 14826 30648 14832 30660
rect 12406 30620 14832 30648
rect 11333 30611 11391 30617
rect 14826 30608 14832 30620
rect 14884 30608 14890 30660
rect 9582 30580 9588 30592
rect 9048 30552 9588 30580
rect 9582 30540 9588 30552
rect 9640 30540 9646 30592
rect 9674 30540 9680 30592
rect 9732 30580 9738 30592
rect 10778 30580 10784 30592
rect 9732 30552 10784 30580
rect 9732 30540 9738 30552
rect 10778 30540 10784 30552
rect 10836 30540 10842 30592
rect 10965 30583 11023 30589
rect 10965 30549 10977 30583
rect 11011 30580 11023 30583
rect 11146 30580 11152 30592
rect 11011 30552 11152 30580
rect 11011 30549 11023 30552
rect 10965 30543 11023 30549
rect 11146 30540 11152 30552
rect 11204 30580 11210 30592
rect 11974 30580 11980 30592
rect 11204 30552 11980 30580
rect 11204 30540 11210 30552
rect 11974 30540 11980 30552
rect 12032 30540 12038 30592
rect 12250 30540 12256 30592
rect 12308 30540 12314 30592
rect 13262 30540 13268 30592
rect 13320 30540 13326 30592
rect 14182 30540 14188 30592
rect 14240 30580 14246 30592
rect 17144 30589 17172 30688
rect 17862 30676 17868 30688
rect 17920 30676 17926 30728
rect 18138 30676 18144 30728
rect 18196 30716 18202 30728
rect 18417 30719 18475 30725
rect 18417 30716 18429 30719
rect 18196 30688 18429 30716
rect 18196 30676 18202 30688
rect 18417 30685 18429 30688
rect 18463 30685 18475 30719
rect 18417 30679 18475 30685
rect 17129 30583 17187 30589
rect 17129 30580 17141 30583
rect 14240 30552 17141 30580
rect 14240 30540 14246 30552
rect 17129 30549 17141 30552
rect 17175 30580 17187 30583
rect 17218 30580 17224 30592
rect 17175 30552 17224 30580
rect 17175 30549 17187 30552
rect 17129 30543 17187 30549
rect 17218 30540 17224 30552
rect 17276 30540 17282 30592
rect 17862 30540 17868 30592
rect 17920 30580 17926 30592
rect 18524 30580 18552 30747
rect 24762 30744 24768 30796
rect 24820 30744 24826 30796
rect 27525 30787 27583 30793
rect 27525 30753 27537 30787
rect 27571 30784 27583 30787
rect 27798 30784 27804 30796
rect 27571 30756 27804 30784
rect 27571 30753 27583 30756
rect 27525 30747 27583 30753
rect 27798 30744 27804 30756
rect 27856 30744 27862 30796
rect 29012 30793 29040 30824
rect 29273 30821 29285 30855
rect 29319 30821 29331 30855
rect 31665 30855 31723 30861
rect 31665 30852 31677 30855
rect 30498 30824 31677 30852
rect 29273 30815 29331 30821
rect 31665 30821 31677 30824
rect 31711 30821 31723 30855
rect 31665 30815 31723 30821
rect 28997 30787 29055 30793
rect 28997 30753 29009 30787
rect 29043 30753 29055 30787
rect 31386 30784 31392 30796
rect 28997 30747 29055 30753
rect 30760 30756 31392 30784
rect 19702 30676 19708 30728
rect 19760 30676 19766 30728
rect 24026 30676 24032 30728
rect 24084 30676 24090 30728
rect 25498 30676 25504 30728
rect 25556 30676 25562 30728
rect 27709 30719 27767 30725
rect 27709 30716 27721 30719
rect 26988 30688 27721 30716
rect 17920 30552 18552 30580
rect 17920 30540 17926 30552
rect 19150 30540 19156 30592
rect 19208 30540 19214 30592
rect 23474 30540 23480 30592
rect 23532 30580 23538 30592
rect 24213 30583 24271 30589
rect 24213 30580 24225 30583
rect 23532 30552 24225 30580
rect 23532 30540 23538 30552
rect 24213 30549 24225 30552
rect 24259 30549 24271 30583
rect 24213 30543 24271 30549
rect 24946 30540 24952 30592
rect 25004 30540 25010 30592
rect 26234 30540 26240 30592
rect 26292 30580 26298 30592
rect 26988 30589 27016 30688
rect 27709 30685 27721 30688
rect 27755 30716 27767 30719
rect 28258 30716 28264 30728
rect 27755 30688 28264 30716
rect 27755 30685 27767 30688
rect 27709 30679 27767 30685
rect 28258 30676 28264 30688
rect 28316 30676 28322 30728
rect 30760 30725 30788 30756
rect 31386 30744 31392 30756
rect 31444 30744 31450 30796
rect 31772 30793 31800 30892
rect 31846 30880 31852 30932
rect 31904 30920 31910 30932
rect 31904 30892 32168 30920
rect 31904 30880 31910 30892
rect 32140 30861 32168 30892
rect 33042 30880 33048 30932
rect 33100 30920 33106 30932
rect 33597 30923 33655 30929
rect 33597 30920 33609 30923
rect 33100 30892 33609 30920
rect 33100 30880 33106 30892
rect 33597 30889 33609 30892
rect 33643 30889 33655 30923
rect 33597 30883 33655 30889
rect 32125 30855 32183 30861
rect 32125 30821 32137 30855
rect 32171 30821 32183 30855
rect 33873 30855 33931 30861
rect 33873 30852 33885 30855
rect 33350 30824 33885 30852
rect 32125 30815 32183 30821
rect 33873 30821 33885 30824
rect 33919 30821 33931 30855
rect 33873 30815 33931 30821
rect 31757 30787 31815 30793
rect 31757 30753 31769 30787
rect 31803 30753 31815 30787
rect 31757 30747 31815 30753
rect 33781 30787 33839 30793
rect 33781 30753 33793 30787
rect 33827 30753 33839 30787
rect 33781 30747 33839 30753
rect 30745 30719 30803 30725
rect 30745 30685 30757 30719
rect 30791 30685 30803 30719
rect 30745 30679 30803 30685
rect 31849 30719 31907 30725
rect 31849 30685 31861 30719
rect 31895 30685 31907 30719
rect 31849 30679 31907 30685
rect 31864 30648 31892 30679
rect 31220 30620 31892 30648
rect 31220 30592 31248 30620
rect 26973 30583 27031 30589
rect 26973 30580 26985 30583
rect 26292 30552 26985 30580
rect 26292 30540 26298 30552
rect 26973 30549 26985 30552
rect 27019 30549 27031 30583
rect 26973 30543 27031 30549
rect 27157 30583 27215 30589
rect 27157 30549 27169 30583
rect 27203 30580 27215 30583
rect 27614 30580 27620 30592
rect 27203 30552 27620 30580
rect 27203 30549 27215 30552
rect 27157 30543 27215 30549
rect 27614 30540 27620 30552
rect 27672 30540 27678 30592
rect 28905 30583 28963 30589
rect 28905 30549 28917 30583
rect 28951 30580 28963 30583
rect 29086 30580 29092 30592
rect 28951 30552 29092 30580
rect 28951 30549 28963 30552
rect 28905 30543 28963 30549
rect 29086 30540 29092 30552
rect 29144 30540 29150 30592
rect 30834 30540 30840 30592
rect 30892 30540 30898 30592
rect 31202 30540 31208 30592
rect 31260 30540 31266 30592
rect 31386 30540 31392 30592
rect 31444 30580 31450 30592
rect 31570 30580 31576 30592
rect 31444 30552 31576 30580
rect 31444 30540 31450 30552
rect 31570 30540 31576 30552
rect 31628 30580 31634 30592
rect 33796 30580 33824 30747
rect 31628 30552 33824 30580
rect 31628 30540 31634 30552
rect 2760 30490 34316 30512
rect 2760 30438 6550 30490
rect 6602 30438 6614 30490
rect 6666 30438 6678 30490
rect 6730 30438 6742 30490
rect 6794 30438 6806 30490
rect 6858 30438 14439 30490
rect 14491 30438 14503 30490
rect 14555 30438 14567 30490
rect 14619 30438 14631 30490
rect 14683 30438 14695 30490
rect 14747 30438 22328 30490
rect 22380 30438 22392 30490
rect 22444 30438 22456 30490
rect 22508 30438 22520 30490
rect 22572 30438 22584 30490
rect 22636 30438 30217 30490
rect 30269 30438 30281 30490
rect 30333 30438 30345 30490
rect 30397 30438 30409 30490
rect 30461 30438 30473 30490
rect 30525 30438 34316 30490
rect 2760 30416 34316 30438
rect 3326 30336 3332 30388
rect 3384 30376 3390 30388
rect 3789 30379 3847 30385
rect 3789 30376 3801 30379
rect 3384 30348 3801 30376
rect 3384 30336 3390 30348
rect 3789 30345 3801 30348
rect 3835 30345 3847 30379
rect 3789 30339 3847 30345
rect 5258 30336 5264 30388
rect 5316 30376 5322 30388
rect 5445 30379 5503 30385
rect 5445 30376 5457 30379
rect 5316 30348 5457 30376
rect 5316 30336 5322 30348
rect 5445 30345 5457 30348
rect 5491 30345 5503 30379
rect 5445 30339 5503 30345
rect 10318 30336 10324 30388
rect 10376 30376 10382 30388
rect 14182 30376 14188 30388
rect 10376 30348 14188 30376
rect 10376 30336 10382 30348
rect 14182 30336 14188 30348
rect 14240 30336 14246 30388
rect 14921 30379 14979 30385
rect 14921 30345 14933 30379
rect 14967 30376 14979 30379
rect 15102 30376 15108 30388
rect 14967 30348 15108 30376
rect 14967 30345 14979 30348
rect 14921 30339 14979 30345
rect 15102 30336 15108 30348
rect 15160 30336 15166 30388
rect 23569 30379 23627 30385
rect 23569 30345 23581 30379
rect 23615 30376 23627 30379
rect 24026 30376 24032 30388
rect 23615 30348 24032 30376
rect 23615 30345 23627 30348
rect 23569 30339 23627 30345
rect 24026 30336 24032 30348
rect 24084 30336 24090 30388
rect 30742 30336 30748 30388
rect 30800 30336 30806 30388
rect 32766 30336 32772 30388
rect 32824 30376 32830 30388
rect 32953 30379 33011 30385
rect 32953 30376 32965 30379
rect 32824 30348 32965 30376
rect 32824 30336 32830 30348
rect 32953 30345 32965 30348
rect 32999 30345 33011 30379
rect 32953 30339 33011 30345
rect 3697 30311 3755 30317
rect 3697 30277 3709 30311
rect 3743 30308 3755 30311
rect 23474 30308 23480 30320
rect 3743 30280 6132 30308
rect 3743 30277 3755 30280
rect 3697 30271 3755 30277
rect 4448 30249 4476 30280
rect 4433 30243 4491 30249
rect 4433 30209 4445 30243
rect 4479 30209 4491 30243
rect 4433 30203 4491 30209
rect 5261 30243 5319 30249
rect 5261 30209 5273 30243
rect 5307 30240 5319 30243
rect 5442 30240 5448 30252
rect 5307 30212 5448 30240
rect 5307 30209 5319 30212
rect 5261 30203 5319 30209
rect 5442 30200 5448 30212
rect 5500 30200 5506 30252
rect 5994 30240 6000 30252
rect 5736 30212 6000 30240
rect 4154 30132 4160 30184
rect 4212 30172 4218 30184
rect 5736 30172 5764 30212
rect 5994 30200 6000 30212
rect 6052 30200 6058 30252
rect 6104 30249 6132 30280
rect 23124 30280 23480 30308
rect 6089 30243 6147 30249
rect 6089 30209 6101 30243
rect 6135 30240 6147 30243
rect 6362 30240 6368 30252
rect 6135 30212 6368 30240
rect 6135 30209 6147 30212
rect 6089 30203 6147 30209
rect 6362 30200 6368 30212
rect 6420 30200 6426 30252
rect 7006 30240 7012 30252
rect 6748 30212 7012 30240
rect 4212 30144 5764 30172
rect 5813 30175 5871 30181
rect 4212 30132 4218 30144
rect 5813 30141 5825 30175
rect 5859 30172 5871 30175
rect 6748 30172 6776 30212
rect 7006 30200 7012 30212
rect 7064 30200 7070 30252
rect 7926 30200 7932 30252
rect 7984 30240 7990 30252
rect 9214 30240 9220 30252
rect 7984 30212 9220 30240
rect 7984 30200 7990 30212
rect 9214 30200 9220 30212
rect 9272 30240 9278 30252
rect 11977 30243 12035 30249
rect 11977 30240 11989 30243
rect 9272 30212 11989 30240
rect 9272 30200 9278 30212
rect 11977 30209 11989 30212
rect 12023 30209 12035 30243
rect 11977 30203 12035 30209
rect 12250 30200 12256 30252
rect 12308 30200 12314 30252
rect 15654 30200 15660 30252
rect 15712 30240 15718 30252
rect 23124 30249 23152 30280
rect 23474 30268 23480 30280
rect 23532 30268 23538 30320
rect 23658 30268 23664 30320
rect 23716 30308 23722 30320
rect 23753 30311 23811 30317
rect 23753 30308 23765 30311
rect 23716 30280 23765 30308
rect 23716 30268 23722 30280
rect 23753 30277 23765 30280
rect 23799 30277 23811 30311
rect 23753 30271 23811 30277
rect 25774 30268 25780 30320
rect 25832 30308 25838 30320
rect 30193 30311 30251 30317
rect 25832 30280 29592 30308
rect 25832 30268 25838 30280
rect 23017 30243 23075 30249
rect 15712 30212 15976 30240
rect 15712 30200 15718 30212
rect 5859 30144 6776 30172
rect 5859 30141 5871 30144
rect 5813 30135 5871 30141
rect 6822 30132 6828 30184
rect 6880 30172 6886 30184
rect 6917 30175 6975 30181
rect 6917 30172 6929 30175
rect 6880 30144 6929 30172
rect 6880 30132 6886 30144
rect 6917 30141 6929 30144
rect 6963 30141 6975 30175
rect 6917 30135 6975 30141
rect 7190 30132 7196 30184
rect 7248 30172 7254 30184
rect 11149 30175 11207 30181
rect 11149 30172 11161 30175
rect 7248 30144 7972 30172
rect 7248 30132 7254 30144
rect 1302 30064 1308 30116
rect 1360 30104 1366 30116
rect 3145 30107 3203 30113
rect 3145 30104 3157 30107
rect 1360 30076 3157 30104
rect 1360 30064 1366 30076
rect 3145 30073 3157 30076
rect 3191 30073 3203 30107
rect 3145 30067 3203 30073
rect 5718 30064 5724 30116
rect 5776 30104 5782 30116
rect 5776 30076 7144 30104
rect 5776 30064 5782 30076
rect 3234 29996 3240 30048
rect 3292 29996 3298 30048
rect 7116 30045 7144 30076
rect 7944 30048 7972 30144
rect 9692 30144 11161 30172
rect 8202 30064 8208 30116
rect 8260 30064 8266 30116
rect 8846 30064 8852 30116
rect 8904 30064 8910 30116
rect 9692 30048 9720 30144
rect 11149 30141 11161 30144
rect 11195 30141 11207 30175
rect 11149 30135 11207 30141
rect 13262 30132 13268 30184
rect 13320 30172 13326 30184
rect 15948 30181 15976 30212
rect 23017 30209 23029 30243
rect 23063 30209 23075 30243
rect 23017 30203 23075 30209
rect 23109 30243 23167 30249
rect 23109 30209 23121 30243
rect 23155 30209 23167 30243
rect 23109 30203 23167 30209
rect 15565 30175 15623 30181
rect 13320 30144 13386 30172
rect 13320 30132 13326 30144
rect 15565 30141 15577 30175
rect 15611 30172 15623 30175
rect 15749 30175 15807 30181
rect 15749 30172 15761 30175
rect 15611 30144 15761 30172
rect 15611 30141 15623 30144
rect 15565 30135 15623 30141
rect 15749 30141 15761 30144
rect 15795 30141 15807 30175
rect 15749 30135 15807 30141
rect 15933 30175 15991 30181
rect 15933 30141 15945 30175
rect 15979 30141 15991 30175
rect 15933 30135 15991 30141
rect 16022 30132 16028 30184
rect 16080 30172 16086 30184
rect 16209 30175 16267 30181
rect 16209 30172 16221 30175
rect 16080 30144 16221 30172
rect 16080 30132 16086 30144
rect 16209 30141 16221 30144
rect 16255 30141 16267 30175
rect 16209 30135 16267 30141
rect 16298 30132 16304 30184
rect 16356 30132 16362 30184
rect 16850 30132 16856 30184
rect 16908 30132 16914 30184
rect 14090 30064 14096 30116
rect 14148 30104 14154 30116
rect 16117 30107 16175 30113
rect 16117 30104 16129 30107
rect 14148 30076 16129 30104
rect 14148 30064 14154 30076
rect 16117 30073 16129 30076
rect 16163 30104 16175 30107
rect 16316 30104 16344 30132
rect 16163 30076 16344 30104
rect 23032 30104 23060 30203
rect 23382 30200 23388 30252
rect 23440 30240 23446 30252
rect 24026 30240 24032 30252
rect 23440 30212 24032 30240
rect 23440 30200 23446 30212
rect 24026 30200 24032 30212
rect 24084 30200 24090 30252
rect 24305 30243 24363 30249
rect 24305 30209 24317 30243
rect 24351 30240 24363 30243
rect 24946 30240 24952 30252
rect 24351 30212 24952 30240
rect 24351 30209 24363 30212
rect 24305 30203 24363 30209
rect 24946 30200 24952 30212
rect 25004 30200 25010 30252
rect 25038 30200 25044 30252
rect 25096 30240 25102 30252
rect 25096 30212 26280 30240
rect 25096 30200 25102 30212
rect 26252 30181 26280 30212
rect 26786 30200 26792 30252
rect 26844 30240 26850 30252
rect 29564 30249 29592 30280
rect 30193 30277 30205 30311
rect 30239 30308 30251 30311
rect 30760 30308 30788 30336
rect 30239 30280 30788 30308
rect 30239 30277 30251 30280
rect 30193 30271 30251 30277
rect 29549 30243 29607 30249
rect 26844 30212 26924 30240
rect 26844 30200 26850 30212
rect 23845 30175 23903 30181
rect 23845 30141 23857 30175
rect 23891 30141 23903 30175
rect 23845 30135 23903 30141
rect 26237 30175 26295 30181
rect 26237 30141 26249 30175
rect 26283 30172 26295 30175
rect 26694 30172 26700 30184
rect 26283 30144 26700 30172
rect 26283 30141 26295 30144
rect 26237 30135 26295 30141
rect 23032 30076 23612 30104
rect 16163 30073 16175 30076
rect 16117 30067 16175 30073
rect 23584 30048 23612 30076
rect 4249 30039 4307 30045
rect 4249 30005 4261 30039
rect 4295 30036 4307 30039
rect 4617 30039 4675 30045
rect 4617 30036 4629 30039
rect 4295 30008 4629 30036
rect 4295 30005 4307 30008
rect 4249 29999 4307 30005
rect 4617 30005 4629 30008
rect 4663 30005 4675 30039
rect 4617 29999 4675 30005
rect 5905 30039 5963 30045
rect 5905 30005 5917 30039
rect 5951 30036 5963 30039
rect 6273 30039 6331 30045
rect 6273 30036 6285 30039
rect 5951 30008 6285 30036
rect 5951 30005 5963 30008
rect 5905 29999 5963 30005
rect 6273 30005 6285 30008
rect 6319 30005 6331 30039
rect 6273 29999 6331 30005
rect 7101 30039 7159 30045
rect 7101 30005 7113 30039
rect 7147 30005 7159 30039
rect 7101 29999 7159 30005
rect 7926 29996 7932 30048
rect 7984 29996 7990 30048
rect 9674 29996 9680 30048
rect 9732 29996 9738 30048
rect 9766 29996 9772 30048
rect 9824 30036 9830 30048
rect 10134 30036 10140 30048
rect 9824 30008 10140 30036
rect 9824 29996 9830 30008
rect 10134 29996 10140 30008
rect 10192 29996 10198 30048
rect 10597 30039 10655 30045
rect 10597 30005 10609 30039
rect 10643 30036 10655 30039
rect 10962 30036 10968 30048
rect 10643 30008 10968 30036
rect 10643 30005 10655 30008
rect 10597 29999 10655 30005
rect 10962 29996 10968 30008
rect 11020 29996 11026 30048
rect 12250 29996 12256 30048
rect 12308 30036 12314 30048
rect 12894 30036 12900 30048
rect 12308 30008 12900 30036
rect 12308 29996 12314 30008
rect 12894 29996 12900 30008
rect 12952 29996 12958 30048
rect 12986 29996 12992 30048
rect 13044 30036 13050 30048
rect 13725 30039 13783 30045
rect 13725 30036 13737 30039
rect 13044 30008 13737 30036
rect 13044 29996 13050 30008
rect 13725 30005 13737 30008
rect 13771 30005 13783 30039
rect 13725 29999 13783 30005
rect 16206 29996 16212 30048
rect 16264 30036 16270 30048
rect 16301 30039 16359 30045
rect 16301 30036 16313 30039
rect 16264 30008 16313 30036
rect 16264 29996 16270 30008
rect 16301 30005 16313 30008
rect 16347 30005 16359 30039
rect 16301 29999 16359 30005
rect 23201 30039 23259 30045
rect 23201 30005 23213 30039
rect 23247 30036 23259 30039
rect 23382 30036 23388 30048
rect 23247 30008 23388 30036
rect 23247 30005 23259 30008
rect 23201 29999 23259 30005
rect 23382 29996 23388 30008
rect 23440 29996 23446 30048
rect 23566 29996 23572 30048
rect 23624 29996 23630 30048
rect 23860 30036 23888 30135
rect 26694 30132 26700 30144
rect 26752 30132 26758 30184
rect 26896 30181 26924 30212
rect 29549 30209 29561 30243
rect 29595 30209 29607 30243
rect 29549 30203 29607 30209
rect 29733 30243 29791 30249
rect 29733 30209 29745 30243
rect 29779 30240 29791 30243
rect 30834 30240 30840 30252
rect 29779 30212 30840 30240
rect 29779 30209 29791 30212
rect 29733 30203 29791 30209
rect 26881 30175 26939 30181
rect 26881 30141 26893 30175
rect 26927 30141 26939 30175
rect 26881 30135 26939 30141
rect 28534 30132 28540 30184
rect 28592 30132 28598 30184
rect 29362 30132 29368 30184
rect 29420 30132 29426 30184
rect 29564 30172 29592 30203
rect 30834 30200 30840 30212
rect 30892 30200 30898 30252
rect 30374 30172 30380 30184
rect 29564 30144 30380 30172
rect 30374 30132 30380 30144
rect 30432 30132 30438 30184
rect 30466 30132 30472 30184
rect 30524 30132 30530 30184
rect 30650 30132 30656 30184
rect 30708 30172 30714 30184
rect 31202 30172 31208 30184
rect 30708 30144 31208 30172
rect 30708 30132 30714 30144
rect 31202 30132 31208 30144
rect 31260 30132 31266 30184
rect 33689 30175 33747 30181
rect 33689 30141 33701 30175
rect 33735 30141 33747 30175
rect 33689 30135 33747 30141
rect 33965 30175 34023 30181
rect 33965 30141 33977 30175
rect 34011 30172 34023 30175
rect 35158 30172 35164 30184
rect 34011 30144 35164 30172
rect 34011 30141 34023 30144
rect 33965 30135 34023 30141
rect 26145 30107 26203 30113
rect 26145 30104 26157 30107
rect 25530 30076 26157 30104
rect 26145 30073 26157 30076
rect 26191 30073 26203 30107
rect 31021 30107 31079 30113
rect 26145 30067 26203 30073
rect 26804 30076 29960 30104
rect 25038 30036 25044 30048
rect 23860 30008 25044 30036
rect 25038 29996 25044 30008
rect 25096 29996 25102 30048
rect 25222 29996 25228 30048
rect 25280 30036 25286 30048
rect 25777 30039 25835 30045
rect 25777 30036 25789 30039
rect 25280 30008 25789 30036
rect 25280 29996 25286 30008
rect 25777 30005 25789 30008
rect 25823 30036 25835 30039
rect 26804 30036 26832 30076
rect 25823 30008 26832 30036
rect 25823 30005 25835 30008
rect 25777 29999 25835 30005
rect 26878 29996 26884 30048
rect 26936 30036 26942 30048
rect 26973 30039 27031 30045
rect 26973 30036 26985 30039
rect 26936 30008 26985 30036
rect 26936 29996 26942 30008
rect 26973 30005 26985 30008
rect 27019 30005 27031 30039
rect 26973 29999 27031 30005
rect 27433 30039 27491 30045
rect 27433 30005 27445 30039
rect 27479 30036 27491 30039
rect 27614 30036 27620 30048
rect 27479 30008 27620 30036
rect 27479 30005 27491 30008
rect 27433 29999 27491 30005
rect 27614 29996 27620 30008
rect 27672 29996 27678 30048
rect 27706 29996 27712 30048
rect 27764 29996 27770 30048
rect 27893 30039 27951 30045
rect 27893 30005 27905 30039
rect 27939 30036 27951 30039
rect 27982 30036 27988 30048
rect 27939 30008 27988 30036
rect 27939 30005 27951 30008
rect 27893 29999 27951 30005
rect 27982 29996 27988 30008
rect 28040 29996 28046 30048
rect 28721 30039 28779 30045
rect 28721 30005 28733 30039
rect 28767 30036 28779 30039
rect 28902 30036 28908 30048
rect 28767 30008 28908 30036
rect 28767 30005 28779 30008
rect 28721 29999 28779 30005
rect 28902 29996 28908 30008
rect 28960 30036 28966 30048
rect 29825 30039 29883 30045
rect 29825 30036 29837 30039
rect 28960 30008 29837 30036
rect 28960 29996 28966 30008
rect 29825 30005 29837 30008
rect 29871 30005 29883 30039
rect 29932 30036 29960 30076
rect 31021 30073 31033 30107
rect 31067 30104 31079 30107
rect 31481 30107 31539 30113
rect 31481 30104 31493 30107
rect 31067 30076 31493 30104
rect 31067 30073 31079 30076
rect 31021 30067 31079 30073
rect 31481 30073 31493 30076
rect 31527 30073 31539 30107
rect 31481 30067 31539 30073
rect 32214 30064 32220 30116
rect 32272 30064 32278 30116
rect 33704 30104 33732 30135
rect 35158 30132 35164 30144
rect 35216 30132 35222 30184
rect 34054 30104 34060 30116
rect 33704 30076 34060 30104
rect 34054 30064 34060 30076
rect 34112 30064 34118 30116
rect 32122 30036 32128 30048
rect 29932 30008 32128 30036
rect 29825 29999 29883 30005
rect 32122 29996 32128 30008
rect 32180 29996 32186 30048
rect 2760 29946 34316 29968
rect 2760 29894 7210 29946
rect 7262 29894 7274 29946
rect 7326 29894 7338 29946
rect 7390 29894 7402 29946
rect 7454 29894 7466 29946
rect 7518 29894 15099 29946
rect 15151 29894 15163 29946
rect 15215 29894 15227 29946
rect 15279 29894 15291 29946
rect 15343 29894 15355 29946
rect 15407 29894 22988 29946
rect 23040 29894 23052 29946
rect 23104 29894 23116 29946
rect 23168 29894 23180 29946
rect 23232 29894 23244 29946
rect 23296 29894 30877 29946
rect 30929 29894 30941 29946
rect 30993 29894 31005 29946
rect 31057 29894 31069 29946
rect 31121 29894 31133 29946
rect 31185 29894 34316 29946
rect 2760 29872 34316 29894
rect 5718 29792 5724 29844
rect 5776 29792 5782 29844
rect 5810 29792 5816 29844
rect 5868 29832 5874 29844
rect 5868 29804 6040 29832
rect 5868 29792 5874 29804
rect 5736 29764 5764 29792
rect 6012 29773 6040 29804
rect 8846 29792 8852 29844
rect 8904 29792 8910 29844
rect 9582 29792 9588 29844
rect 9640 29792 9646 29844
rect 9769 29835 9827 29841
rect 9769 29801 9781 29835
rect 9815 29832 9827 29835
rect 10318 29832 10324 29844
rect 9815 29804 10324 29832
rect 9815 29801 9827 29804
rect 9769 29795 9827 29801
rect 10318 29792 10324 29804
rect 10376 29832 10382 29844
rect 11054 29832 11060 29844
rect 10376 29804 11060 29832
rect 10376 29792 10382 29804
rect 11054 29792 11060 29804
rect 11112 29792 11118 29844
rect 12161 29835 12219 29841
rect 12161 29801 12173 29835
rect 12207 29832 12219 29835
rect 12618 29832 12624 29844
rect 12207 29804 12624 29832
rect 12207 29801 12219 29804
rect 12161 29795 12219 29801
rect 12618 29792 12624 29804
rect 12676 29792 12682 29844
rect 13173 29835 13231 29841
rect 13173 29801 13185 29835
rect 13219 29832 13231 29835
rect 13538 29832 13544 29844
rect 13219 29804 13544 29832
rect 13219 29801 13231 29804
rect 13173 29795 13231 29801
rect 13538 29792 13544 29804
rect 13596 29792 13602 29844
rect 14090 29792 14096 29844
rect 14148 29792 14154 29844
rect 14274 29792 14280 29844
rect 14332 29832 14338 29844
rect 14461 29835 14519 29841
rect 14461 29832 14473 29835
rect 14332 29804 14473 29832
rect 14332 29792 14338 29804
rect 14461 29801 14473 29804
rect 14507 29801 14519 29835
rect 14461 29795 14519 29801
rect 15473 29835 15531 29841
rect 15473 29801 15485 29835
rect 15519 29832 15531 29835
rect 16022 29832 16028 29844
rect 15519 29804 16028 29832
rect 15519 29801 15531 29804
rect 15473 29795 15531 29801
rect 16022 29792 16028 29804
rect 16080 29792 16086 29844
rect 16485 29835 16543 29841
rect 16485 29801 16497 29835
rect 16531 29832 16543 29835
rect 16850 29832 16856 29844
rect 16531 29804 16856 29832
rect 16531 29801 16543 29804
rect 16485 29795 16543 29801
rect 16850 29792 16856 29804
rect 16908 29792 16914 29844
rect 24857 29835 24915 29841
rect 24857 29801 24869 29835
rect 24903 29832 24915 29835
rect 25222 29832 25228 29844
rect 24903 29804 25228 29832
rect 24903 29801 24915 29804
rect 24857 29795 24915 29801
rect 25222 29792 25228 29804
rect 25280 29792 25286 29844
rect 25317 29835 25375 29841
rect 25317 29801 25329 29835
rect 25363 29832 25375 29835
rect 25498 29832 25504 29844
rect 25363 29804 25504 29832
rect 25363 29801 25375 29804
rect 25317 29795 25375 29801
rect 25498 29792 25504 29804
rect 25556 29792 25562 29844
rect 27709 29835 27767 29841
rect 27709 29801 27721 29835
rect 27755 29832 27767 29835
rect 27798 29832 27804 29844
rect 27755 29804 27804 29832
rect 27755 29801 27767 29804
rect 27709 29795 27767 29801
rect 27798 29792 27804 29804
rect 27856 29792 27862 29844
rect 28534 29792 28540 29844
rect 28592 29832 28598 29844
rect 28629 29835 28687 29841
rect 28629 29832 28641 29835
rect 28592 29804 28641 29832
rect 28592 29792 28598 29804
rect 28629 29801 28641 29804
rect 28675 29801 28687 29835
rect 28629 29795 28687 29801
rect 28902 29792 28908 29844
rect 28960 29792 28966 29844
rect 30466 29792 30472 29844
rect 30524 29832 30530 29844
rect 31113 29835 31171 29841
rect 31113 29832 31125 29835
rect 30524 29804 31125 29832
rect 30524 29792 30530 29804
rect 31113 29801 31125 29804
rect 31159 29801 31171 29835
rect 31113 29795 31171 29801
rect 32490 29792 32496 29844
rect 32548 29832 32554 29844
rect 32677 29835 32735 29841
rect 32677 29832 32689 29835
rect 32548 29804 32689 29832
rect 32548 29792 32554 29804
rect 32677 29801 32689 29804
rect 32723 29801 32735 29835
rect 32677 29795 32735 29801
rect 33042 29792 33048 29844
rect 33100 29832 33106 29844
rect 33137 29835 33195 29841
rect 33137 29832 33149 29835
rect 33100 29804 33149 29832
rect 33100 29792 33106 29804
rect 33137 29801 33149 29804
rect 33183 29801 33195 29835
rect 33137 29795 33195 29801
rect 5566 29736 5764 29764
rect 5997 29767 6055 29773
rect 5997 29733 6009 29767
rect 6043 29733 6055 29767
rect 5997 29727 6055 29733
rect 4433 29699 4491 29705
rect 4433 29665 4445 29699
rect 4479 29696 4491 29699
rect 4706 29696 4712 29708
rect 4479 29668 4712 29696
rect 4479 29665 4491 29668
rect 4433 29659 4491 29665
rect 4706 29656 4712 29668
rect 4764 29656 4770 29708
rect 6273 29699 6331 29705
rect 6273 29665 6285 29699
rect 6319 29696 6331 29699
rect 6319 29668 7604 29696
rect 6319 29665 6331 29668
rect 6273 29659 6331 29665
rect 7576 29640 7604 29668
rect 7926 29656 7932 29708
rect 7984 29696 7990 29708
rect 8757 29699 8815 29705
rect 8757 29696 8769 29699
rect 7984 29668 8769 29696
rect 7984 29656 7990 29668
rect 8757 29665 8769 29668
rect 8803 29696 8815 29699
rect 9600 29696 9628 29792
rect 9674 29724 9680 29776
rect 9732 29764 9738 29776
rect 11885 29767 11943 29773
rect 9732 29736 10732 29764
rect 9732 29724 9738 29736
rect 8803 29668 9628 29696
rect 8803 29665 8815 29668
rect 8757 29659 8815 29665
rect 10410 29656 10416 29708
rect 10468 29656 10474 29708
rect 10502 29656 10508 29708
rect 10560 29696 10566 29708
rect 10704 29705 10732 29736
rect 11885 29733 11897 29767
rect 11931 29764 11943 29767
rect 12710 29764 12716 29776
rect 11931 29736 12716 29764
rect 11931 29733 11943 29736
rect 11885 29727 11943 29733
rect 10597 29699 10655 29705
rect 10597 29696 10609 29699
rect 10560 29668 10609 29696
rect 10560 29656 10566 29668
rect 10597 29665 10609 29668
rect 10643 29665 10655 29699
rect 10597 29659 10655 29665
rect 10689 29699 10747 29705
rect 10689 29665 10701 29699
rect 10735 29696 10747 29699
rect 10778 29696 10784 29708
rect 10735 29668 10784 29696
rect 10735 29665 10747 29668
rect 10689 29659 10747 29665
rect 10778 29656 10784 29668
rect 10836 29656 10842 29708
rect 12084 29705 12112 29736
rect 12710 29724 12716 29736
rect 12768 29724 12774 29776
rect 12894 29724 12900 29776
rect 12952 29764 12958 29776
rect 14185 29767 14243 29773
rect 12952 29736 13584 29764
rect 12952 29724 12958 29736
rect 11977 29699 12035 29705
rect 11977 29665 11989 29699
rect 12023 29665 12035 29699
rect 11977 29659 12035 29665
rect 12069 29699 12127 29705
rect 12069 29665 12081 29699
rect 12115 29665 12127 29699
rect 12069 29659 12127 29665
rect 4065 29631 4123 29637
rect 4065 29597 4077 29631
rect 4111 29597 4123 29631
rect 4065 29591 4123 29597
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29628 4583 29631
rect 5626 29628 5632 29640
rect 4571 29600 5632 29628
rect 4571 29597 4583 29600
rect 4525 29591 4583 29597
rect 4080 29560 4108 29591
rect 5626 29588 5632 29600
rect 5684 29628 5690 29640
rect 6822 29628 6828 29640
rect 5684 29600 6828 29628
rect 5684 29588 5690 29600
rect 6822 29588 6828 29600
rect 6880 29588 6886 29640
rect 6914 29588 6920 29640
rect 6972 29588 6978 29640
rect 7558 29588 7564 29640
rect 7616 29588 7622 29640
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 9858 29588 9864 29640
rect 9916 29588 9922 29640
rect 10045 29631 10103 29637
rect 10045 29597 10057 29631
rect 10091 29628 10103 29631
rect 10962 29628 10968 29640
rect 10091 29600 10968 29628
rect 10091 29597 10103 29600
rect 10045 29591 10103 29597
rect 10962 29588 10968 29600
rect 11020 29588 11026 29640
rect 11992 29628 12020 29659
rect 12250 29656 12256 29708
rect 12308 29656 12314 29708
rect 12345 29699 12403 29705
rect 12345 29665 12357 29699
rect 12391 29696 12403 29699
rect 13357 29699 13415 29705
rect 13357 29696 13369 29699
rect 12391 29668 13369 29696
rect 12391 29665 12403 29668
rect 12345 29659 12403 29665
rect 13357 29665 13369 29668
rect 13403 29665 13415 29699
rect 13357 29659 13415 29665
rect 12360 29628 12388 29659
rect 11992 29600 12388 29628
rect 4982 29560 4988 29572
rect 4080 29532 4988 29560
rect 4982 29520 4988 29532
rect 5040 29520 5046 29572
rect 8312 29560 8340 29588
rect 12084 29572 12112 29600
rect 12986 29588 12992 29640
rect 13044 29588 13050 29640
rect 13449 29631 13507 29637
rect 13449 29597 13461 29631
rect 13495 29597 13507 29631
rect 13556 29628 13584 29736
rect 14185 29733 14197 29767
rect 14231 29764 14243 29767
rect 14826 29764 14832 29776
rect 14231 29736 14832 29764
rect 14231 29733 14243 29736
rect 14185 29727 14243 29733
rect 14826 29724 14832 29736
rect 14884 29724 14890 29776
rect 18325 29767 18383 29773
rect 18325 29764 18337 29767
rect 15212 29736 18337 29764
rect 13817 29699 13875 29705
rect 13817 29665 13829 29699
rect 13863 29696 13875 29699
rect 13906 29696 13912 29708
rect 13863 29668 13912 29696
rect 13863 29665 13875 29668
rect 13817 29659 13875 29665
rect 13906 29656 13912 29668
rect 13964 29656 13970 29708
rect 14277 29699 14335 29705
rect 14277 29665 14289 29699
rect 14323 29696 14335 29699
rect 15010 29696 15016 29708
rect 14323 29668 15016 29696
rect 14323 29665 14335 29668
rect 14277 29659 14335 29665
rect 15010 29656 15016 29668
rect 15068 29656 15074 29708
rect 15212 29705 15240 29736
rect 18325 29733 18337 29736
rect 18371 29733 18383 29767
rect 26234 29764 26240 29776
rect 18325 29727 18383 29733
rect 24780 29736 26240 29764
rect 15197 29699 15255 29705
rect 15197 29665 15209 29699
rect 15243 29665 15255 29699
rect 15197 29659 15255 29665
rect 15381 29699 15439 29705
rect 15381 29665 15393 29699
rect 15427 29665 15439 29699
rect 15381 29659 15439 29665
rect 15396 29628 15424 29659
rect 15470 29656 15476 29708
rect 15528 29696 15534 29708
rect 15565 29699 15623 29705
rect 15565 29696 15577 29699
rect 15528 29668 15577 29696
rect 15528 29656 15534 29668
rect 15565 29665 15577 29668
rect 15611 29696 15623 29699
rect 16117 29699 16175 29705
rect 16117 29696 16129 29699
rect 15611 29668 16129 29696
rect 15611 29665 15623 29668
rect 15565 29659 15623 29665
rect 16117 29665 16129 29668
rect 16163 29665 16175 29699
rect 16117 29659 16175 29665
rect 17586 29656 17592 29708
rect 17644 29656 17650 29708
rect 24780 29640 24808 29736
rect 26234 29724 26240 29736
rect 26292 29724 26298 29776
rect 26878 29724 26884 29776
rect 26936 29724 26942 29776
rect 27448 29736 28856 29764
rect 24949 29699 25007 29705
rect 24949 29665 24961 29699
rect 24995 29696 25007 29699
rect 25130 29696 25136 29708
rect 24995 29668 25136 29696
rect 24995 29665 25007 29668
rect 24949 29659 25007 29665
rect 25130 29656 25136 29668
rect 25188 29656 25194 29708
rect 13556 29600 15424 29628
rect 15933 29631 15991 29637
rect 13449 29591 13507 29597
rect 15933 29597 15945 29631
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 18969 29631 19027 29637
rect 18969 29597 18981 29631
rect 19015 29628 19027 29631
rect 20254 29628 20260 29640
rect 19015 29600 20260 29628
rect 19015 29597 19027 29600
rect 18969 29591 19027 29597
rect 9401 29563 9459 29569
rect 9401 29560 9413 29563
rect 8312 29532 9413 29560
rect 9401 29529 9413 29532
rect 9447 29529 9459 29563
rect 9401 29523 9459 29529
rect 12066 29520 12072 29572
rect 12124 29520 12130 29572
rect 12434 29520 12440 29572
rect 12492 29560 12498 29572
rect 13464 29560 13492 29591
rect 13814 29560 13820 29572
rect 12492 29532 13400 29560
rect 13464 29532 13820 29560
rect 12492 29520 12498 29532
rect 5442 29452 5448 29504
rect 5500 29492 5506 29504
rect 6365 29495 6423 29501
rect 6365 29492 6377 29495
rect 5500 29464 6377 29492
rect 5500 29452 5506 29464
rect 6365 29461 6377 29464
rect 6411 29461 6423 29495
rect 6365 29455 6423 29461
rect 10226 29452 10232 29504
rect 10284 29452 10290 29504
rect 13372 29501 13400 29532
rect 13814 29520 13820 29532
rect 13872 29520 13878 29572
rect 13909 29563 13967 29569
rect 13909 29529 13921 29563
rect 13955 29560 13967 29563
rect 13998 29560 14004 29572
rect 13955 29532 14004 29560
rect 13955 29529 13967 29532
rect 13909 29523 13967 29529
rect 13998 29520 14004 29532
rect 14056 29560 14062 29572
rect 15948 29560 15976 29591
rect 20254 29588 20260 29600
rect 20312 29588 20318 29640
rect 24762 29588 24768 29640
rect 24820 29588 24826 29640
rect 25869 29631 25927 29637
rect 25869 29597 25881 29631
rect 25915 29597 25927 29631
rect 25869 29591 25927 29597
rect 17405 29563 17463 29569
rect 17405 29560 17417 29563
rect 14056 29532 17417 29560
rect 14056 29520 14062 29532
rect 17405 29529 17417 29532
rect 17451 29529 17463 29563
rect 17405 29523 17463 29529
rect 23566 29520 23572 29572
rect 23624 29560 23630 29572
rect 24121 29563 24179 29569
rect 24121 29560 24133 29563
rect 23624 29532 24133 29560
rect 23624 29520 23630 29532
rect 24121 29529 24133 29532
rect 24167 29560 24179 29563
rect 25774 29560 25780 29572
rect 24167 29532 25780 29560
rect 24167 29529 24179 29532
rect 24121 29523 24179 29529
rect 25774 29520 25780 29532
rect 25832 29520 25838 29572
rect 13357 29495 13415 29501
rect 13357 29461 13369 29495
rect 13403 29461 13415 29495
rect 13357 29455 13415 29461
rect 14734 29452 14740 29504
rect 14792 29492 14798 29504
rect 15013 29495 15071 29501
rect 15013 29492 15025 29495
rect 14792 29464 15025 29492
rect 14792 29452 14798 29464
rect 15013 29461 15025 29464
rect 15059 29492 15071 29495
rect 21174 29492 21180 29504
rect 15059 29464 21180 29492
rect 15059 29461 15071 29464
rect 15013 29455 15071 29461
rect 21174 29452 21180 29464
rect 21232 29452 21238 29504
rect 23474 29452 23480 29504
rect 23532 29492 23538 29504
rect 23661 29495 23719 29501
rect 23661 29492 23673 29495
rect 23532 29464 23673 29492
rect 23532 29452 23538 29464
rect 23661 29461 23673 29464
rect 23707 29461 23719 29495
rect 23661 29455 23719 29461
rect 24489 29495 24547 29501
rect 24489 29461 24501 29495
rect 24535 29492 24547 29495
rect 24762 29492 24768 29504
rect 24535 29464 24768 29492
rect 24535 29461 24547 29464
rect 24489 29455 24547 29461
rect 24762 29452 24768 29464
rect 24820 29492 24826 29504
rect 24946 29492 24952 29504
rect 24820 29464 24952 29492
rect 24820 29452 24826 29464
rect 24946 29452 24952 29464
rect 25004 29452 25010 29504
rect 25884 29492 25912 29591
rect 26142 29588 26148 29640
rect 26200 29588 26206 29640
rect 26234 29588 26240 29640
rect 26292 29628 26298 29640
rect 27448 29628 27476 29736
rect 27890 29656 27896 29708
rect 27948 29696 27954 29708
rect 28828 29705 28856 29736
rect 28920 29705 28948 29792
rect 29086 29724 29092 29776
rect 29144 29764 29150 29776
rect 29273 29767 29331 29773
rect 29273 29764 29285 29767
rect 29144 29736 29285 29764
rect 29144 29724 29150 29736
rect 29273 29733 29285 29736
rect 29319 29733 29331 29767
rect 29273 29727 29331 29733
rect 30374 29724 30380 29776
rect 30432 29764 30438 29776
rect 31662 29764 31668 29776
rect 30432 29736 31668 29764
rect 30432 29724 30438 29736
rect 31662 29724 31668 29736
rect 31720 29764 31726 29776
rect 31720 29736 32168 29764
rect 31720 29724 31726 29736
rect 28813 29699 28871 29705
rect 27948 29668 28764 29696
rect 27948 29656 27954 29668
rect 26292 29600 27476 29628
rect 27617 29631 27675 29637
rect 26292 29588 26298 29600
rect 27617 29597 27629 29631
rect 27663 29628 27675 29631
rect 28261 29631 28319 29637
rect 28261 29628 28273 29631
rect 27663 29600 28273 29628
rect 27663 29597 27675 29600
rect 27617 29591 27675 29597
rect 28261 29597 28273 29600
rect 28307 29597 28319 29631
rect 28736 29628 28764 29668
rect 28813 29665 28825 29699
rect 28859 29665 28871 29699
rect 28813 29659 28871 29665
rect 28905 29699 28963 29705
rect 28905 29665 28917 29699
rect 28951 29665 28963 29699
rect 28905 29659 28963 29665
rect 28997 29699 29055 29705
rect 28997 29665 29009 29699
rect 29043 29665 29055 29699
rect 28997 29659 29055 29665
rect 29181 29699 29239 29705
rect 29181 29665 29193 29699
rect 29227 29665 29239 29699
rect 29181 29659 29239 29665
rect 29012 29628 29040 29659
rect 28736 29600 29040 29628
rect 28261 29591 28319 29597
rect 27706 29520 27712 29572
rect 27764 29560 27770 29572
rect 29196 29560 29224 29659
rect 30098 29656 30104 29708
rect 30156 29696 30162 29708
rect 31481 29699 31539 29705
rect 31481 29696 31493 29699
rect 30156 29668 31493 29696
rect 30156 29656 30162 29668
rect 31481 29665 31493 29668
rect 31527 29665 31539 29699
rect 31481 29659 31539 29665
rect 31573 29699 31631 29705
rect 31573 29665 31585 29699
rect 31619 29696 31631 29699
rect 31941 29699 31999 29705
rect 31941 29696 31953 29699
rect 31619 29668 31953 29696
rect 31619 29665 31631 29668
rect 31573 29659 31631 29665
rect 31941 29665 31953 29668
rect 31987 29665 31999 29699
rect 31941 29659 31999 29665
rect 31665 29631 31723 29637
rect 31665 29597 31677 29631
rect 31711 29628 31723 29631
rect 32030 29628 32036 29640
rect 31711 29600 32036 29628
rect 31711 29597 31723 29600
rect 31665 29591 31723 29597
rect 32030 29588 32036 29600
rect 32088 29588 32094 29640
rect 32140 29628 32168 29736
rect 32585 29699 32643 29705
rect 32585 29665 32597 29699
rect 32631 29696 32643 29699
rect 32766 29696 32772 29708
rect 32631 29668 32772 29696
rect 32631 29665 32643 29668
rect 32585 29659 32643 29665
rect 32766 29656 32772 29668
rect 32824 29656 32830 29708
rect 33042 29656 33048 29708
rect 33100 29656 33106 29708
rect 33229 29631 33287 29637
rect 33229 29628 33241 29631
rect 32140 29600 33241 29628
rect 33229 29597 33241 29600
rect 33275 29597 33287 29631
rect 33229 29591 33287 29597
rect 27764 29532 29224 29560
rect 27764 29520 27770 29532
rect 27522 29492 27528 29504
rect 25884 29464 27528 29492
rect 27522 29452 27528 29464
rect 27580 29452 27586 29504
rect 30561 29495 30619 29501
rect 30561 29461 30573 29495
rect 30607 29492 30619 29495
rect 30650 29492 30656 29504
rect 30607 29464 30656 29492
rect 30607 29461 30619 29464
rect 30561 29455 30619 29461
rect 30650 29452 30656 29464
rect 30708 29452 30714 29504
rect 2760 29402 34316 29424
rect 2760 29350 6550 29402
rect 6602 29350 6614 29402
rect 6666 29350 6678 29402
rect 6730 29350 6742 29402
rect 6794 29350 6806 29402
rect 6858 29350 14439 29402
rect 14491 29350 14503 29402
rect 14555 29350 14567 29402
rect 14619 29350 14631 29402
rect 14683 29350 14695 29402
rect 14747 29350 22328 29402
rect 22380 29350 22392 29402
rect 22444 29350 22456 29402
rect 22508 29350 22520 29402
rect 22572 29350 22584 29402
rect 22636 29350 30217 29402
rect 30269 29350 30281 29402
rect 30333 29350 30345 29402
rect 30397 29350 30409 29402
rect 30461 29350 30473 29402
rect 30525 29350 34316 29402
rect 2760 29328 34316 29350
rect 3053 29291 3111 29297
rect 3053 29257 3065 29291
rect 3099 29288 3111 29291
rect 4522 29288 4528 29300
rect 3099 29260 4528 29288
rect 3099 29257 3111 29260
rect 3053 29251 3111 29257
rect 4522 29248 4528 29260
rect 4580 29288 4586 29300
rect 4580 29260 5672 29288
rect 4580 29248 4586 29260
rect 5442 29180 5448 29232
rect 5500 29180 5506 29232
rect 4525 29155 4583 29161
rect 4525 29121 4537 29155
rect 4571 29152 4583 29155
rect 5460 29152 5488 29180
rect 4571 29124 5488 29152
rect 4571 29121 4583 29124
rect 4525 29115 4583 29121
rect 5534 29112 5540 29164
rect 5592 29112 5598 29164
rect 5644 29152 5672 29260
rect 5718 29248 5724 29300
rect 5776 29248 5782 29300
rect 6181 29291 6239 29297
rect 6181 29257 6193 29291
rect 6227 29288 6239 29291
rect 6914 29288 6920 29300
rect 6227 29260 6920 29288
rect 6227 29257 6239 29260
rect 6181 29251 6239 29257
rect 6914 29248 6920 29260
rect 6972 29248 6978 29300
rect 7024 29260 11928 29288
rect 5736 29220 5764 29248
rect 6457 29223 6515 29229
rect 6457 29220 6469 29223
rect 5736 29192 6469 29220
rect 6457 29189 6469 29192
rect 6503 29189 6515 29223
rect 6457 29183 6515 29189
rect 5721 29155 5779 29161
rect 5721 29152 5733 29155
rect 5644 29124 5733 29152
rect 5721 29121 5733 29124
rect 5767 29121 5779 29155
rect 5721 29115 5779 29121
rect 4801 29087 4859 29093
rect 4801 29053 4813 29087
rect 4847 29053 4859 29087
rect 4801 29047 4859 29053
rect 4816 29016 4844 29047
rect 4982 29044 4988 29096
rect 5040 29084 5046 29096
rect 5077 29087 5135 29093
rect 5077 29084 5089 29087
rect 5040 29056 5089 29084
rect 5040 29044 5046 29056
rect 5077 29053 5089 29056
rect 5123 29053 5135 29087
rect 5077 29047 5135 29053
rect 5166 29044 5172 29096
rect 5224 29084 5230 29096
rect 7024 29084 7052 29260
rect 11900 29220 11928 29260
rect 11974 29248 11980 29300
rect 12032 29248 12038 29300
rect 13078 29288 13084 29300
rect 12084 29260 13084 29288
rect 12084 29220 12112 29260
rect 13078 29248 13084 29260
rect 13136 29248 13142 29300
rect 14090 29248 14096 29300
rect 14148 29248 14154 29300
rect 15010 29288 15016 29300
rect 14936 29260 15016 29288
rect 11900 29192 12112 29220
rect 12253 29223 12311 29229
rect 12253 29189 12265 29223
rect 12299 29220 12311 29223
rect 12299 29192 12434 29220
rect 12299 29189 12311 29192
rect 12253 29183 12311 29189
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7558 29152 7564 29164
rect 7331 29124 7564 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7558 29112 7564 29124
rect 7616 29112 7622 29164
rect 9033 29155 9091 29161
rect 9033 29121 9045 29155
rect 9079 29121 9091 29155
rect 9033 29115 9091 29121
rect 5224 29056 7052 29084
rect 9048 29084 9076 29115
rect 10134 29112 10140 29164
rect 10192 29152 10198 29164
rect 12406 29152 12434 29192
rect 12894 29180 12900 29232
rect 12952 29220 12958 29232
rect 13633 29223 13691 29229
rect 13633 29220 13645 29223
rect 12952 29192 13645 29220
rect 12952 29180 12958 29192
rect 13633 29189 13645 29192
rect 13679 29189 13691 29223
rect 13633 29183 13691 29189
rect 12621 29155 12679 29161
rect 12621 29152 12633 29155
rect 10192 29124 11836 29152
rect 12406 29124 12633 29152
rect 10192 29112 10198 29124
rect 9493 29087 9551 29093
rect 9493 29084 9505 29087
rect 9048 29056 9505 29084
rect 5224 29044 5230 29056
rect 9493 29053 9505 29056
rect 9539 29084 9551 29087
rect 11609 29087 11667 29093
rect 10796 29084 11008 29086
rect 11609 29084 11621 29087
rect 9539 29058 11621 29084
rect 9539 29056 10824 29058
rect 10980 29056 11621 29058
rect 9539 29053 9551 29056
rect 9493 29047 9551 29053
rect 11609 29053 11621 29056
rect 11655 29053 11667 29087
rect 11609 29047 11667 29053
rect 11701 29087 11759 29093
rect 11701 29053 11713 29087
rect 11747 29053 11759 29087
rect 11701 29047 11759 29053
rect 5813 29019 5871 29025
rect 4094 28988 4476 29016
rect 4816 28988 5580 29016
rect 4448 28948 4476 28988
rect 5552 28960 5580 28988
rect 5813 28985 5825 29019
rect 5859 29016 5871 29019
rect 6362 29016 6368 29028
rect 5859 28988 6368 29016
rect 5859 28985 5871 28988
rect 5813 28979 5871 28985
rect 6362 28976 6368 28988
rect 6420 28976 6426 29028
rect 7561 29019 7619 29025
rect 7561 28985 7573 29019
rect 7607 29016 7619 29019
rect 7607 28988 7972 29016
rect 7607 28985 7619 28988
rect 7561 28979 7619 28985
rect 4985 28951 5043 28957
rect 4985 28948 4997 28951
rect 4448 28920 4997 28948
rect 4985 28917 4997 28920
rect 5031 28917 5043 28951
rect 4985 28911 5043 28917
rect 5534 28908 5540 28960
rect 5592 28908 5598 28960
rect 7944 28948 7972 28988
rect 8294 28976 8300 29028
rect 8352 28976 8358 29028
rect 10594 28976 10600 29028
rect 10652 28976 10658 29028
rect 11716 29016 11744 29047
rect 11440 28988 11744 29016
rect 11808 29016 11836 29124
rect 12621 29121 12633 29124
rect 12667 29121 12679 29155
rect 12621 29115 12679 29121
rect 13722 29112 13728 29164
rect 13780 29152 13786 29164
rect 13909 29155 13967 29161
rect 13909 29152 13921 29155
rect 13780 29124 13921 29152
rect 13780 29112 13786 29124
rect 13909 29121 13921 29124
rect 13955 29121 13967 29155
rect 13909 29115 13967 29121
rect 14090 29112 14096 29164
rect 14148 29152 14154 29164
rect 14461 29155 14519 29161
rect 14461 29152 14473 29155
rect 14148 29124 14473 29152
rect 14148 29112 14154 29124
rect 14461 29121 14473 29124
rect 14507 29152 14519 29155
rect 14642 29152 14648 29164
rect 14507 29124 14648 29152
rect 14507 29121 14519 29124
rect 14461 29115 14519 29121
rect 14642 29112 14648 29124
rect 14700 29112 14706 29164
rect 14826 29112 14832 29164
rect 14884 29112 14890 29164
rect 14936 29161 14964 29260
rect 15010 29248 15016 29260
rect 15068 29248 15074 29300
rect 15105 29291 15163 29297
rect 15105 29257 15117 29291
rect 15151 29288 15163 29291
rect 15654 29288 15660 29300
rect 15151 29260 15660 29288
rect 15151 29257 15163 29260
rect 15105 29251 15163 29257
rect 15654 29248 15660 29260
rect 15712 29248 15718 29300
rect 17586 29248 17592 29300
rect 17644 29248 17650 29300
rect 19429 29291 19487 29297
rect 19429 29257 19441 29291
rect 19475 29288 19487 29291
rect 19702 29288 19708 29300
rect 19475 29260 19708 29288
rect 19475 29257 19487 29260
rect 19429 29251 19487 29257
rect 19702 29248 19708 29260
rect 19760 29248 19766 29300
rect 22554 29248 22560 29300
rect 22612 29288 22618 29300
rect 23382 29288 23388 29300
rect 22612 29260 23388 29288
rect 22612 29248 22618 29260
rect 23382 29248 23388 29260
rect 23440 29288 23446 29300
rect 23753 29291 23811 29297
rect 23753 29288 23765 29291
rect 23440 29260 23765 29288
rect 23440 29248 23446 29260
rect 23753 29257 23765 29260
rect 23799 29257 23811 29291
rect 23753 29251 23811 29257
rect 25038 29248 25044 29300
rect 25096 29248 25102 29300
rect 26142 29248 26148 29300
rect 26200 29288 26206 29300
rect 26605 29291 26663 29297
rect 26605 29288 26617 29291
rect 26200 29260 26617 29288
rect 26200 29248 26206 29260
rect 26605 29257 26617 29260
rect 26651 29257 26663 29291
rect 26605 29251 26663 29257
rect 29362 29248 29368 29300
rect 29420 29288 29426 29300
rect 29457 29291 29515 29297
rect 29457 29288 29469 29291
rect 29420 29260 29469 29288
rect 29420 29248 29426 29260
rect 29457 29257 29469 29260
rect 29503 29257 29515 29291
rect 29457 29251 29515 29257
rect 32214 29248 32220 29300
rect 32272 29288 32278 29300
rect 32401 29291 32459 29297
rect 32401 29288 32413 29291
rect 32272 29260 32413 29288
rect 32272 29248 32278 29260
rect 32401 29257 32413 29260
rect 32447 29257 32459 29291
rect 32401 29251 32459 29257
rect 18984 29192 21404 29220
rect 14936 29155 15004 29161
rect 14936 29124 14958 29155
rect 14946 29121 14958 29124
rect 14992 29121 15004 29155
rect 14946 29115 15004 29121
rect 15838 29112 15844 29164
rect 15896 29112 15902 29164
rect 16117 29155 16175 29161
rect 16117 29121 16129 29155
rect 16163 29152 16175 29155
rect 16206 29152 16212 29164
rect 16163 29124 16212 29152
rect 16163 29121 16175 29124
rect 16117 29115 16175 29121
rect 16206 29112 16212 29124
rect 16264 29112 16270 29164
rect 16482 29112 16488 29164
rect 16540 29152 16546 29164
rect 18984 29152 19012 29192
rect 16540 29124 19012 29152
rect 21269 29155 21327 29161
rect 16540 29112 16546 29124
rect 21269 29121 21281 29155
rect 21315 29121 21327 29155
rect 21376 29152 21404 29192
rect 23017 29155 23075 29161
rect 21376 29124 22968 29152
rect 21269 29115 21327 29121
rect 12066 29044 12072 29096
rect 12124 29044 12130 29096
rect 13817 29087 13875 29093
rect 13817 29053 13829 29087
rect 13863 29084 13875 29087
rect 13998 29084 14004 29096
rect 13863 29056 14004 29084
rect 13863 29053 13875 29056
rect 13817 29047 13875 29053
rect 13998 29044 14004 29056
rect 14056 29044 14062 29096
rect 14737 29087 14795 29093
rect 14737 29053 14749 29087
rect 14783 29084 14795 29087
rect 14783 29056 14964 29084
rect 14783 29053 14795 29056
rect 14737 29047 14795 29053
rect 14936 29028 14964 29056
rect 17678 29044 17684 29096
rect 17736 29044 17742 29096
rect 19702 29044 19708 29096
rect 19760 29084 19766 29096
rect 19760 29056 20944 29084
rect 19760 29044 19766 29056
rect 11808 28988 13676 29016
rect 8478 28948 8484 28960
rect 7944 28920 8484 28948
rect 8478 28908 8484 28920
rect 8536 28908 8542 28960
rect 9677 28951 9735 28957
rect 9677 28917 9689 28951
rect 9723 28948 9735 28951
rect 10410 28948 10416 28960
rect 9723 28920 10416 28948
rect 9723 28917 9735 28920
rect 9677 28911 9735 28917
rect 10410 28908 10416 28920
rect 10468 28948 10474 28960
rect 10686 28948 10692 28960
rect 10468 28920 10692 28948
rect 10468 28908 10474 28920
rect 10686 28908 10692 28920
rect 10744 28948 10750 28960
rect 10781 28951 10839 28957
rect 10781 28948 10793 28951
rect 10744 28920 10793 28948
rect 10744 28908 10750 28920
rect 10781 28917 10793 28920
rect 10827 28917 10839 28951
rect 10781 28911 10839 28917
rect 10870 28908 10876 28960
rect 10928 28908 10934 28960
rect 10962 28908 10968 28960
rect 11020 28908 11026 28960
rect 11146 28908 11152 28960
rect 11204 28908 11210 28960
rect 11330 28908 11336 28960
rect 11388 28948 11394 28960
rect 11440 28948 11468 28988
rect 11388 28920 11468 28948
rect 11388 28908 11394 28920
rect 12986 28908 12992 28960
rect 13044 28948 13050 28960
rect 13265 28951 13323 28957
rect 13265 28948 13277 28951
rect 13044 28920 13277 28948
rect 13044 28908 13050 28920
rect 13265 28917 13277 28920
rect 13311 28917 13323 28951
rect 13648 28948 13676 28988
rect 13722 28976 13728 29028
rect 13780 29016 13786 29028
rect 14277 29019 14335 29025
rect 14277 29016 14289 29019
rect 13780 28988 14289 29016
rect 13780 28976 13786 28988
rect 14277 28985 14289 28988
rect 14323 28985 14335 29019
rect 14277 28979 14335 28985
rect 14366 28976 14372 29028
rect 14424 28976 14430 29028
rect 14918 28976 14924 29028
rect 14976 28976 14982 29028
rect 17126 28976 17132 29028
rect 17184 28976 17190 29028
rect 17954 28976 17960 29028
rect 18012 28976 18018 29028
rect 19613 29019 19671 29025
rect 19613 29016 19625 29019
rect 19182 28988 19625 29016
rect 19613 28985 19625 28988
rect 19659 28985 19671 29019
rect 19613 28979 19671 28985
rect 14384 28948 14412 28976
rect 20916 28960 20944 29056
rect 21284 29028 21312 29115
rect 22940 29084 22968 29124
rect 23017 29121 23029 29155
rect 23063 29152 23075 29155
rect 23109 29155 23167 29161
rect 23109 29152 23121 29155
rect 23063 29124 23121 29152
rect 23063 29121 23075 29124
rect 23017 29115 23075 29121
rect 23109 29121 23121 29124
rect 23155 29121 23167 29155
rect 24397 29155 24455 29161
rect 24397 29152 24409 29155
rect 23109 29115 23167 29121
rect 23492 29124 24409 29152
rect 23492 29096 23520 29124
rect 24397 29121 24409 29124
rect 24443 29121 24455 29155
rect 24397 29115 24455 29121
rect 23474 29084 23480 29096
rect 22940 29056 23480 29084
rect 23474 29044 23480 29056
rect 23532 29044 23538 29096
rect 23750 29044 23756 29096
rect 23808 29084 23814 29096
rect 23845 29087 23903 29093
rect 23845 29084 23857 29087
rect 23808 29056 23857 29084
rect 23808 29044 23814 29056
rect 23845 29053 23857 29056
rect 23891 29053 23903 29087
rect 23845 29047 23903 29053
rect 24765 29087 24823 29093
rect 24765 29053 24777 29087
rect 24811 29084 24823 29087
rect 25056 29084 25084 29248
rect 27522 29112 27528 29164
rect 27580 29152 27586 29164
rect 27709 29155 27767 29161
rect 27709 29152 27721 29155
rect 27580 29124 27721 29152
rect 27580 29112 27586 29124
rect 27709 29121 27721 29124
rect 27755 29121 27767 29155
rect 27709 29115 27767 29121
rect 27982 29112 27988 29164
rect 28040 29112 28046 29164
rect 28442 29112 28448 29164
rect 28500 29152 28506 29164
rect 29549 29155 29607 29161
rect 29549 29152 29561 29155
rect 28500 29124 29561 29152
rect 28500 29112 28506 29124
rect 29549 29121 29561 29124
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 24811 29056 25084 29084
rect 24811 29053 24823 29056
rect 24765 29047 24823 29053
rect 21266 28976 21272 29028
rect 21324 28976 21330 29028
rect 21542 28976 21548 29028
rect 21600 28976 21606 29028
rect 22830 29016 22836 29028
rect 22770 28988 22836 29016
rect 22830 28976 22836 28988
rect 22888 28976 22894 29028
rect 23382 28976 23388 29028
rect 23440 29016 23446 29028
rect 24780 29016 24808 29047
rect 27246 29044 27252 29096
rect 27304 29044 27310 29096
rect 30929 29087 30987 29093
rect 30929 29053 30941 29087
rect 30975 29084 30987 29087
rect 31202 29084 31208 29096
rect 30975 29056 31208 29084
rect 30975 29053 30987 29056
rect 30929 29047 30987 29053
rect 31202 29044 31208 29056
rect 31260 29044 31266 29096
rect 31846 29044 31852 29096
rect 31904 29044 31910 29096
rect 32033 29087 32091 29093
rect 32033 29084 32045 29087
rect 31956 29056 32045 29084
rect 23440 28988 24808 29016
rect 23440 28976 23446 28988
rect 26786 28976 26792 29028
rect 26844 29016 26850 29028
rect 26844 28988 27660 29016
rect 26844 28976 26850 28988
rect 13648 28920 14412 28948
rect 13265 28911 13323 28917
rect 20898 28908 20904 28960
rect 20956 28908 20962 28960
rect 24670 28908 24676 28960
rect 24728 28908 24734 28960
rect 26142 28908 26148 28960
rect 26200 28948 26206 28960
rect 26421 28951 26479 28957
rect 26421 28948 26433 28951
rect 26200 28920 26433 28948
rect 26200 28908 26206 28920
rect 26421 28917 26433 28920
rect 26467 28948 26479 28951
rect 27430 28948 27436 28960
rect 26467 28920 27436 28948
rect 26467 28917 26479 28920
rect 26421 28911 26479 28917
rect 27430 28908 27436 28920
rect 27488 28948 27494 28960
rect 27525 28951 27583 28957
rect 27525 28948 27537 28951
rect 27488 28920 27537 28948
rect 27488 28908 27494 28920
rect 27525 28917 27537 28920
rect 27571 28917 27583 28951
rect 27632 28948 27660 28988
rect 28994 28976 29000 29028
rect 29052 28976 29058 29028
rect 30098 28976 30104 29028
rect 30156 29016 30162 29028
rect 30285 29019 30343 29025
rect 30285 29016 30297 29019
rect 30156 28988 30297 29016
rect 30156 28976 30162 28988
rect 30285 28985 30297 28988
rect 30331 28985 30343 29019
rect 30285 28979 30343 28985
rect 28258 28948 28264 28960
rect 27632 28920 28264 28948
rect 27525 28911 27583 28917
rect 28258 28908 28264 28920
rect 28316 28908 28322 28960
rect 29362 28908 29368 28960
rect 29420 28948 29426 28960
rect 30193 28951 30251 28957
rect 30193 28948 30205 28951
rect 29420 28920 30205 28948
rect 29420 28908 29426 28920
rect 30193 28917 30205 28920
rect 30239 28917 30251 28951
rect 30193 28911 30251 28917
rect 31294 28908 31300 28960
rect 31352 28908 31358 28960
rect 31386 28908 31392 28960
rect 31444 28948 31450 28960
rect 31956 28948 31984 29056
rect 32033 29053 32045 29056
rect 32079 29084 32091 29087
rect 32493 29087 32551 29093
rect 32493 29084 32505 29087
rect 32079 29056 32505 29084
rect 32079 29053 32091 29056
rect 32033 29047 32091 29053
rect 32493 29053 32505 29056
rect 32539 29053 32551 29087
rect 32493 29047 32551 29053
rect 31444 28920 31984 28948
rect 31444 28908 31450 28920
rect 32030 28908 32036 28960
rect 32088 28948 32094 28960
rect 32125 28951 32183 28957
rect 32125 28948 32137 28951
rect 32088 28920 32137 28948
rect 32088 28908 32094 28920
rect 32125 28917 32137 28920
rect 32171 28917 32183 28951
rect 32508 28948 32536 29047
rect 32582 29044 32588 29096
rect 32640 29044 32646 29096
rect 33778 28976 33784 29028
rect 33836 28976 33842 29028
rect 33134 28948 33140 28960
rect 32508 28920 33140 28948
rect 32125 28911 32183 28917
rect 33134 28908 33140 28920
rect 33192 28908 33198 28960
rect 2760 28858 34316 28880
rect 2760 28806 7210 28858
rect 7262 28806 7274 28858
rect 7326 28806 7338 28858
rect 7390 28806 7402 28858
rect 7454 28806 7466 28858
rect 7518 28806 15099 28858
rect 15151 28806 15163 28858
rect 15215 28806 15227 28858
rect 15279 28806 15291 28858
rect 15343 28806 15355 28858
rect 15407 28806 22988 28858
rect 23040 28806 23052 28858
rect 23104 28806 23116 28858
rect 23168 28806 23180 28858
rect 23232 28806 23244 28858
rect 23296 28806 30877 28858
rect 30929 28806 30941 28858
rect 30993 28806 31005 28858
rect 31057 28806 31069 28858
rect 31121 28806 31133 28858
rect 31185 28806 34316 28858
rect 2760 28784 34316 28806
rect 5534 28744 5540 28756
rect 5184 28716 5540 28744
rect 5184 28676 5212 28716
rect 5534 28704 5540 28716
rect 5592 28744 5598 28756
rect 5592 28716 7604 28744
rect 5592 28704 5598 28716
rect 7576 28688 7604 28716
rect 7926 28704 7932 28756
rect 7984 28704 7990 28756
rect 8294 28704 8300 28756
rect 8352 28704 8358 28756
rect 8478 28704 8484 28756
rect 8536 28704 8542 28756
rect 10226 28704 10232 28756
rect 10284 28704 10290 28756
rect 10689 28747 10747 28753
rect 10689 28744 10701 28747
rect 10336 28716 10701 28744
rect 5092 28648 5212 28676
rect 1302 28568 1308 28620
rect 1360 28608 1366 28620
rect 3237 28611 3295 28617
rect 3237 28608 3249 28611
rect 1360 28580 3249 28608
rect 1360 28568 1366 28580
rect 3237 28577 3249 28580
rect 3283 28577 3295 28611
rect 3237 28571 3295 28577
rect 4430 28568 4436 28620
rect 4488 28568 4494 28620
rect 5092 28617 5120 28648
rect 7558 28636 7564 28688
rect 7616 28636 7622 28688
rect 5077 28611 5135 28617
rect 5077 28577 5089 28611
rect 5123 28577 5135 28611
rect 7745 28611 7803 28617
rect 7745 28608 7757 28611
rect 6486 28580 7757 28608
rect 5077 28571 5135 28577
rect 7745 28577 7757 28580
rect 7791 28577 7803 28611
rect 7745 28571 7803 28577
rect 7837 28611 7895 28617
rect 7837 28577 7849 28611
rect 7883 28608 7895 28611
rect 7944 28608 7972 28704
rect 10042 28636 10048 28688
rect 10100 28636 10106 28688
rect 10244 28676 10272 28704
rect 10336 28688 10364 28716
rect 10689 28713 10701 28716
rect 10735 28713 10747 28747
rect 10689 28707 10747 28713
rect 10778 28704 10784 28756
rect 10836 28744 10842 28756
rect 10962 28744 10968 28756
rect 10836 28716 10968 28744
rect 10836 28704 10842 28716
rect 10962 28704 10968 28716
rect 11020 28704 11026 28756
rect 13630 28704 13636 28756
rect 13688 28744 13694 28756
rect 14274 28744 14280 28756
rect 13688 28716 14280 28744
rect 13688 28704 13694 28716
rect 14274 28704 14280 28716
rect 14332 28744 14338 28756
rect 14461 28747 14519 28753
rect 14461 28744 14473 28747
rect 14332 28716 14473 28744
rect 14332 28704 14338 28716
rect 14461 28713 14473 28716
rect 14507 28713 14519 28747
rect 14461 28707 14519 28713
rect 14826 28704 14832 28756
rect 14884 28744 14890 28756
rect 15013 28747 15071 28753
rect 15013 28744 15025 28747
rect 14884 28716 15025 28744
rect 14884 28704 14890 28716
rect 15013 28713 15025 28716
rect 15059 28713 15071 28747
rect 16117 28747 16175 28753
rect 16117 28744 16129 28747
rect 15013 28707 15071 28713
rect 15488 28716 16129 28744
rect 10152 28648 10272 28676
rect 8202 28608 8208 28620
rect 7883 28580 8208 28608
rect 7883 28577 7895 28580
rect 7837 28571 7895 28577
rect 8202 28568 8208 28580
rect 8260 28568 8266 28620
rect 9125 28611 9183 28617
rect 9125 28577 9137 28611
rect 9171 28608 9183 28611
rect 9953 28611 10011 28617
rect 9953 28608 9965 28611
rect 9171 28580 9965 28608
rect 9171 28577 9183 28580
rect 9125 28571 9183 28577
rect 9953 28577 9965 28580
rect 9999 28577 10011 28611
rect 9953 28571 10011 28577
rect 5350 28500 5356 28552
rect 5408 28500 5414 28552
rect 6825 28543 6883 28549
rect 6825 28509 6837 28543
rect 6871 28540 6883 28543
rect 6917 28543 6975 28549
rect 6917 28540 6929 28543
rect 6871 28512 6929 28540
rect 6871 28509 6883 28512
rect 6825 28503 6883 28509
rect 6917 28509 6929 28512
rect 6963 28509 6975 28543
rect 6917 28503 6975 28509
rect 7006 28500 7012 28552
rect 7064 28540 7070 28552
rect 7561 28543 7619 28549
rect 7561 28540 7573 28543
rect 7064 28512 7573 28540
rect 7064 28500 7070 28512
rect 7561 28509 7573 28512
rect 7607 28509 7619 28543
rect 7561 28503 7619 28509
rect 9858 28500 9864 28552
rect 9916 28500 9922 28552
rect 10060 28540 10088 28636
rect 10152 28617 10180 28648
rect 10318 28636 10324 28688
rect 10376 28636 10382 28688
rect 10410 28636 10416 28688
rect 10468 28685 10474 28688
rect 10468 28679 10497 28685
rect 10485 28645 10497 28679
rect 12345 28679 12403 28685
rect 12345 28676 12357 28679
rect 10468 28639 10497 28645
rect 10704 28648 11560 28676
rect 10468 28636 10474 28639
rect 10704 28620 10732 28648
rect 10137 28611 10195 28617
rect 10137 28577 10149 28611
rect 10183 28577 10195 28611
rect 10137 28571 10195 28577
rect 10229 28611 10287 28617
rect 10229 28577 10241 28611
rect 10275 28577 10287 28611
rect 10229 28571 10287 28577
rect 10597 28611 10655 28617
rect 10597 28577 10609 28611
rect 10643 28608 10655 28611
rect 10686 28608 10692 28620
rect 10643 28580 10692 28608
rect 10643 28577 10655 28580
rect 10597 28571 10655 28577
rect 10244 28540 10272 28571
rect 10686 28568 10692 28580
rect 10744 28568 10750 28620
rect 10781 28611 10839 28617
rect 10781 28577 10793 28611
rect 10827 28577 10839 28611
rect 10781 28571 10839 28577
rect 10060 28512 10272 28540
rect 10502 28500 10508 28552
rect 10560 28540 10566 28552
rect 10796 28540 10824 28571
rect 10962 28568 10968 28620
rect 11020 28608 11026 28620
rect 11330 28608 11336 28620
rect 11020 28580 11336 28608
rect 11020 28568 11026 28580
rect 11330 28568 11336 28580
rect 11388 28608 11394 28620
rect 11532 28617 11560 28648
rect 11624 28648 12357 28676
rect 11425 28611 11483 28617
rect 11425 28608 11437 28611
rect 11388 28580 11437 28608
rect 11388 28568 11394 28580
rect 11425 28577 11437 28580
rect 11471 28577 11483 28611
rect 11425 28571 11483 28577
rect 11517 28611 11575 28617
rect 11517 28577 11529 28611
rect 11563 28577 11575 28611
rect 11517 28571 11575 28577
rect 11624 28540 11652 28648
rect 12345 28645 12357 28648
rect 12391 28645 12403 28679
rect 15381 28679 15439 28685
rect 15381 28676 15393 28679
rect 12345 28639 12403 28645
rect 14660 28648 15393 28676
rect 11885 28611 11943 28617
rect 11885 28577 11897 28611
rect 11931 28577 11943 28611
rect 11885 28571 11943 28577
rect 12621 28611 12679 28617
rect 12621 28577 12633 28611
rect 12667 28608 12679 28611
rect 13630 28608 13636 28620
rect 12667 28580 13636 28608
rect 12667 28577 12679 28580
rect 12621 28571 12679 28577
rect 10560 28512 11652 28540
rect 10560 28500 10566 28512
rect 10594 28432 10600 28484
rect 10652 28472 10658 28484
rect 11900 28472 11928 28571
rect 13630 28568 13636 28580
rect 13688 28568 13694 28620
rect 14660 28617 14688 28648
rect 15381 28645 15393 28648
rect 15427 28645 15439 28679
rect 15381 28639 15439 28645
rect 14645 28611 14703 28617
rect 14645 28577 14657 28611
rect 14691 28577 14703 28611
rect 14645 28571 14703 28577
rect 14734 28568 14740 28620
rect 14792 28568 14798 28620
rect 14918 28568 14924 28620
rect 14976 28568 14982 28620
rect 15010 28568 15016 28620
rect 15068 28608 15074 28620
rect 15105 28611 15163 28617
rect 15105 28608 15117 28611
rect 15068 28580 15117 28608
rect 15068 28568 15074 28580
rect 15105 28577 15117 28580
rect 15151 28608 15163 28611
rect 15488 28608 15516 28716
rect 16117 28713 16129 28716
rect 16163 28713 16175 28747
rect 16117 28707 16175 28713
rect 16574 28704 16580 28756
rect 16632 28704 16638 28756
rect 17126 28704 17132 28756
rect 17184 28704 17190 28756
rect 17954 28704 17960 28756
rect 18012 28744 18018 28756
rect 18325 28747 18383 28753
rect 18325 28744 18337 28747
rect 18012 28716 18337 28744
rect 18012 28704 18018 28716
rect 18325 28713 18337 28716
rect 18371 28713 18383 28747
rect 18325 28707 18383 28713
rect 19076 28716 19472 28744
rect 16485 28679 16543 28685
rect 16485 28676 16497 28679
rect 15151 28580 15516 28608
rect 15580 28648 16497 28676
rect 15151 28577 15163 28580
rect 15105 28571 15163 28577
rect 12434 28500 12440 28552
rect 12492 28500 12498 28552
rect 13725 28543 13783 28549
rect 13725 28540 13737 28543
rect 12820 28512 13737 28540
rect 12820 28481 12848 28512
rect 13725 28509 13737 28512
rect 13771 28509 13783 28543
rect 13725 28503 13783 28509
rect 15289 28543 15347 28549
rect 15289 28509 15301 28543
rect 15335 28540 15347 28543
rect 15470 28540 15476 28552
rect 15335 28512 15476 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 15470 28500 15476 28512
rect 15528 28500 15534 28552
rect 10652 28444 11928 28472
rect 12069 28475 12127 28481
rect 10652 28432 10658 28444
rect 12069 28441 12081 28475
rect 12115 28472 12127 28475
rect 12805 28475 12863 28481
rect 12115 28444 12756 28472
rect 12115 28441 12127 28444
rect 12069 28435 12127 28441
rect 9214 28364 9220 28416
rect 9272 28364 9278 28416
rect 10870 28364 10876 28416
rect 10928 28404 10934 28416
rect 11606 28404 11612 28416
rect 10928 28376 11612 28404
rect 10928 28364 10934 28376
rect 11606 28364 11612 28376
rect 11664 28404 11670 28416
rect 11793 28407 11851 28413
rect 11793 28404 11805 28407
rect 11664 28376 11805 28404
rect 11664 28364 11670 28376
rect 11793 28373 11805 28376
rect 11839 28373 11851 28407
rect 11793 28367 11851 28373
rect 12618 28364 12624 28416
rect 12676 28364 12682 28416
rect 12728 28404 12756 28444
rect 12805 28441 12817 28475
rect 12851 28441 12863 28475
rect 12805 28435 12863 28441
rect 12912 28444 13400 28472
rect 12912 28404 12940 28444
rect 13372 28416 13400 28444
rect 13814 28432 13820 28484
rect 13872 28472 13878 28484
rect 14366 28472 14372 28484
rect 13872 28444 14372 28472
rect 13872 28432 13878 28444
rect 14366 28432 14372 28444
rect 14424 28432 14430 28484
rect 12728 28376 12940 28404
rect 13170 28364 13176 28416
rect 13228 28364 13234 28416
rect 13354 28364 13360 28416
rect 13412 28364 13418 28416
rect 13906 28364 13912 28416
rect 13964 28404 13970 28416
rect 15580 28404 15608 28648
rect 16485 28645 16497 28648
rect 16531 28645 16543 28679
rect 16485 28639 16543 28645
rect 15838 28568 15844 28620
rect 15896 28608 15902 28620
rect 16301 28611 16359 28617
rect 16301 28608 16313 28611
rect 15896 28580 16313 28608
rect 15896 28568 15902 28580
rect 16301 28577 16313 28580
rect 16347 28577 16359 28611
rect 16301 28571 16359 28577
rect 16390 28568 16396 28620
rect 16448 28568 16454 28620
rect 16592 28608 16620 28704
rect 18141 28679 18199 28685
rect 18141 28645 18153 28679
rect 18187 28676 18199 28679
rect 19076 28676 19104 28716
rect 18187 28648 19104 28676
rect 18187 28645 18199 28648
rect 18141 28639 18199 28645
rect 19150 28636 19156 28688
rect 19208 28676 19214 28688
rect 19444 28685 19472 28716
rect 21542 28704 21548 28756
rect 21600 28704 21606 28756
rect 21928 28716 22784 28744
rect 21928 28688 21956 28716
rect 19337 28679 19395 28685
rect 19337 28676 19349 28679
rect 19208 28648 19349 28676
rect 19208 28636 19214 28648
rect 19337 28645 19349 28648
rect 19383 28645 19395 28679
rect 19337 28639 19395 28645
rect 19429 28679 19487 28685
rect 19429 28645 19441 28679
rect 19475 28676 19487 28679
rect 19702 28676 19708 28688
rect 19475 28648 19708 28676
rect 19475 28645 19487 28648
rect 19429 28639 19487 28645
rect 19702 28636 19708 28648
rect 19760 28636 19766 28688
rect 21910 28636 21916 28688
rect 21968 28636 21974 28688
rect 22554 28636 22560 28688
rect 22612 28636 22618 28688
rect 17221 28611 17279 28617
rect 17221 28608 17233 28611
rect 16592 28580 17233 28608
rect 17221 28577 17233 28580
rect 17267 28577 17279 28611
rect 17221 28571 17279 28577
rect 19242 28568 19248 28620
rect 19300 28568 19306 28620
rect 19610 28568 19616 28620
rect 19668 28568 19674 28620
rect 21082 28568 21088 28620
rect 21140 28608 21146 28620
rect 22465 28611 22523 28617
rect 22465 28608 22477 28611
rect 21140 28580 22477 28608
rect 21140 28568 21146 28580
rect 22465 28577 22477 28580
rect 22511 28608 22523 28611
rect 22511 28580 22600 28608
rect 22511 28577 22523 28580
rect 22465 28571 22523 28577
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28540 16083 28543
rect 18969 28543 19027 28549
rect 16071 28512 16436 28540
rect 16071 28509 16083 28512
rect 16025 28503 16083 28509
rect 16408 28472 16436 28512
rect 18969 28509 18981 28543
rect 19015 28540 19027 28543
rect 22189 28543 22247 28549
rect 19015 28512 19104 28540
rect 19015 28509 19027 28512
rect 18969 28503 19027 28509
rect 19076 28481 19104 28512
rect 22189 28509 22201 28543
rect 22235 28540 22247 28543
rect 22235 28512 22324 28540
rect 22235 28509 22247 28512
rect 22189 28503 22247 28509
rect 22296 28481 22324 28512
rect 16669 28475 16727 28481
rect 16669 28472 16681 28475
rect 16408 28444 16681 28472
rect 16669 28441 16681 28444
rect 16715 28472 16727 28475
rect 19061 28475 19119 28481
rect 16715 28444 17540 28472
rect 16715 28441 16727 28444
rect 16669 28435 16727 28441
rect 17512 28416 17540 28444
rect 19061 28441 19073 28475
rect 19107 28441 19119 28475
rect 19061 28435 19119 28441
rect 22281 28475 22339 28481
rect 22281 28441 22293 28475
rect 22327 28441 22339 28475
rect 22572 28472 22600 28580
rect 22646 28568 22652 28620
rect 22704 28568 22710 28620
rect 22756 28608 22784 28716
rect 22830 28704 22836 28756
rect 22888 28744 22894 28756
rect 23017 28747 23075 28753
rect 23017 28744 23029 28747
rect 22888 28716 23029 28744
rect 22888 28704 22894 28716
rect 23017 28713 23029 28716
rect 23063 28713 23075 28747
rect 23017 28707 23075 28713
rect 23382 28704 23388 28756
rect 23440 28704 23446 28756
rect 27246 28704 27252 28756
rect 27304 28744 27310 28756
rect 27433 28747 27491 28753
rect 27433 28744 27445 28747
rect 27304 28716 27445 28744
rect 27304 28704 27310 28716
rect 27433 28713 27445 28716
rect 27479 28713 27491 28747
rect 27433 28707 27491 28713
rect 27798 28704 27804 28756
rect 27856 28704 27862 28756
rect 28258 28704 28264 28756
rect 28316 28704 28322 28756
rect 28813 28747 28871 28753
rect 28813 28713 28825 28747
rect 28859 28744 28871 28747
rect 28994 28744 29000 28756
rect 28859 28716 29000 28744
rect 28859 28713 28871 28716
rect 28813 28707 28871 28713
rect 28994 28704 29000 28716
rect 29052 28704 29058 28756
rect 30929 28747 30987 28753
rect 30929 28713 30941 28747
rect 30975 28744 30987 28747
rect 31202 28744 31208 28756
rect 30975 28716 31208 28744
rect 30975 28713 30987 28716
rect 30929 28707 30987 28713
rect 31202 28704 31208 28716
rect 31260 28704 31266 28756
rect 22830 28608 22836 28620
rect 22756 28580 22836 28608
rect 22830 28568 22836 28580
rect 22888 28568 22894 28620
rect 23109 28611 23167 28617
rect 23109 28577 23121 28611
rect 23155 28608 23167 28611
rect 23400 28608 23428 28704
rect 23474 28636 23480 28688
rect 23532 28636 23538 28688
rect 24670 28636 24676 28688
rect 24728 28636 24734 28688
rect 26878 28636 26884 28688
rect 26936 28636 26942 28688
rect 27709 28679 27767 28685
rect 27448 28648 27660 28676
rect 27448 28620 27476 28648
rect 23155 28580 23428 28608
rect 23155 28577 23167 28580
rect 23109 28571 23167 28577
rect 27430 28568 27436 28620
rect 27488 28568 27494 28620
rect 27522 28568 27528 28620
rect 27580 28568 27586 28620
rect 27632 28617 27660 28648
rect 27709 28645 27721 28679
rect 27755 28676 27767 28679
rect 27816 28676 27844 28704
rect 27755 28648 27844 28676
rect 27755 28645 27767 28648
rect 27709 28639 27767 28645
rect 27617 28611 27675 28617
rect 27617 28577 27629 28611
rect 27663 28577 27675 28611
rect 27617 28571 27675 28577
rect 27798 28568 27804 28620
rect 27856 28568 27862 28620
rect 27890 28568 27896 28620
rect 27948 28608 27954 28620
rect 27985 28611 28043 28617
rect 27985 28608 27997 28611
rect 27948 28580 27997 28608
rect 27948 28568 27954 28580
rect 27985 28577 27997 28580
rect 28031 28577 28043 28611
rect 28276 28608 28304 28704
rect 31294 28636 31300 28688
rect 31352 28636 31358 28688
rect 32030 28636 32036 28688
rect 32088 28636 32094 28688
rect 28626 28608 28632 28620
rect 28276 28580 28632 28608
rect 27985 28571 28043 28577
rect 28626 28568 28632 28580
rect 28684 28608 28690 28620
rect 28721 28611 28779 28617
rect 28721 28608 28733 28611
rect 28684 28580 28733 28608
rect 28684 28568 28690 28580
rect 28721 28577 28733 28580
rect 28767 28577 28779 28611
rect 28721 28571 28779 28577
rect 30558 28568 30564 28620
rect 30616 28568 30622 28620
rect 33134 28568 33140 28620
rect 33192 28608 33198 28620
rect 33781 28611 33839 28617
rect 33781 28608 33793 28611
rect 33192 28580 33793 28608
rect 33192 28568 33198 28580
rect 33781 28577 33793 28580
rect 33827 28577 33839 28611
rect 33781 28571 33839 28577
rect 24762 28540 24768 28552
rect 22756 28512 24768 28540
rect 22756 28472 22784 28512
rect 24762 28500 24768 28512
rect 24820 28500 24826 28552
rect 25222 28500 25228 28552
rect 25280 28500 25286 28552
rect 25501 28543 25559 28549
rect 25501 28509 25513 28543
rect 25547 28540 25559 28543
rect 25593 28543 25651 28549
rect 25593 28540 25605 28543
rect 25547 28512 25605 28540
rect 25547 28509 25559 28512
rect 25501 28503 25559 28509
rect 25593 28509 25605 28512
rect 25639 28509 25651 28543
rect 25593 28503 25651 28509
rect 22572 28444 22784 28472
rect 22281 28435 22339 28441
rect 13964 28376 15608 28404
rect 13964 28364 13970 28376
rect 17494 28364 17500 28416
rect 17552 28364 17558 28416
rect 24026 28364 24032 28416
rect 24084 28404 24090 28416
rect 25516 28404 25544 28503
rect 25866 28500 25872 28552
rect 25924 28500 25930 28552
rect 27540 28540 27568 28568
rect 29178 28540 29184 28552
rect 27540 28512 29184 28540
rect 29178 28500 29184 28512
rect 29236 28500 29242 28552
rect 29454 28500 29460 28552
rect 29512 28500 29518 28552
rect 30650 28540 30656 28552
rect 30484 28512 30656 28540
rect 27341 28475 27399 28481
rect 27341 28441 27353 28475
rect 27387 28472 27399 28475
rect 28442 28472 28448 28484
rect 27387 28444 28448 28472
rect 27387 28441 27399 28444
rect 27341 28435 27399 28441
rect 28442 28432 28448 28444
rect 28500 28432 28506 28484
rect 24084 28376 25544 28404
rect 24084 28364 24090 28376
rect 27798 28364 27804 28416
rect 27856 28404 27862 28416
rect 28261 28407 28319 28413
rect 28261 28404 28273 28407
rect 27856 28376 28273 28404
rect 27856 28364 27862 28376
rect 28261 28373 28273 28376
rect 28307 28373 28319 28407
rect 29196 28404 29224 28500
rect 30484 28404 30512 28512
rect 30650 28500 30656 28512
rect 30708 28540 30714 28552
rect 31018 28540 31024 28552
rect 30708 28512 31024 28540
rect 30708 28500 30714 28512
rect 31018 28500 31024 28512
rect 31076 28500 31082 28552
rect 33410 28500 33416 28552
rect 33468 28500 33474 28552
rect 29196 28376 30512 28404
rect 28261 28367 28319 28373
rect 32306 28364 32312 28416
rect 32364 28404 32370 28416
rect 32582 28404 32588 28416
rect 32364 28376 32588 28404
rect 32364 28364 32370 28376
rect 32582 28364 32588 28376
rect 32640 28404 32646 28416
rect 32769 28407 32827 28413
rect 32769 28404 32781 28407
rect 32640 28376 32781 28404
rect 32640 28364 32646 28376
rect 32769 28373 32781 28376
rect 32815 28373 32827 28407
rect 32769 28367 32827 28373
rect 32858 28364 32864 28416
rect 32916 28364 32922 28416
rect 33870 28364 33876 28416
rect 33928 28364 33934 28416
rect 2760 28314 34316 28336
rect 2760 28262 6550 28314
rect 6602 28262 6614 28314
rect 6666 28262 6678 28314
rect 6730 28262 6742 28314
rect 6794 28262 6806 28314
rect 6858 28262 14439 28314
rect 14491 28262 14503 28314
rect 14555 28262 14567 28314
rect 14619 28262 14631 28314
rect 14683 28262 14695 28314
rect 14747 28262 22328 28314
rect 22380 28262 22392 28314
rect 22444 28262 22456 28314
rect 22508 28262 22520 28314
rect 22572 28262 22584 28314
rect 22636 28262 30217 28314
rect 30269 28262 30281 28314
rect 30333 28262 30345 28314
rect 30397 28262 30409 28314
rect 30461 28262 30473 28314
rect 30525 28262 34316 28314
rect 2760 28240 34316 28262
rect 5261 28203 5319 28209
rect 5261 28169 5273 28203
rect 5307 28200 5319 28203
rect 5350 28200 5356 28212
rect 5307 28172 5356 28200
rect 5307 28169 5319 28172
rect 5261 28163 5319 28169
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 7732 28203 7790 28209
rect 7732 28169 7744 28203
rect 7778 28200 7790 28203
rect 9214 28200 9220 28212
rect 7778 28172 9220 28200
rect 7778 28169 7790 28172
rect 7732 28163 7790 28169
rect 9214 28160 9220 28172
rect 9272 28160 9278 28212
rect 9858 28160 9864 28212
rect 9916 28200 9922 28212
rect 10597 28203 10655 28209
rect 10597 28200 10609 28203
rect 9916 28172 10609 28200
rect 9916 28160 9922 28172
rect 10597 28169 10609 28172
rect 10643 28169 10655 28203
rect 10597 28163 10655 28169
rect 12069 28203 12127 28209
rect 12069 28169 12081 28203
rect 12115 28200 12127 28203
rect 12434 28200 12440 28212
rect 12115 28172 12440 28200
rect 12115 28169 12127 28172
rect 12069 28163 12127 28169
rect 12434 28160 12440 28172
rect 12492 28160 12498 28212
rect 12986 28160 12992 28212
rect 13044 28160 13050 28212
rect 13170 28160 13176 28212
rect 13228 28160 13234 28212
rect 13541 28203 13599 28209
rect 13541 28169 13553 28203
rect 13587 28200 13599 28203
rect 13633 28203 13691 28209
rect 13633 28200 13645 28203
rect 13587 28172 13645 28200
rect 13587 28169 13599 28172
rect 13541 28163 13599 28169
rect 13633 28169 13645 28172
rect 13679 28169 13691 28203
rect 13633 28163 13691 28169
rect 14090 28160 14096 28212
rect 14148 28160 14154 28212
rect 15746 28200 15752 28212
rect 14292 28172 15752 28200
rect 9953 28135 10011 28141
rect 9953 28101 9965 28135
rect 9999 28101 10011 28135
rect 9953 28095 10011 28101
rect 10873 28135 10931 28141
rect 10873 28101 10885 28135
rect 10919 28132 10931 28135
rect 11974 28132 11980 28144
rect 10919 28104 11980 28132
rect 10919 28101 10931 28104
rect 10873 28095 10931 28101
rect 7834 28064 7840 28076
rect 5644 28036 7840 28064
rect 3970 27956 3976 28008
rect 4028 27956 4034 28008
rect 5644 28005 5672 28036
rect 7834 28024 7840 28036
rect 7892 28024 7898 28076
rect 9217 28067 9275 28073
rect 9217 28033 9229 28067
rect 9263 28064 9275 28067
rect 9263 28036 9812 28064
rect 9263 28033 9275 28036
rect 9217 28027 9275 28033
rect 9784 28005 9812 28036
rect 4709 27999 4767 28005
rect 4709 27965 4721 27999
rect 4755 27965 4767 27999
rect 4709 27959 4767 27965
rect 5629 27999 5687 28005
rect 5629 27965 5641 27999
rect 5675 27965 5687 27999
rect 5629 27959 5687 27965
rect 7469 27999 7527 28005
rect 7469 27965 7481 27999
rect 7515 27965 7527 27999
rect 7469 27959 7527 27965
rect 9769 27999 9827 28005
rect 9769 27965 9781 27999
rect 9815 27965 9827 27999
rect 9968 27996 9996 28095
rect 11974 28092 11980 28104
rect 12032 28132 12038 28144
rect 12250 28132 12256 28144
rect 12032 28104 12256 28132
rect 12032 28092 12038 28104
rect 12250 28092 12256 28104
rect 12308 28092 12314 28144
rect 10965 28067 11023 28073
rect 10965 28033 10977 28067
rect 11011 28064 11023 28067
rect 11146 28064 11152 28076
rect 11011 28036 11152 28064
rect 11011 28033 11023 28036
rect 10965 28027 11023 28033
rect 11146 28024 11152 28036
rect 11204 28024 11210 28076
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28064 12955 28067
rect 13188 28064 13216 28160
rect 12943 28036 13216 28064
rect 12943 28033 12955 28036
rect 12897 28027 12955 28033
rect 13354 28024 13360 28076
rect 13412 28024 13418 28076
rect 13630 28024 13636 28076
rect 13688 28064 13694 28076
rect 13909 28067 13967 28073
rect 13909 28064 13921 28067
rect 13688 28036 13921 28064
rect 13688 28024 13694 28036
rect 13909 28033 13921 28036
rect 13955 28064 13967 28067
rect 14292 28064 14320 28172
rect 15746 28160 15752 28172
rect 15804 28200 15810 28212
rect 16390 28200 16396 28212
rect 15804 28172 16396 28200
rect 15804 28160 15810 28172
rect 16390 28160 16396 28172
rect 16448 28160 16454 28212
rect 17494 28160 17500 28212
rect 17552 28160 17558 28212
rect 20898 28160 20904 28212
rect 20956 28200 20962 28212
rect 23382 28200 23388 28212
rect 20956 28172 23388 28200
rect 20956 28160 20962 28172
rect 23382 28160 23388 28172
rect 23440 28160 23446 28212
rect 24026 28160 24032 28212
rect 24084 28200 24090 28212
rect 24213 28203 24271 28209
rect 24213 28200 24225 28203
rect 24084 28172 24225 28200
rect 24084 28160 24090 28172
rect 24213 28169 24225 28172
rect 24259 28169 24271 28203
rect 24213 28163 24271 28169
rect 24688 28172 25176 28200
rect 22830 28092 22836 28144
rect 22888 28132 22894 28144
rect 24688 28132 24716 28172
rect 22888 28104 24716 28132
rect 25148 28132 25176 28172
rect 25222 28160 25228 28212
rect 25280 28200 25286 28212
rect 25409 28203 25467 28209
rect 25409 28200 25421 28203
rect 25280 28172 25421 28200
rect 25280 28160 25286 28172
rect 25409 28169 25421 28172
rect 25455 28169 25467 28203
rect 25409 28163 25467 28169
rect 25866 28160 25872 28212
rect 25924 28200 25930 28212
rect 26053 28203 26111 28209
rect 26053 28200 26065 28203
rect 25924 28172 26065 28200
rect 25924 28160 25930 28172
rect 26053 28169 26065 28172
rect 26099 28169 26111 28203
rect 26053 28163 26111 28169
rect 26789 28203 26847 28209
rect 26789 28169 26801 28203
rect 26835 28200 26847 28203
rect 26878 28200 26884 28212
rect 26835 28172 26884 28200
rect 26835 28169 26847 28172
rect 26789 28163 26847 28169
rect 26878 28160 26884 28172
rect 26936 28160 26942 28212
rect 28350 28160 28356 28212
rect 28408 28200 28414 28212
rect 28810 28200 28816 28212
rect 28408 28172 28816 28200
rect 28408 28160 28414 28172
rect 28810 28160 28816 28172
rect 28868 28200 28874 28212
rect 29181 28203 29239 28209
rect 29181 28200 29193 28203
rect 28868 28172 29193 28200
rect 28868 28160 28874 28172
rect 29181 28169 29193 28172
rect 29227 28169 29239 28203
rect 29181 28163 29239 28169
rect 29270 28160 29276 28212
rect 29328 28160 29334 28212
rect 29454 28160 29460 28212
rect 29512 28200 29518 28212
rect 29917 28203 29975 28209
rect 29917 28200 29929 28203
rect 29512 28172 29929 28200
rect 29512 28160 29518 28172
rect 29917 28169 29929 28172
rect 29963 28169 29975 28203
rect 29917 28163 29975 28169
rect 31205 28203 31263 28209
rect 31205 28169 31217 28203
rect 31251 28200 31263 28203
rect 31846 28200 31852 28212
rect 31251 28172 31852 28200
rect 31251 28169 31263 28172
rect 31205 28163 31263 28169
rect 31846 28160 31852 28172
rect 31904 28160 31910 28212
rect 25148 28104 26556 28132
rect 22888 28092 22894 28104
rect 13955 28036 14320 28064
rect 13955 28033 13967 28036
rect 13909 28027 13967 28033
rect 14366 28024 14372 28076
rect 14424 28024 14430 28076
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28064 15807 28067
rect 15795 28036 17724 28064
rect 15795 28033 15807 28036
rect 15749 28027 15807 28033
rect 17696 28008 17724 28036
rect 25038 28024 25044 28076
rect 25096 28064 25102 28076
rect 26528 28064 26556 28104
rect 28902 28092 28908 28144
rect 28960 28132 28966 28144
rect 29288 28132 29316 28160
rect 28960 28104 29316 28132
rect 28960 28092 28966 28104
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 25096 28036 26464 28064
rect 25096 28024 25102 28036
rect 10781 27999 10839 28005
rect 10781 27996 10793 27999
rect 9968 27968 10793 27996
rect 9769 27959 9827 27965
rect 10781 27965 10793 27968
rect 10827 27996 10839 27999
rect 10870 27996 10876 28008
rect 10827 27968 10876 27996
rect 10827 27965 10839 27968
rect 10781 27959 10839 27965
rect 4724 27928 4752 27959
rect 6730 27928 6736 27940
rect 4724 27900 6736 27928
rect 6730 27888 6736 27900
rect 6788 27888 6794 27940
rect 7377 27931 7435 27937
rect 7377 27897 7389 27931
rect 7423 27928 7435 27931
rect 7484 27928 7512 27959
rect 7423 27900 7512 27928
rect 7423 27897 7435 27900
rect 7377 27891 7435 27897
rect 4522 27820 4528 27872
rect 4580 27820 4586 27872
rect 7484 27860 7512 27900
rect 8386 27888 8392 27940
rect 8444 27888 8450 27940
rect 9784 27928 9812 27959
rect 10870 27956 10876 27968
rect 10928 27956 10934 28008
rect 11057 27999 11115 28005
rect 11057 27965 11069 27999
rect 11103 27965 11115 27999
rect 11057 27959 11115 27965
rect 10502 27928 10508 27940
rect 9784 27900 10508 27928
rect 10502 27888 10508 27900
rect 10560 27888 10566 27940
rect 11072 27928 11100 27959
rect 11238 27956 11244 28008
rect 11296 27956 11302 28008
rect 11422 27956 11428 28008
rect 11480 27956 11486 28008
rect 12713 27999 12771 28005
rect 12713 27965 12725 27999
rect 12759 27996 12771 27999
rect 13262 27996 13268 28008
rect 12759 27968 13268 27996
rect 12759 27965 12771 27968
rect 12713 27959 12771 27965
rect 13262 27956 13268 27968
rect 13320 27956 13326 28008
rect 13538 27956 13544 28008
rect 13596 27956 13602 28008
rect 13817 27999 13875 28005
rect 13817 27965 13829 27999
rect 13863 27965 13875 27999
rect 13817 27959 13875 27965
rect 11330 27928 11336 27940
rect 11072 27900 11336 27928
rect 11330 27888 11336 27900
rect 11388 27888 11394 27940
rect 12894 27888 12900 27940
rect 12952 27928 12958 27940
rect 12989 27931 13047 27937
rect 12989 27928 13001 27931
rect 12952 27900 13001 27928
rect 12952 27888 12958 27900
rect 12989 27897 13001 27900
rect 13035 27897 13047 27931
rect 13832 27928 13860 27959
rect 13998 27956 14004 28008
rect 14056 27956 14062 28008
rect 14274 27956 14280 28008
rect 14332 27996 14338 28008
rect 14553 27999 14611 28005
rect 14553 27996 14565 27999
rect 14332 27968 14565 27996
rect 14332 27956 14338 27968
rect 14553 27965 14565 27968
rect 14599 27965 14611 27999
rect 14553 27959 14611 27965
rect 17678 27956 17684 28008
rect 17736 27956 17742 28008
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27996 19671 27999
rect 20070 27996 20076 28008
rect 19659 27968 20076 27996
rect 19659 27965 19671 27968
rect 19613 27959 19671 27965
rect 20070 27956 20076 27968
rect 20128 27956 20134 28008
rect 20898 27956 20904 28008
rect 20956 27996 20962 28008
rect 21085 27999 21143 28005
rect 21085 27996 21097 27999
rect 20956 27968 21097 27996
rect 20956 27956 20962 27968
rect 21085 27965 21097 27968
rect 21131 27965 21143 27999
rect 21085 27959 21143 27965
rect 24210 27956 24216 28008
rect 24268 27996 24274 28008
rect 24765 27999 24823 28005
rect 24765 27996 24777 27999
rect 24268 27968 24777 27996
rect 24268 27956 24274 27968
rect 24765 27965 24777 27968
rect 24811 27965 24823 27999
rect 26142 27996 26148 28008
rect 24765 27959 24823 27965
rect 25700 27968 26148 27996
rect 14016 27928 14044 27956
rect 13832 27900 14044 27928
rect 14093 27931 14151 27937
rect 12989 27891 13047 27897
rect 14093 27897 14105 27931
rect 14139 27928 14151 27931
rect 15470 27928 15476 27940
rect 14139 27900 15476 27928
rect 14139 27897 14151 27900
rect 14093 27891 14151 27897
rect 15470 27888 15476 27900
rect 15528 27888 15534 27940
rect 16022 27888 16028 27940
rect 16080 27888 16086 27940
rect 16758 27888 16764 27940
rect 16816 27888 16822 27940
rect 22925 27931 22983 27937
rect 22925 27928 22937 27931
rect 22756 27900 22937 27928
rect 7558 27860 7564 27872
rect 7484 27832 7564 27860
rect 7558 27820 7564 27832
rect 7616 27860 7622 27872
rect 8018 27860 8024 27872
rect 7616 27832 8024 27860
rect 7616 27820 7622 27832
rect 8018 27820 8024 27832
rect 8076 27820 8082 27872
rect 11698 27820 11704 27872
rect 11756 27860 11762 27872
rect 12529 27863 12587 27869
rect 12529 27860 12541 27863
rect 11756 27832 12541 27860
rect 11756 27820 11762 27832
rect 12529 27829 12541 27832
rect 12575 27829 12587 27863
rect 12529 27823 12587 27829
rect 13078 27820 13084 27872
rect 13136 27820 13142 27872
rect 13814 27820 13820 27872
rect 13872 27860 13878 27872
rect 13998 27860 14004 27872
rect 13872 27832 14004 27860
rect 13872 27820 13878 27832
rect 13998 27820 14004 27832
rect 14056 27820 14062 27872
rect 14642 27820 14648 27872
rect 14700 27820 14706 27872
rect 15013 27863 15071 27869
rect 15013 27829 15025 27863
rect 15059 27860 15071 27863
rect 15562 27860 15568 27872
rect 15059 27832 15568 27860
rect 15059 27829 15071 27832
rect 15013 27823 15071 27829
rect 15562 27820 15568 27832
rect 15620 27820 15626 27872
rect 17770 27820 17776 27872
rect 17828 27820 17834 27872
rect 18046 27820 18052 27872
rect 18104 27860 18110 27872
rect 18969 27863 19027 27869
rect 18969 27860 18981 27863
rect 18104 27832 18981 27860
rect 18104 27820 18110 27832
rect 18969 27829 18981 27832
rect 19015 27829 19027 27863
rect 18969 27823 19027 27829
rect 20990 27820 20996 27872
rect 21048 27820 21054 27872
rect 21910 27820 21916 27872
rect 21968 27820 21974 27872
rect 22186 27820 22192 27872
rect 22244 27860 22250 27872
rect 22281 27863 22339 27869
rect 22281 27860 22293 27863
rect 22244 27832 22293 27860
rect 22244 27820 22250 27832
rect 22281 27829 22293 27832
rect 22327 27860 22339 27863
rect 22554 27860 22560 27872
rect 22327 27832 22560 27860
rect 22327 27829 22339 27832
rect 22281 27823 22339 27829
rect 22554 27820 22560 27832
rect 22612 27820 22618 27872
rect 22646 27820 22652 27872
rect 22704 27860 22710 27872
rect 22756 27869 22784 27900
rect 22925 27897 22937 27900
rect 22971 27897 22983 27931
rect 22925 27891 22983 27897
rect 22741 27863 22799 27869
rect 22741 27860 22753 27863
rect 22704 27832 22753 27860
rect 22704 27820 22710 27832
rect 22741 27829 22753 27832
rect 22787 27829 22799 27863
rect 22741 27823 22799 27829
rect 25130 27820 25136 27872
rect 25188 27860 25194 27872
rect 25700 27869 25728 27968
rect 26142 27956 26148 27968
rect 26200 27996 26206 28008
rect 26436 28005 26464 28036
rect 26528 28036 27169 28064
rect 26237 27999 26295 28005
rect 26237 27996 26249 27999
rect 26200 27968 26249 27996
rect 26200 27956 26206 27968
rect 26237 27965 26249 27968
rect 26283 27965 26295 27999
rect 26237 27959 26295 27965
rect 26421 27999 26479 28005
rect 26421 27965 26433 27999
rect 26467 27965 26479 27999
rect 26528 27996 26556 28036
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 29089 28067 29147 28073
rect 29089 28033 29101 28067
rect 29135 28064 29147 28067
rect 29733 28067 29791 28073
rect 29733 28064 29745 28067
rect 29135 28036 29745 28064
rect 29135 28033 29147 28036
rect 29089 28027 29147 28033
rect 29733 28033 29745 28036
rect 29779 28033 29791 28067
rect 31386 28064 31392 28076
rect 29733 28027 29791 28033
rect 30024 28036 31392 28064
rect 30024 28008 30052 28036
rect 26605 27999 26663 28005
rect 26605 27996 26617 27999
rect 26528 27968 26617 27996
rect 26421 27959 26479 27965
rect 26605 27965 26617 27968
rect 26651 27965 26663 27999
rect 26605 27959 26663 27965
rect 26694 27956 26700 28008
rect 26752 27956 26758 28008
rect 27341 27999 27399 28005
rect 27341 27965 27353 27999
rect 27387 27965 27399 27999
rect 27341 27959 27399 27965
rect 26329 27931 26387 27937
rect 26329 27897 26341 27931
rect 26375 27928 26387 27931
rect 27356 27928 27384 27959
rect 28718 27956 28724 28008
rect 28776 27956 28782 28008
rect 30006 27956 30012 28008
rect 30064 27956 30070 28008
rect 30374 27956 30380 28008
rect 30432 27996 30438 28008
rect 30852 28005 30880 28036
rect 31386 28024 31392 28036
rect 31444 28024 31450 28076
rect 31662 28024 31668 28076
rect 31720 28064 31726 28076
rect 31757 28067 31815 28073
rect 31757 28064 31769 28067
rect 31720 28036 31769 28064
rect 31720 28024 31726 28036
rect 31757 28033 31769 28036
rect 31803 28033 31815 28067
rect 31757 28027 31815 28033
rect 32401 28067 32459 28073
rect 32401 28033 32413 28067
rect 32447 28064 32459 28067
rect 32858 28064 32864 28076
rect 32447 28036 32864 28064
rect 32447 28033 32459 28036
rect 32401 28027 32459 28033
rect 32858 28024 32864 28036
rect 32916 28024 32922 28076
rect 30469 27999 30527 28005
rect 30469 27996 30481 27999
rect 30432 27968 30481 27996
rect 30432 27956 30438 27968
rect 30469 27965 30481 27968
rect 30515 27965 30527 27999
rect 30469 27959 30527 27965
rect 30837 27999 30895 28005
rect 30837 27965 30849 27999
rect 30883 27965 30895 27999
rect 30837 27959 30895 27965
rect 31018 27956 31024 28008
rect 31076 27996 31082 28008
rect 32125 27999 32183 28005
rect 32125 27996 32137 27999
rect 31076 27968 32137 27996
rect 31076 27956 31082 27968
rect 32125 27965 32137 27968
rect 32171 27965 32183 27999
rect 33870 27996 33876 28008
rect 33534 27968 33876 27996
rect 32125 27959 32183 27965
rect 33870 27956 33876 27968
rect 33928 27956 33934 28008
rect 27522 27928 27528 27940
rect 26375 27900 26556 27928
rect 27356 27900 27528 27928
rect 26375 27897 26387 27900
rect 26329 27891 26387 27897
rect 25685 27863 25743 27869
rect 25685 27860 25697 27863
rect 25188 27832 25697 27860
rect 25188 27820 25194 27832
rect 25685 27829 25697 27832
rect 25731 27829 25743 27863
rect 26528 27860 26556 27900
rect 27522 27888 27528 27900
rect 27580 27888 27586 27940
rect 27614 27888 27620 27940
rect 27672 27888 27678 27940
rect 31573 27931 31631 27937
rect 31573 27928 31585 27931
rect 29380 27900 31585 27928
rect 29380 27872 29408 27900
rect 31573 27897 31585 27900
rect 31619 27897 31631 27931
rect 31573 27891 31631 27897
rect 31665 27931 31723 27937
rect 31665 27897 31677 27931
rect 31711 27928 31723 27931
rect 32306 27928 32312 27940
rect 31711 27900 32312 27928
rect 31711 27897 31723 27900
rect 31665 27891 31723 27897
rect 32306 27888 32312 27900
rect 32364 27888 32370 27940
rect 32674 27888 32680 27940
rect 32732 27888 32738 27940
rect 29362 27860 29368 27872
rect 26528 27832 29368 27860
rect 25685 27823 25743 27829
rect 29362 27820 29368 27832
rect 29420 27820 29426 27872
rect 30650 27820 30656 27872
rect 30708 27860 30714 27872
rect 30745 27863 30803 27869
rect 30745 27860 30757 27863
rect 30708 27832 30757 27860
rect 30708 27820 30714 27832
rect 30745 27829 30757 27832
rect 30791 27829 30803 27863
rect 32692 27860 32720 27888
rect 33873 27863 33931 27869
rect 33873 27860 33885 27863
rect 32692 27832 33885 27860
rect 30745 27823 30803 27829
rect 33873 27829 33885 27832
rect 33919 27829 33931 27863
rect 33873 27823 33931 27829
rect 2760 27770 34316 27792
rect 2760 27718 7210 27770
rect 7262 27718 7274 27770
rect 7326 27718 7338 27770
rect 7390 27718 7402 27770
rect 7454 27718 7466 27770
rect 7518 27718 15099 27770
rect 15151 27718 15163 27770
rect 15215 27718 15227 27770
rect 15279 27718 15291 27770
rect 15343 27718 15355 27770
rect 15407 27718 22988 27770
rect 23040 27718 23052 27770
rect 23104 27718 23116 27770
rect 23168 27718 23180 27770
rect 23232 27718 23244 27770
rect 23296 27718 30877 27770
rect 30929 27718 30941 27770
rect 30993 27718 31005 27770
rect 31057 27718 31069 27770
rect 31121 27718 31133 27770
rect 31185 27718 34316 27770
rect 2760 27696 34316 27718
rect 6730 27616 6736 27668
rect 6788 27616 6794 27668
rect 8202 27616 8208 27668
rect 8260 27616 8266 27668
rect 8386 27616 8392 27668
rect 8444 27616 8450 27668
rect 11057 27659 11115 27665
rect 11057 27625 11069 27659
rect 11103 27656 11115 27659
rect 11146 27656 11152 27668
rect 11103 27628 11152 27656
rect 11103 27625 11115 27628
rect 11057 27619 11115 27625
rect 11146 27616 11152 27628
rect 11204 27616 11210 27668
rect 11238 27616 11244 27668
rect 11296 27656 11302 27668
rect 11517 27659 11575 27665
rect 11517 27656 11529 27659
rect 11296 27628 11529 27656
rect 11296 27616 11302 27628
rect 11517 27625 11529 27628
rect 11563 27625 11575 27659
rect 11517 27619 11575 27625
rect 11606 27616 11612 27668
rect 11664 27616 11670 27668
rect 12618 27616 12624 27668
rect 12676 27656 12682 27668
rect 12676 27628 14320 27656
rect 12676 27616 12682 27628
rect 4522 27548 4528 27600
rect 4580 27548 4586 27600
rect 4816 27560 5580 27588
rect 4816 27529 4844 27560
rect 5552 27532 5580 27560
rect 7006 27548 7012 27600
rect 7064 27548 7070 27600
rect 4801 27523 4859 27529
rect 3436 27452 3464 27506
rect 4801 27489 4813 27523
rect 4847 27489 4859 27523
rect 4801 27483 4859 27489
rect 5074 27480 5080 27532
rect 5132 27480 5138 27532
rect 5534 27480 5540 27532
rect 5592 27480 5598 27532
rect 6917 27523 6975 27529
rect 6917 27489 6929 27523
rect 6963 27489 6975 27523
rect 6917 27483 6975 27489
rect 4985 27455 5043 27461
rect 4985 27452 4997 27455
rect 3436 27424 4997 27452
rect 4985 27421 4997 27424
rect 5031 27421 5043 27455
rect 4985 27415 5043 27421
rect 5258 27412 5264 27464
rect 5316 27412 5322 27464
rect 5350 27412 5356 27464
rect 5408 27452 5414 27464
rect 5997 27455 6055 27461
rect 5997 27452 6009 27455
rect 5408 27424 6009 27452
rect 5408 27412 5414 27424
rect 5997 27421 6009 27424
rect 6043 27421 6055 27455
rect 6932 27452 6960 27483
rect 7098 27480 7104 27532
rect 7156 27480 7162 27532
rect 7285 27523 7343 27529
rect 7285 27489 7297 27523
rect 7331 27520 7343 27523
rect 7558 27520 7564 27532
rect 7331 27492 7564 27520
rect 7331 27489 7343 27492
rect 7285 27483 7343 27489
rect 7558 27480 7564 27492
rect 7616 27480 7622 27532
rect 8220 27520 8248 27616
rect 10962 27548 10968 27600
rect 11020 27588 11026 27600
rect 11425 27591 11483 27597
rect 11020 27560 11342 27588
rect 11020 27548 11026 27560
rect 8297 27523 8355 27529
rect 8297 27520 8309 27523
rect 8220 27492 8309 27520
rect 8297 27489 8309 27492
rect 8343 27520 8355 27523
rect 9493 27523 9551 27529
rect 9493 27520 9505 27523
rect 8343 27492 9505 27520
rect 8343 27489 8355 27492
rect 8297 27483 8355 27489
rect 9493 27489 9505 27492
rect 9539 27489 9551 27523
rect 9493 27483 9551 27489
rect 9950 27480 9956 27532
rect 10008 27520 10014 27532
rect 10778 27520 10784 27532
rect 10008 27492 10784 27520
rect 10008 27480 10014 27492
rect 10778 27480 10784 27492
rect 10836 27520 10842 27532
rect 11314 27529 11342 27560
rect 11425 27557 11437 27591
rect 11471 27588 11483 27591
rect 11624 27588 11652 27616
rect 11471 27560 11652 27588
rect 11471 27557 11483 27560
rect 11425 27551 11483 27557
rect 11974 27548 11980 27600
rect 12032 27588 12038 27600
rect 12437 27591 12495 27597
rect 12437 27588 12449 27591
rect 12032 27560 12449 27588
rect 12032 27548 12038 27560
rect 12437 27557 12449 27560
rect 12483 27557 12495 27591
rect 12437 27551 12495 27557
rect 13906 27548 13912 27600
rect 13964 27588 13970 27600
rect 14001 27591 14059 27597
rect 14001 27588 14013 27591
rect 13964 27560 14013 27588
rect 13964 27548 13970 27560
rect 14001 27557 14013 27560
rect 14047 27557 14059 27591
rect 14001 27551 14059 27557
rect 14090 27548 14096 27600
rect 14148 27588 14154 27600
rect 14201 27591 14259 27597
rect 14201 27588 14213 27591
rect 14148 27560 14213 27588
rect 14148 27548 14154 27560
rect 14201 27557 14213 27560
rect 14247 27557 14259 27591
rect 14292 27588 14320 27628
rect 14366 27616 14372 27668
rect 14424 27616 14430 27668
rect 14476 27628 15240 27656
rect 14476 27588 14504 27628
rect 14292 27560 14504 27588
rect 14201 27551 14259 27557
rect 10873 27523 10931 27529
rect 10873 27520 10885 27523
rect 10836 27492 10885 27520
rect 10836 27480 10842 27492
rect 10873 27489 10885 27492
rect 10919 27520 10931 27523
rect 11314 27523 11391 27529
rect 10919 27492 11100 27520
rect 10919 27489 10931 27492
rect 10873 27483 10931 27489
rect 11072 27486 11100 27492
rect 11314 27490 11345 27523
rect 11333 27489 11345 27490
rect 11379 27489 11391 27523
rect 11790 27520 11796 27532
rect 11751 27492 11796 27520
rect 10689 27455 10747 27461
rect 6932 27424 7696 27452
rect 5997 27415 6055 27421
rect 3053 27319 3111 27325
rect 3053 27285 3065 27319
rect 3099 27316 3111 27319
rect 4430 27316 4436 27328
rect 3099 27288 4436 27316
rect 3099 27285 3111 27288
rect 3053 27279 3111 27285
rect 4430 27276 4436 27288
rect 4488 27276 4494 27328
rect 5810 27276 5816 27328
rect 5868 27276 5874 27328
rect 5994 27276 6000 27328
rect 6052 27316 6058 27328
rect 7668 27325 7696 27424
rect 10689 27421 10701 27455
rect 10735 27452 10747 27455
rect 10962 27452 10968 27464
rect 10735 27424 10968 27452
rect 10735 27421 10747 27424
rect 10689 27415 10747 27421
rect 10962 27412 10968 27424
rect 11020 27412 11026 27464
rect 11072 27458 11284 27486
rect 11333 27483 11391 27489
rect 11790 27480 11796 27492
rect 11848 27518 11854 27532
rect 12069 27523 12127 27529
rect 12069 27520 12081 27523
rect 11900 27518 12081 27520
rect 11848 27492 12081 27518
rect 11848 27490 11928 27492
rect 11848 27480 11854 27490
rect 12069 27489 12081 27492
rect 12115 27489 12127 27523
rect 12069 27483 12127 27489
rect 12158 27480 12164 27532
rect 12216 27520 12222 27532
rect 12529 27523 12587 27529
rect 12529 27520 12541 27523
rect 12216 27492 12541 27520
rect 12216 27480 12222 27492
rect 12529 27489 12541 27492
rect 12575 27520 12587 27523
rect 13449 27523 13507 27529
rect 13449 27520 13461 27523
rect 12575 27492 13461 27520
rect 12575 27489 12587 27492
rect 12529 27483 12587 27489
rect 13449 27489 13461 27492
rect 13495 27489 13507 27523
rect 13449 27483 13507 27489
rect 13633 27523 13691 27529
rect 13633 27489 13645 27523
rect 13679 27520 13691 27523
rect 14366 27520 14372 27532
rect 13679 27492 14372 27520
rect 13679 27489 13691 27492
rect 13633 27483 13691 27489
rect 14366 27480 14372 27492
rect 14424 27480 14430 27532
rect 15212 27529 15240 27628
rect 15470 27616 15476 27668
rect 15528 27616 15534 27668
rect 15562 27616 15568 27668
rect 15620 27616 15626 27668
rect 16022 27616 16028 27668
rect 16080 27656 16086 27668
rect 16209 27659 16267 27665
rect 16209 27656 16221 27659
rect 16080 27628 16221 27656
rect 16080 27616 16086 27628
rect 16209 27625 16221 27628
rect 16255 27625 16267 27659
rect 16209 27619 16267 27625
rect 16574 27616 16580 27668
rect 16632 27616 16638 27668
rect 16758 27616 16764 27668
rect 16816 27616 16822 27668
rect 17034 27616 17040 27668
rect 17092 27656 17098 27668
rect 17770 27656 17776 27668
rect 17092 27628 17776 27656
rect 17092 27616 17098 27628
rect 17770 27616 17776 27628
rect 17828 27616 17834 27668
rect 18046 27616 18052 27668
rect 18104 27616 18110 27668
rect 18141 27659 18199 27665
rect 18141 27625 18153 27659
rect 18187 27625 18199 27659
rect 18141 27619 18199 27625
rect 15381 27591 15439 27597
rect 15381 27557 15393 27591
rect 15427 27588 15439 27591
rect 15488 27588 15516 27616
rect 15427 27560 15516 27588
rect 15427 27557 15439 27560
rect 15381 27551 15439 27557
rect 15197 27523 15255 27529
rect 15197 27489 15209 27523
rect 15243 27489 15255 27523
rect 15580 27520 15608 27616
rect 16117 27523 16175 27529
rect 16117 27520 16129 27523
rect 15580 27492 16129 27520
rect 15197 27483 15255 27489
rect 16117 27489 16129 27492
rect 16163 27489 16175 27523
rect 16592 27520 16620 27616
rect 17218 27548 17224 27600
rect 17276 27548 17282 27600
rect 17681 27591 17739 27597
rect 17681 27557 17693 27591
rect 17727 27588 17739 27591
rect 18064 27588 18092 27616
rect 17727 27560 18092 27588
rect 18156 27588 18184 27619
rect 20070 27616 20076 27668
rect 20128 27616 20134 27668
rect 28166 27656 28172 27668
rect 27540 27628 28172 27656
rect 18601 27591 18659 27597
rect 18601 27588 18613 27591
rect 18156 27560 18613 27588
rect 17727 27557 17739 27560
rect 17681 27551 17739 27557
rect 18601 27557 18613 27560
rect 18647 27557 18659 27591
rect 18601 27551 18659 27557
rect 19058 27548 19064 27600
rect 19116 27548 19122 27600
rect 20990 27548 20996 27600
rect 21048 27548 21054 27600
rect 21818 27548 21824 27600
rect 21876 27588 21882 27600
rect 22925 27591 22983 27597
rect 22925 27588 22937 27591
rect 21876 27560 22937 27588
rect 21876 27548 21882 27560
rect 22925 27557 22937 27560
rect 22971 27557 22983 27591
rect 22925 27551 22983 27557
rect 16669 27523 16727 27529
rect 16669 27520 16681 27523
rect 16592 27492 16681 27520
rect 16117 27483 16175 27489
rect 16669 27489 16681 27492
rect 16715 27489 16727 27523
rect 16669 27483 16727 27489
rect 11256 27452 11284 27458
rect 12253 27455 12311 27461
rect 12253 27452 12265 27455
rect 11256 27424 12265 27452
rect 12253 27421 12265 27424
rect 12299 27421 12311 27455
rect 12253 27415 12311 27421
rect 13541 27455 13599 27461
rect 13541 27421 13553 27455
rect 13587 27452 13599 27455
rect 14642 27452 14648 27464
rect 13587 27424 14648 27452
rect 13587 27421 13599 27424
rect 13541 27415 13599 27421
rect 12268 27384 12296 27415
rect 14642 27412 14648 27424
rect 14700 27412 14706 27464
rect 15212 27452 15240 27483
rect 15838 27452 15844 27464
rect 15212 27424 15844 27452
rect 15838 27412 15844 27424
rect 15896 27452 15902 27464
rect 15933 27455 15991 27461
rect 15933 27452 15945 27455
rect 15896 27424 15945 27452
rect 15896 27412 15902 27424
rect 15933 27421 15945 27424
rect 15979 27421 15991 27455
rect 15933 27415 15991 27421
rect 17218 27412 17224 27464
rect 17276 27452 17282 27464
rect 17497 27455 17555 27461
rect 17497 27452 17509 27455
rect 17276 27424 17509 27452
rect 17276 27412 17282 27424
rect 17497 27421 17509 27424
rect 17543 27421 17555 27455
rect 17497 27415 17555 27421
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 14918 27384 14924 27396
rect 11072 27356 12204 27384
rect 12268 27356 14924 27384
rect 11072 27328 11100 27356
rect 6641 27319 6699 27325
rect 6641 27316 6653 27319
rect 6052 27288 6653 27316
rect 6052 27276 6058 27288
rect 6641 27285 6653 27288
rect 6687 27285 6699 27319
rect 6641 27279 6699 27285
rect 7653 27319 7711 27325
rect 7653 27285 7665 27319
rect 7699 27316 7711 27319
rect 7742 27316 7748 27328
rect 7699 27288 7748 27316
rect 7699 27285 7711 27288
rect 7653 27279 7711 27285
rect 7742 27276 7748 27288
rect 7800 27276 7806 27328
rect 9582 27276 9588 27328
rect 9640 27276 9646 27328
rect 11054 27276 11060 27328
rect 11112 27276 11118 27328
rect 11514 27276 11520 27328
rect 11572 27316 11578 27328
rect 11885 27319 11943 27325
rect 11885 27316 11897 27319
rect 11572 27288 11897 27316
rect 11572 27276 11578 27288
rect 11885 27285 11897 27288
rect 11931 27285 11943 27319
rect 12176 27316 12204 27356
rect 13814 27316 13820 27328
rect 12176 27288 13820 27316
rect 11885 27279 11943 27285
rect 13814 27276 13820 27288
rect 13872 27276 13878 27328
rect 14200 27325 14228 27356
rect 14918 27344 14924 27356
rect 14976 27344 14982 27396
rect 14185 27319 14243 27325
rect 14185 27285 14197 27319
rect 14231 27285 14243 27319
rect 14185 27279 14243 27285
rect 14274 27276 14280 27328
rect 14332 27316 14338 27328
rect 14645 27319 14703 27325
rect 14645 27316 14657 27319
rect 14332 27288 14657 27316
rect 14332 27276 14338 27288
rect 14645 27285 14657 27288
rect 14691 27316 14703 27319
rect 15470 27316 15476 27328
rect 14691 27288 15476 27316
rect 14691 27285 14703 27288
rect 14645 27279 14703 27285
rect 15470 27276 15476 27288
rect 15528 27276 15534 27328
rect 18340 27316 18368 27415
rect 19242 27412 19248 27464
rect 19300 27452 19306 27464
rect 21082 27452 21088 27464
rect 19300 27424 21088 27452
rect 19300 27412 19306 27424
rect 21082 27412 21088 27424
rect 21140 27412 21146 27464
rect 21726 27412 21732 27464
rect 21784 27412 21790 27464
rect 22005 27455 22063 27461
rect 22005 27421 22017 27455
rect 22051 27421 22063 27455
rect 22940 27452 22968 27551
rect 23382 27548 23388 27600
rect 23440 27548 23446 27600
rect 23750 27548 23756 27600
rect 23808 27548 23814 27600
rect 23845 27591 23903 27597
rect 23845 27557 23857 27591
rect 23891 27588 23903 27591
rect 24670 27588 24676 27600
rect 23891 27560 24676 27588
rect 23891 27557 23903 27560
rect 23845 27551 23903 27557
rect 24670 27548 24676 27560
rect 24728 27588 24734 27600
rect 25041 27591 25099 27597
rect 25041 27588 25053 27591
rect 24728 27560 25053 27588
rect 24728 27548 24734 27560
rect 25041 27557 25053 27560
rect 25087 27557 25099 27591
rect 25041 27551 25099 27557
rect 26142 27548 26148 27600
rect 26200 27588 26206 27600
rect 27540 27588 27568 27628
rect 28166 27616 28172 27628
rect 28224 27616 28230 27668
rect 28718 27616 28724 27668
rect 28776 27616 28782 27668
rect 29104 27628 30236 27656
rect 26200 27560 27568 27588
rect 26200 27548 26206 27560
rect 23109 27523 23167 27529
rect 23109 27489 23121 27523
rect 23155 27520 23167 27523
rect 23400 27520 23428 27548
rect 23155 27492 23428 27520
rect 23155 27489 23167 27492
rect 23109 27483 23167 27489
rect 24210 27480 24216 27532
rect 24268 27480 24274 27532
rect 27540 27529 27568 27560
rect 27617 27591 27675 27597
rect 27617 27557 27629 27591
rect 27663 27588 27675 27591
rect 28350 27588 28356 27600
rect 27663 27560 28356 27588
rect 27663 27557 27675 27560
rect 27617 27551 27675 27557
rect 28350 27548 28356 27560
rect 28408 27548 28414 27600
rect 29104 27588 29132 27628
rect 28828 27560 29132 27588
rect 29181 27591 29239 27597
rect 24949 27523 25007 27529
rect 24949 27489 24961 27523
rect 24995 27520 25007 27523
rect 26513 27523 26571 27529
rect 26513 27520 26525 27523
rect 24995 27492 26525 27520
rect 24995 27489 25007 27492
rect 24949 27483 25007 27489
rect 26513 27489 26525 27492
rect 26559 27489 26571 27523
rect 26513 27483 26571 27489
rect 27525 27523 27583 27529
rect 27525 27489 27537 27523
rect 27571 27489 27583 27523
rect 27525 27483 27583 27489
rect 27706 27480 27712 27532
rect 27764 27480 27770 27532
rect 27893 27523 27951 27529
rect 27893 27489 27905 27523
rect 27939 27489 27951 27523
rect 27893 27483 27951 27489
rect 23569 27455 23627 27461
rect 23569 27452 23581 27455
rect 22940 27424 23581 27452
rect 22005 27415 22063 27421
rect 23569 27421 23581 27424
rect 23615 27421 23627 27455
rect 23569 27415 23627 27421
rect 19996 27356 20760 27384
rect 18966 27316 18972 27328
rect 18340 27288 18972 27316
rect 18966 27276 18972 27288
rect 19024 27316 19030 27328
rect 19996 27316 20024 27356
rect 19024 27288 20024 27316
rect 19024 27276 19030 27288
rect 20254 27276 20260 27328
rect 20312 27276 20318 27328
rect 20732 27316 20760 27356
rect 22020 27328 22048 27415
rect 24228 27393 24256 27480
rect 24302 27412 24308 27464
rect 24360 27412 24366 27464
rect 24854 27412 24860 27464
rect 24912 27452 24918 27464
rect 25593 27455 25651 27461
rect 25593 27452 25605 27455
rect 24912 27424 25605 27452
rect 24912 27412 24918 27424
rect 25593 27421 25605 27424
rect 25639 27421 25651 27455
rect 25593 27415 25651 27421
rect 26326 27412 26332 27464
rect 26384 27412 26390 27464
rect 27154 27412 27160 27464
rect 27212 27452 27218 27464
rect 27908 27452 27936 27483
rect 28626 27480 28632 27532
rect 28684 27520 28690 27532
rect 28828 27529 28856 27560
rect 29181 27557 29193 27591
rect 29227 27588 29239 27591
rect 30098 27588 30104 27600
rect 29227 27560 30104 27588
rect 29227 27557 29239 27560
rect 29181 27551 29239 27557
rect 30098 27548 30104 27560
rect 30156 27548 30162 27600
rect 30208 27588 30236 27628
rect 30558 27616 30564 27668
rect 30616 27616 30622 27668
rect 31662 27616 31668 27668
rect 31720 27656 31726 27668
rect 32030 27656 32036 27668
rect 31720 27628 32036 27656
rect 31720 27616 31726 27628
rect 32030 27616 32036 27628
rect 32088 27656 32094 27668
rect 32490 27656 32496 27668
rect 32088 27628 32496 27656
rect 32088 27616 32094 27628
rect 32490 27616 32496 27628
rect 32548 27616 32554 27668
rect 32674 27616 32680 27668
rect 32732 27656 32738 27668
rect 33137 27659 33195 27665
rect 33137 27656 33149 27659
rect 32732 27628 33149 27656
rect 32732 27616 32738 27628
rect 33137 27625 33149 27628
rect 33183 27625 33195 27659
rect 33137 27619 33195 27625
rect 30576 27588 30604 27616
rect 31297 27591 31355 27597
rect 31297 27588 31309 27591
rect 30208 27560 30512 27588
rect 30576 27560 31309 27588
rect 28813 27523 28871 27529
rect 28813 27520 28825 27523
rect 28684 27492 28825 27520
rect 28684 27480 28690 27492
rect 28813 27489 28825 27492
rect 28859 27489 28871 27523
rect 28813 27483 28871 27489
rect 28902 27480 28908 27532
rect 28960 27480 28966 27532
rect 29089 27523 29147 27529
rect 29089 27489 29101 27523
rect 29135 27489 29147 27523
rect 29089 27483 29147 27489
rect 29104 27452 29132 27483
rect 29270 27480 29276 27532
rect 29328 27480 29334 27532
rect 30374 27520 30380 27532
rect 29472 27492 30380 27520
rect 27212 27424 29132 27452
rect 27212 27412 27218 27424
rect 24213 27387 24271 27393
rect 24213 27353 24225 27387
rect 24259 27353 24271 27387
rect 27341 27387 27399 27393
rect 24213 27347 24271 27353
rect 26712 27356 27292 27384
rect 26712 27328 26740 27356
rect 21266 27316 21272 27328
rect 20732 27288 21272 27316
rect 21266 27276 21272 27288
rect 21324 27316 21330 27328
rect 22002 27316 22008 27328
rect 21324 27288 22008 27316
rect 21324 27276 21330 27288
rect 22002 27276 22008 27288
rect 22060 27276 22066 27328
rect 23201 27319 23259 27325
rect 23201 27285 23213 27319
rect 23247 27316 23259 27319
rect 23290 27316 23296 27328
rect 23247 27288 23296 27316
rect 23247 27285 23259 27288
rect 23201 27279 23259 27285
rect 23290 27276 23296 27288
rect 23348 27276 23354 27328
rect 24118 27276 24124 27328
rect 24176 27316 24182 27328
rect 25777 27319 25835 27325
rect 25777 27316 25789 27319
rect 24176 27288 25789 27316
rect 24176 27276 24182 27288
rect 25777 27285 25789 27288
rect 25823 27285 25835 27319
rect 25777 27279 25835 27285
rect 26694 27276 26700 27328
rect 26752 27276 26758 27328
rect 27062 27276 27068 27328
rect 27120 27276 27126 27328
rect 27264 27316 27292 27356
rect 27341 27353 27353 27387
rect 27387 27384 27399 27387
rect 27614 27384 27620 27396
rect 27387 27356 27620 27384
rect 27387 27353 27399 27356
rect 27341 27347 27399 27353
rect 27614 27344 27620 27356
rect 27672 27344 27678 27396
rect 29472 27393 29500 27492
rect 30374 27480 30380 27492
rect 30432 27480 30438 27532
rect 30484 27520 30512 27560
rect 31297 27557 31309 27560
rect 31343 27557 31355 27591
rect 31297 27551 31355 27557
rect 31386 27548 31392 27600
rect 31444 27588 31450 27600
rect 33045 27591 33103 27597
rect 33045 27588 33057 27591
rect 31444 27560 33057 27588
rect 31444 27548 31450 27560
rect 33045 27557 33057 27560
rect 33091 27557 33103 27591
rect 33045 27551 33103 27557
rect 31205 27523 31263 27529
rect 31205 27520 31217 27523
rect 30484 27492 31217 27520
rect 31205 27489 31217 27492
rect 31251 27489 31263 27523
rect 31205 27483 31263 27489
rect 31849 27523 31907 27529
rect 31849 27489 31861 27523
rect 31895 27489 31907 27523
rect 33965 27523 34023 27529
rect 31849 27483 31907 27489
rect 32140 27492 33272 27520
rect 29546 27412 29552 27464
rect 29604 27412 29610 27464
rect 30098 27412 30104 27464
rect 30156 27412 30162 27464
rect 30558 27412 30564 27464
rect 30616 27412 30622 27464
rect 29457 27387 29515 27393
rect 27724 27356 29408 27384
rect 27724 27316 27752 27356
rect 27264 27288 27752 27316
rect 28166 27276 28172 27328
rect 28224 27316 28230 27328
rect 29270 27316 29276 27328
rect 28224 27288 29276 27316
rect 28224 27276 28230 27288
rect 29270 27276 29276 27288
rect 29328 27276 29334 27328
rect 29380 27316 29408 27356
rect 29457 27353 29469 27387
rect 29503 27353 29515 27387
rect 31864 27384 31892 27483
rect 32140 27464 32168 27492
rect 33060 27464 33088 27492
rect 31941 27455 31999 27461
rect 31941 27421 31953 27455
rect 31987 27421 31999 27455
rect 31941 27415 31999 27421
rect 29457 27347 29515 27353
rect 30116 27356 31892 27384
rect 31956 27384 31984 27415
rect 32030 27412 32036 27464
rect 32088 27412 32094 27464
rect 32122 27412 32128 27464
rect 32180 27412 32186 27464
rect 32398 27412 32404 27464
rect 32456 27412 32462 27464
rect 33042 27412 33048 27464
rect 33100 27412 33106 27464
rect 33244 27461 33272 27492
rect 33965 27489 33977 27523
rect 34011 27520 34023 27523
rect 34011 27492 35204 27520
rect 34011 27489 34023 27492
rect 33965 27483 34023 27489
rect 33229 27455 33287 27461
rect 33229 27421 33241 27455
rect 33275 27421 33287 27455
rect 33229 27415 33287 27421
rect 33410 27412 33416 27464
rect 33468 27412 33474 27464
rect 32416 27384 32444 27412
rect 32582 27384 32588 27396
rect 31956 27356 32588 27384
rect 30116 27316 30144 27356
rect 32582 27344 32588 27356
rect 32640 27344 32646 27396
rect 32677 27387 32735 27393
rect 32677 27353 32689 27387
rect 32723 27384 32735 27387
rect 33428 27384 33456 27412
rect 35176 27396 35204 27492
rect 32723 27356 33456 27384
rect 32723 27353 32735 27356
rect 32677 27347 32735 27353
rect 35158 27344 35164 27396
rect 35216 27344 35222 27396
rect 29380 27288 30144 27316
rect 30742 27276 30748 27328
rect 30800 27316 30806 27328
rect 31113 27319 31171 27325
rect 31113 27316 31125 27319
rect 30800 27288 31125 27316
rect 30800 27276 30806 27288
rect 31113 27285 31125 27288
rect 31159 27316 31171 27319
rect 31386 27316 31392 27328
rect 31159 27288 31392 27316
rect 31159 27285 31171 27288
rect 31113 27279 31171 27285
rect 31386 27276 31392 27288
rect 31444 27276 31450 27328
rect 31481 27319 31539 27325
rect 31481 27285 31493 27319
rect 31527 27316 31539 27319
rect 32030 27316 32036 27328
rect 31527 27288 32036 27316
rect 31527 27285 31539 27288
rect 31481 27279 31539 27285
rect 32030 27276 32036 27288
rect 32088 27276 32094 27328
rect 33778 27276 33784 27328
rect 33836 27276 33842 27328
rect 2760 27226 34316 27248
rect 2760 27174 6550 27226
rect 6602 27174 6614 27226
rect 6666 27174 6678 27226
rect 6730 27174 6742 27226
rect 6794 27174 6806 27226
rect 6858 27174 14439 27226
rect 14491 27174 14503 27226
rect 14555 27174 14567 27226
rect 14619 27174 14631 27226
rect 14683 27174 14695 27226
rect 14747 27174 22328 27226
rect 22380 27174 22392 27226
rect 22444 27174 22456 27226
rect 22508 27174 22520 27226
rect 22572 27174 22584 27226
rect 22636 27174 30217 27226
rect 30269 27174 30281 27226
rect 30333 27174 30345 27226
rect 30397 27174 30409 27226
rect 30461 27174 30473 27226
rect 30525 27174 34316 27226
rect 2760 27152 34316 27174
rect 3970 27072 3976 27124
rect 4028 27072 4034 27124
rect 5258 27072 5264 27124
rect 5316 27112 5322 27124
rect 5445 27115 5503 27121
rect 5445 27112 5457 27115
rect 5316 27084 5457 27112
rect 5316 27072 5322 27084
rect 5445 27081 5457 27084
rect 5491 27081 5503 27115
rect 5445 27075 5503 27081
rect 6086 27072 6092 27124
rect 6144 27112 6150 27124
rect 6362 27112 6368 27124
rect 6144 27084 6368 27112
rect 6144 27072 6150 27084
rect 6362 27072 6368 27084
rect 6420 27112 6426 27124
rect 6917 27115 6975 27121
rect 6917 27112 6929 27115
rect 6420 27084 6929 27112
rect 6420 27072 6426 27084
rect 6917 27081 6929 27084
rect 6963 27081 6975 27115
rect 6917 27075 6975 27081
rect 7834 27072 7840 27124
rect 7892 27072 7898 27124
rect 8202 27072 8208 27124
rect 8260 27072 8266 27124
rect 10042 27072 10048 27124
rect 10100 27072 10106 27124
rect 10321 27115 10379 27121
rect 10321 27081 10333 27115
rect 10367 27112 10379 27115
rect 11422 27112 11428 27124
rect 10367 27084 11428 27112
rect 10367 27081 10379 27084
rect 10321 27075 10379 27081
rect 11422 27072 11428 27084
rect 11480 27072 11486 27124
rect 12618 27112 12624 27124
rect 12406 27084 12624 27112
rect 5626 27044 5632 27056
rect 4540 27016 5632 27044
rect 4430 26936 4436 26988
rect 4488 26936 4494 26988
rect 4540 26985 4568 27016
rect 5626 27004 5632 27016
rect 5684 27044 5690 27056
rect 5684 27016 6040 27044
rect 5684 27004 5690 27016
rect 4525 26979 4583 26985
rect 4525 26945 4537 26979
rect 4571 26945 4583 26979
rect 4525 26939 4583 26945
rect 1302 26868 1308 26920
rect 1360 26908 1366 26920
rect 3053 26911 3111 26917
rect 3053 26908 3065 26911
rect 1360 26880 3065 26908
rect 1360 26868 1366 26880
rect 3053 26877 3065 26880
rect 3099 26877 3111 26911
rect 3053 26871 3111 26877
rect 3881 26911 3939 26917
rect 3881 26877 3893 26911
rect 3927 26908 3939 26911
rect 4540 26908 4568 26939
rect 4614 26936 4620 26988
rect 4672 26976 4678 26988
rect 6012 26985 6040 27016
rect 5905 26979 5963 26985
rect 5905 26976 5917 26979
rect 4672 26948 5917 26976
rect 4672 26936 4678 26948
rect 5905 26945 5917 26948
rect 5951 26945 5963 26979
rect 5905 26939 5963 26945
rect 5997 26979 6055 26985
rect 5997 26945 6009 26979
rect 6043 26945 6055 26979
rect 8220 26976 8248 27072
rect 5997 26939 6055 26945
rect 7208 26948 8248 26976
rect 10060 26976 10088 27072
rect 11149 27047 11207 27053
rect 11149 27013 11161 27047
rect 11195 27044 11207 27047
rect 11330 27044 11336 27056
rect 11195 27016 11336 27044
rect 11195 27013 11207 27016
rect 11149 27007 11207 27013
rect 11330 27004 11336 27016
rect 11388 27004 11394 27056
rect 11514 27044 11520 27056
rect 11440 27016 11520 27044
rect 10060 26948 11008 26976
rect 4890 26908 4896 26920
rect 3927 26880 4896 26908
rect 3927 26877 3939 26880
rect 3881 26871 3939 26877
rect 4890 26868 4896 26880
rect 4948 26868 4954 26920
rect 5813 26911 5871 26917
rect 5813 26877 5825 26911
rect 5859 26908 5871 26911
rect 6178 26908 6184 26920
rect 5859 26880 6184 26908
rect 5859 26877 5871 26880
rect 5813 26871 5871 26877
rect 6178 26868 6184 26880
rect 6236 26868 6242 26920
rect 6270 26868 6276 26920
rect 6328 26868 6334 26920
rect 7208 26917 7236 26948
rect 7193 26911 7251 26917
rect 7193 26877 7205 26911
rect 7239 26877 7251 26911
rect 7193 26871 7251 26877
rect 8018 26868 8024 26920
rect 8076 26908 8082 26920
rect 8573 26911 8631 26917
rect 8573 26908 8585 26911
rect 8076 26880 8585 26908
rect 8076 26868 8082 26880
rect 8573 26877 8585 26880
rect 8619 26877 8631 26911
rect 8573 26871 8631 26877
rect 10594 26868 10600 26920
rect 10652 26908 10658 26920
rect 10722 26911 10780 26917
rect 10722 26908 10734 26911
rect 10652 26880 10734 26908
rect 10652 26868 10658 26880
rect 10722 26877 10734 26880
rect 10768 26877 10780 26911
rect 10980 26908 11008 26948
rect 11054 26936 11060 26988
rect 11112 26976 11118 26988
rect 11241 26979 11299 26985
rect 11241 26976 11253 26979
rect 11112 26948 11253 26976
rect 11112 26936 11118 26948
rect 11241 26945 11253 26948
rect 11287 26945 11299 26979
rect 11241 26939 11299 26945
rect 11440 26917 11468 27016
rect 11514 27004 11520 27016
rect 11572 27004 11578 27056
rect 12406 27044 12434 27084
rect 12618 27072 12624 27084
rect 12676 27072 12682 27124
rect 13817 27115 13875 27121
rect 13817 27081 13829 27115
rect 13863 27081 13875 27115
rect 13817 27075 13875 27081
rect 14001 27115 14059 27121
rect 14001 27081 14013 27115
rect 14047 27112 14059 27115
rect 14090 27112 14096 27124
rect 14047 27084 14096 27112
rect 14047 27081 14059 27084
rect 14001 27075 14059 27081
rect 11624 27016 12434 27044
rect 13832 27044 13860 27075
rect 14090 27072 14096 27084
rect 14148 27072 14154 27124
rect 14826 27072 14832 27124
rect 14884 27112 14890 27124
rect 14884 27084 15148 27112
rect 14884 27072 14890 27084
rect 14274 27044 14280 27056
rect 13832 27016 14280 27044
rect 11425 26911 11483 26917
rect 11425 26908 11437 26911
rect 10980 26880 11437 26908
rect 10722 26871 10780 26877
rect 11425 26877 11437 26880
rect 11471 26877 11483 26911
rect 11425 26871 11483 26877
rect 11517 26911 11575 26917
rect 11517 26877 11529 26911
rect 11563 26908 11575 26911
rect 11624 26908 11652 27016
rect 14274 27004 14280 27016
rect 14332 27004 14338 27056
rect 11790 26936 11796 26988
rect 11848 26976 11854 26988
rect 13078 26976 13084 26988
rect 11848 26948 13084 26976
rect 11848 26936 11854 26948
rect 13078 26936 13084 26948
rect 13136 26976 13142 26988
rect 13265 26979 13323 26985
rect 13265 26976 13277 26979
rect 13136 26948 13277 26976
rect 13136 26936 13142 26948
rect 13265 26945 13277 26948
rect 13311 26945 13323 26979
rect 13265 26939 13323 26945
rect 13814 26936 13820 26988
rect 13872 26936 13878 26988
rect 11563 26880 11652 26908
rect 11701 26911 11759 26917
rect 11563 26877 11575 26880
rect 11517 26871 11575 26877
rect 11701 26877 11713 26911
rect 11747 26877 11759 26911
rect 11701 26871 11759 26877
rect 4341 26843 4399 26849
rect 4341 26809 4353 26843
rect 4387 26840 4399 26843
rect 5534 26840 5540 26852
rect 4387 26812 5540 26840
rect 4387 26809 4399 26812
rect 4341 26803 4399 26809
rect 5534 26800 5540 26812
rect 5592 26800 5598 26852
rect 5718 26800 5724 26852
rect 5776 26840 5782 26852
rect 5776 26812 7144 26840
rect 5776 26800 5782 26812
rect 3237 26775 3295 26781
rect 3237 26741 3249 26775
rect 3283 26772 3295 26775
rect 3602 26772 3608 26784
rect 3283 26744 3608 26772
rect 3283 26741 3295 26744
rect 3237 26735 3295 26741
rect 3602 26732 3608 26744
rect 3660 26732 3666 26784
rect 4890 26732 4896 26784
rect 4948 26772 4954 26784
rect 7116 26781 7144 26812
rect 8846 26800 8852 26852
rect 8904 26800 8910 26852
rect 9582 26800 9588 26852
rect 9640 26800 9646 26852
rect 10410 26800 10416 26852
rect 10468 26840 10474 26852
rect 11716 26840 11744 26871
rect 12434 26868 12440 26920
rect 12492 26908 12498 26920
rect 12529 26911 12587 26917
rect 12529 26908 12541 26911
rect 12492 26880 12541 26908
rect 12492 26868 12498 26880
rect 12529 26877 12541 26880
rect 12575 26877 12587 26911
rect 12529 26871 12587 26877
rect 13848 26883 13876 26936
rect 14292 26917 14320 27004
rect 14369 26979 14427 26985
rect 14369 26945 14381 26979
rect 14415 26976 14427 26979
rect 15013 26979 15071 26985
rect 15013 26976 15025 26979
rect 14415 26948 15025 26976
rect 14415 26945 14427 26948
rect 14369 26939 14427 26945
rect 15013 26945 15025 26948
rect 15059 26945 15071 26979
rect 15120 26976 15148 27084
rect 15838 27072 15844 27124
rect 15896 27072 15902 27124
rect 15930 27072 15936 27124
rect 15988 27112 15994 27124
rect 18601 27115 18659 27121
rect 15988 27084 17540 27112
rect 15988 27072 15994 27084
rect 15197 27047 15255 27053
rect 15197 27013 15209 27047
rect 15243 27044 15255 27047
rect 17512 27044 17540 27084
rect 18601 27081 18613 27115
rect 18647 27112 18659 27115
rect 19058 27112 19064 27124
rect 18647 27084 19064 27112
rect 18647 27081 18659 27084
rect 18601 27075 18659 27081
rect 19058 27072 19064 27084
rect 19116 27072 19122 27124
rect 20901 27115 20959 27121
rect 20901 27081 20913 27115
rect 20947 27112 20959 27115
rect 21726 27112 21732 27124
rect 20947 27084 21732 27112
rect 20947 27081 20959 27084
rect 20901 27075 20959 27081
rect 21726 27072 21732 27084
rect 21784 27072 21790 27124
rect 21818 27072 21824 27124
rect 21876 27072 21882 27124
rect 22002 27072 22008 27124
rect 22060 27112 22066 27124
rect 22820 27115 22878 27121
rect 22060 27084 22600 27112
rect 22060 27072 22066 27084
rect 21836 27044 21864 27072
rect 15243 27016 16252 27044
rect 17512 27016 21864 27044
rect 15243 27013 15255 27016
rect 15197 27007 15255 27013
rect 16224 26976 16252 27016
rect 17313 26979 17371 26985
rect 17313 26976 17325 26979
rect 15120 26948 15608 26976
rect 16224 26948 17325 26976
rect 15013 26939 15071 26945
rect 14277 26911 14335 26917
rect 13848 26877 13921 26883
rect 10468 26812 13492 26840
rect 10468 26800 10474 26812
rect 5169 26775 5227 26781
rect 5169 26772 5181 26775
rect 4948 26744 5181 26772
rect 4948 26732 4954 26744
rect 5169 26741 5181 26744
rect 5215 26741 5227 26775
rect 5169 26735 5227 26741
rect 7101 26775 7159 26781
rect 7101 26741 7113 26775
rect 7147 26741 7159 26775
rect 7101 26735 7159 26741
rect 7190 26732 7196 26784
rect 7248 26772 7254 26784
rect 7469 26775 7527 26781
rect 7469 26772 7481 26775
rect 7248 26744 7481 26772
rect 7248 26732 7254 26744
rect 7469 26741 7481 26744
rect 7515 26741 7527 26775
rect 7469 26735 7527 26741
rect 10594 26732 10600 26784
rect 10652 26732 10658 26784
rect 10796 26781 10824 26812
rect 10781 26775 10839 26781
rect 10781 26741 10793 26775
rect 10827 26741 10839 26775
rect 10781 26735 10839 26741
rect 11882 26732 11888 26784
rect 11940 26732 11946 26784
rect 11974 26732 11980 26784
rect 12032 26732 12038 26784
rect 12710 26732 12716 26784
rect 12768 26732 12774 26784
rect 13464 26772 13492 26812
rect 13630 26800 13636 26852
rect 13688 26800 13694 26852
rect 13848 26843 13875 26877
rect 13909 26843 13921 26877
rect 14277 26877 14289 26911
rect 14323 26877 14335 26911
rect 14277 26871 14335 26877
rect 14553 26911 14611 26917
rect 14553 26877 14565 26911
rect 14599 26908 14611 26911
rect 14921 26911 14979 26917
rect 14921 26908 14933 26911
rect 14599 26880 14780 26908
rect 14599 26877 14611 26880
rect 14553 26871 14611 26877
rect 13848 26840 13921 26843
rect 14642 26840 14648 26852
rect 13848 26812 14648 26840
rect 14642 26800 14648 26812
rect 14700 26800 14706 26852
rect 14752 26784 14780 26880
rect 14844 26880 14933 26908
rect 14844 26852 14872 26880
rect 14921 26877 14933 26880
rect 14967 26877 14979 26911
rect 14921 26871 14979 26877
rect 15470 26868 15476 26920
rect 15528 26868 15534 26920
rect 15580 26917 15608 26948
rect 17313 26945 17325 26948
rect 17359 26945 17371 26979
rect 17313 26939 17371 26945
rect 17589 26979 17647 26985
rect 17589 26945 17601 26979
rect 17635 26976 17647 26979
rect 17678 26976 17684 26988
rect 17635 26948 17684 26976
rect 17635 26945 17647 26948
rect 17589 26939 17647 26945
rect 17678 26936 17684 26948
rect 17736 26936 17742 26988
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 21910 26976 21916 26988
rect 18104 26948 21916 26976
rect 18104 26936 18110 26948
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 22572 26985 22600 27084
rect 22820 27081 22832 27115
rect 22866 27112 22878 27115
rect 24118 27112 24124 27124
rect 22866 27084 24124 27112
rect 22866 27081 22878 27084
rect 22820 27075 22878 27081
rect 24118 27072 24124 27084
rect 24176 27072 24182 27124
rect 24305 27115 24363 27121
rect 24305 27081 24317 27115
rect 24351 27112 24363 27115
rect 24854 27112 24860 27124
rect 24351 27084 24860 27112
rect 24351 27081 24363 27084
rect 24305 27075 24363 27081
rect 24854 27072 24860 27084
rect 24912 27072 24918 27124
rect 24949 27115 25007 27121
rect 24949 27081 24961 27115
rect 24995 27112 25007 27115
rect 26326 27112 26332 27124
rect 24995 27084 26332 27112
rect 24995 27081 25007 27084
rect 24949 27075 25007 27081
rect 26326 27072 26332 27084
rect 26384 27072 26390 27124
rect 27801 27115 27859 27121
rect 27801 27081 27813 27115
rect 27847 27112 27859 27115
rect 30558 27112 30564 27124
rect 27847 27084 30564 27112
rect 27847 27081 27859 27084
rect 27801 27075 27859 27081
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 32582 27072 32588 27124
rect 32640 27112 32646 27124
rect 32953 27115 33011 27121
rect 32953 27112 32965 27115
rect 32640 27084 32965 27112
rect 32640 27072 32646 27084
rect 32953 27081 32965 27084
rect 32999 27081 33011 27115
rect 32953 27075 33011 27081
rect 33042 27072 33048 27124
rect 33100 27112 33106 27124
rect 33505 27115 33563 27121
rect 33505 27112 33517 27115
rect 33100 27084 33517 27112
rect 33100 27072 33106 27084
rect 33505 27081 33517 27084
rect 33551 27081 33563 27115
rect 33505 27075 33563 27081
rect 28353 27047 28411 27053
rect 28353 27044 28365 27047
rect 27356 27016 28365 27044
rect 22557 26979 22615 26985
rect 22557 26945 22569 26979
rect 22603 26976 22615 26979
rect 24026 26976 24032 26988
rect 22603 26948 24032 26976
rect 22603 26945 22615 26948
rect 22557 26939 22615 26945
rect 24026 26936 24032 26948
rect 24084 26976 24090 26988
rect 26053 26979 26111 26985
rect 26053 26976 26065 26979
rect 24084 26948 26065 26976
rect 24084 26936 24090 26948
rect 26053 26945 26065 26948
rect 26099 26945 26111 26979
rect 26053 26939 26111 26945
rect 27062 26936 27068 26988
rect 27120 26976 27126 26988
rect 27356 26976 27384 27016
rect 28353 27013 28365 27016
rect 28399 27013 28411 27047
rect 28353 27007 28411 27013
rect 31021 27047 31079 27053
rect 31021 27013 31033 27047
rect 31067 27044 31079 27047
rect 31067 27016 31340 27044
rect 31067 27013 31079 27016
rect 31021 27007 31079 27013
rect 27120 26948 27384 26976
rect 27120 26936 27126 26948
rect 28074 26936 28080 26988
rect 28132 26976 28138 26988
rect 29089 26979 29147 26985
rect 29089 26976 29101 26979
rect 28132 26948 29101 26976
rect 28132 26936 28138 26948
rect 29089 26945 29101 26948
rect 29135 26945 29147 26979
rect 29089 26939 29147 26945
rect 29178 26936 29184 26988
rect 29236 26976 29242 26988
rect 29273 26979 29331 26985
rect 29273 26976 29285 26979
rect 29236 26948 29285 26976
rect 29236 26936 29242 26948
rect 29273 26945 29285 26948
rect 29319 26976 29331 26979
rect 31205 26979 31263 26985
rect 31205 26976 31217 26979
rect 29319 26948 31217 26976
rect 29319 26945 29331 26948
rect 29273 26939 29331 26945
rect 31205 26945 31217 26948
rect 31251 26945 31263 26979
rect 31312 26976 31340 27016
rect 33134 27004 33140 27056
rect 33192 27004 33198 27056
rect 31846 26976 31852 26988
rect 31312 26948 31852 26976
rect 31205 26939 31263 26945
rect 31846 26936 31852 26948
rect 31904 26976 31910 26988
rect 32214 26976 32220 26988
rect 31904 26948 32220 26976
rect 31904 26936 31910 26948
rect 32214 26936 32220 26948
rect 32272 26936 32278 26988
rect 15565 26911 15623 26917
rect 15565 26877 15577 26911
rect 15611 26877 15623 26911
rect 15565 26871 15623 26877
rect 18693 26911 18751 26917
rect 18693 26877 18705 26911
rect 18739 26908 18751 26911
rect 20898 26908 20904 26920
rect 18739 26880 20904 26908
rect 18739 26877 18751 26880
rect 18693 26871 18751 26877
rect 20898 26868 20904 26880
rect 20956 26868 20962 26920
rect 21082 26868 21088 26920
rect 21140 26868 21146 26920
rect 21174 26868 21180 26920
rect 21232 26868 21238 26920
rect 21358 26868 21364 26920
rect 21416 26908 21422 26920
rect 21453 26911 21511 26917
rect 21453 26908 21465 26911
rect 21416 26880 21465 26908
rect 21416 26868 21422 26880
rect 21453 26877 21465 26880
rect 21499 26877 21511 26911
rect 21453 26871 21511 26877
rect 24397 26911 24455 26917
rect 24397 26877 24409 26911
rect 24443 26908 24455 26911
rect 24486 26908 24492 26920
rect 24443 26880 24492 26908
rect 24443 26877 24455 26880
rect 24397 26871 24455 26877
rect 14826 26800 14832 26852
rect 14884 26800 14890 26852
rect 15289 26843 15347 26849
rect 15289 26809 15301 26843
rect 15335 26840 15347 26843
rect 15654 26840 15660 26852
rect 15335 26812 15660 26840
rect 15335 26809 15347 26812
rect 15289 26803 15347 26809
rect 15654 26800 15660 26812
rect 15712 26800 15718 26852
rect 16298 26800 16304 26852
rect 16356 26800 16362 26852
rect 17218 26800 17224 26852
rect 17276 26840 17282 26852
rect 19058 26840 19064 26852
rect 17276 26812 19064 26840
rect 17276 26800 17282 26812
rect 19058 26800 19064 26812
rect 19116 26800 19122 26852
rect 21269 26843 21327 26849
rect 21269 26809 21281 26843
rect 21315 26840 21327 26843
rect 21634 26840 21640 26852
rect 21315 26812 21640 26840
rect 21315 26809 21327 26812
rect 21269 26803 21327 26809
rect 14182 26772 14188 26784
rect 13464 26744 14188 26772
rect 14182 26732 14188 26744
rect 14240 26732 14246 26784
rect 14734 26732 14740 26784
rect 14792 26772 14798 26784
rect 15387 26775 15445 26781
rect 15387 26772 15399 26775
rect 14792 26744 15399 26772
rect 14792 26732 14798 26744
rect 15387 26741 15399 26744
rect 15433 26741 15445 26775
rect 15387 26735 15445 26741
rect 20717 26775 20775 26781
rect 20717 26741 20729 26775
rect 20763 26772 20775 26775
rect 21284 26772 21312 26803
rect 21634 26800 21640 26812
rect 21692 26800 21698 26852
rect 23290 26800 23296 26852
rect 23348 26800 23354 26852
rect 20763 26744 21312 26772
rect 20763 26741 20775 26744
rect 20717 26735 20775 26741
rect 21910 26732 21916 26784
rect 21968 26772 21974 26784
rect 22186 26772 22192 26784
rect 21968 26744 22192 26772
rect 21968 26732 21974 26744
rect 22186 26732 22192 26744
rect 22244 26732 22250 26784
rect 22465 26775 22523 26781
rect 22465 26741 22477 26775
rect 22511 26772 22523 26775
rect 24412 26772 24440 26871
rect 24486 26868 24492 26880
rect 24544 26868 24550 26920
rect 24670 26868 24676 26920
rect 24728 26868 24734 26920
rect 24762 26868 24768 26920
rect 24820 26910 24826 26920
rect 24820 26882 24900 26910
rect 24820 26868 24826 26882
rect 24578 26800 24584 26852
rect 24636 26800 24642 26852
rect 24872 26840 24900 26882
rect 25682 26868 25688 26920
rect 25740 26868 25746 26920
rect 27893 26911 27951 26917
rect 27893 26877 27905 26911
rect 27939 26877 27951 26911
rect 27893 26871 27951 26877
rect 26234 26840 26240 26852
rect 24872 26812 26240 26840
rect 26234 26800 26240 26812
rect 26292 26800 26298 26852
rect 26326 26800 26332 26852
rect 26384 26800 26390 26852
rect 26878 26800 26884 26852
rect 26936 26800 26942 26852
rect 22511 26744 24440 26772
rect 22511 26741 22523 26744
rect 22465 26735 22523 26741
rect 24854 26732 24860 26784
rect 24912 26772 24918 26784
rect 25133 26775 25191 26781
rect 25133 26772 25145 26775
rect 24912 26744 25145 26772
rect 24912 26732 24918 26744
rect 25133 26741 25145 26744
rect 25179 26741 25191 26775
rect 25133 26735 25191 26741
rect 26970 26732 26976 26784
rect 27028 26772 27034 26784
rect 27908 26772 27936 26871
rect 28626 26868 28632 26920
rect 28684 26868 28690 26920
rect 30650 26868 30656 26920
rect 30708 26868 30714 26920
rect 33152 26908 33180 27004
rect 33229 26911 33287 26917
rect 33229 26908 33241 26911
rect 33152 26880 33241 26908
rect 33229 26877 33241 26880
rect 33275 26908 33287 26911
rect 33410 26908 33416 26920
rect 33275 26880 33416 26908
rect 33275 26877 33287 26880
rect 33229 26871 33287 26877
rect 33410 26868 33416 26880
rect 33468 26868 33474 26920
rect 28721 26843 28779 26849
rect 28721 26809 28733 26843
rect 28767 26840 28779 26843
rect 28767 26812 29316 26840
rect 28767 26809 28779 26812
rect 28721 26803 28779 26809
rect 29288 26784 29316 26812
rect 29546 26800 29552 26852
rect 29604 26800 29610 26852
rect 31478 26800 31484 26852
rect 31536 26800 31542 26852
rect 33137 26843 33195 26849
rect 33137 26840 33149 26843
rect 32706 26812 33149 26840
rect 33137 26809 33149 26812
rect 33183 26809 33195 26843
rect 33137 26803 33195 26809
rect 27028 26744 27936 26772
rect 27028 26732 27034 26744
rect 27982 26732 27988 26784
rect 28040 26772 28046 26784
rect 28077 26775 28135 26781
rect 28077 26772 28089 26775
rect 28040 26744 28089 26772
rect 28040 26732 28046 26744
rect 28077 26741 28089 26744
rect 28123 26741 28135 26775
rect 28077 26735 28135 26741
rect 29270 26732 29276 26784
rect 29328 26732 29334 26784
rect 32490 26732 32496 26784
rect 32548 26772 32554 26784
rect 33873 26775 33931 26781
rect 33873 26772 33885 26775
rect 32548 26744 33885 26772
rect 32548 26732 32554 26744
rect 33873 26741 33885 26744
rect 33919 26741 33931 26775
rect 33873 26735 33931 26741
rect 2760 26682 34316 26704
rect 2760 26630 7210 26682
rect 7262 26630 7274 26682
rect 7326 26630 7338 26682
rect 7390 26630 7402 26682
rect 7454 26630 7466 26682
rect 7518 26630 15099 26682
rect 15151 26630 15163 26682
rect 15215 26630 15227 26682
rect 15279 26630 15291 26682
rect 15343 26630 15355 26682
rect 15407 26630 22988 26682
rect 23040 26630 23052 26682
rect 23104 26630 23116 26682
rect 23168 26630 23180 26682
rect 23232 26630 23244 26682
rect 23296 26630 30877 26682
rect 30929 26630 30941 26682
rect 30993 26630 31005 26682
rect 31057 26630 31069 26682
rect 31121 26630 31133 26682
rect 31185 26630 34316 26682
rect 2760 26608 34316 26630
rect 4525 26571 4583 26577
rect 4525 26537 4537 26571
rect 4571 26568 4583 26571
rect 4614 26568 4620 26580
rect 4571 26540 4620 26568
rect 4571 26537 4583 26540
rect 4525 26531 4583 26537
rect 4614 26528 4620 26540
rect 4672 26528 4678 26580
rect 5718 26528 5724 26580
rect 5776 26528 5782 26580
rect 5810 26528 5816 26580
rect 5868 26528 5874 26580
rect 6178 26528 6184 26580
rect 6236 26568 6242 26580
rect 7101 26571 7159 26577
rect 7101 26568 7113 26571
rect 6236 26540 7113 26568
rect 6236 26528 6242 26540
rect 7101 26537 7113 26540
rect 7147 26537 7159 26571
rect 7101 26531 7159 26537
rect 8846 26528 8852 26580
rect 8904 26568 8910 26580
rect 9309 26571 9367 26577
rect 9309 26568 9321 26571
rect 8904 26540 9321 26568
rect 8904 26528 8910 26540
rect 9309 26537 9321 26540
rect 9355 26537 9367 26571
rect 9309 26531 9367 26537
rect 10686 26528 10692 26580
rect 10744 26528 10750 26580
rect 11422 26528 11428 26580
rect 11480 26528 11486 26580
rect 11882 26528 11888 26580
rect 11940 26568 11946 26580
rect 12437 26571 12495 26577
rect 12437 26568 12449 26571
rect 11940 26540 12449 26568
rect 11940 26528 11946 26540
rect 12437 26537 12449 26540
rect 12483 26537 12495 26571
rect 12437 26531 12495 26537
rect 13630 26528 13636 26580
rect 13688 26528 13694 26580
rect 13722 26528 13728 26580
rect 13780 26528 13786 26580
rect 13817 26571 13875 26577
rect 13817 26537 13829 26571
rect 13863 26568 13875 26571
rect 13906 26568 13912 26580
rect 13863 26540 13912 26568
rect 13863 26537 13875 26540
rect 13817 26531 13875 26537
rect 13906 26528 13912 26540
rect 13964 26528 13970 26580
rect 14090 26528 14096 26580
rect 14148 26528 14154 26580
rect 15381 26571 15439 26577
rect 15381 26537 15393 26571
rect 15427 26568 15439 26571
rect 15746 26568 15752 26580
rect 15427 26540 15752 26568
rect 15427 26537 15439 26540
rect 15381 26531 15439 26537
rect 15746 26528 15752 26540
rect 15804 26528 15810 26580
rect 16298 26528 16304 26580
rect 16356 26568 16362 26580
rect 16485 26571 16543 26577
rect 16485 26568 16497 26571
rect 16356 26540 16497 26568
rect 16356 26528 16362 26540
rect 16485 26537 16497 26540
rect 16531 26537 16543 26571
rect 16485 26531 16543 26537
rect 17497 26571 17555 26577
rect 17497 26537 17509 26571
rect 17543 26568 17555 26571
rect 17586 26568 17592 26580
rect 17543 26540 17592 26568
rect 17543 26537 17555 26540
rect 17497 26531 17555 26537
rect 17586 26528 17592 26540
rect 17644 26528 17650 26580
rect 22925 26571 22983 26577
rect 22925 26537 22937 26571
rect 22971 26568 22983 26571
rect 24578 26568 24584 26580
rect 22971 26540 24584 26568
rect 22971 26537 22983 26540
rect 22925 26531 22983 26537
rect 5736 26500 5764 26528
rect 5566 26472 5764 26500
rect 5828 26500 5856 26528
rect 5997 26503 6055 26509
rect 5997 26500 6009 26503
rect 5828 26472 6009 26500
rect 5997 26469 6009 26472
rect 6043 26469 6055 26503
rect 5997 26463 6055 26469
rect 4246 26392 4252 26444
rect 4304 26392 4310 26444
rect 6273 26435 6331 26441
rect 6273 26401 6285 26435
rect 6319 26432 6331 26435
rect 8018 26432 8024 26444
rect 6319 26404 8024 26432
rect 6319 26401 6331 26404
rect 6273 26395 6331 26401
rect 8018 26392 8024 26404
rect 8076 26392 8082 26444
rect 10873 26435 10931 26441
rect 10873 26401 10885 26435
rect 10919 26432 10931 26435
rect 11440 26432 11468 26528
rect 12345 26503 12403 26509
rect 12345 26469 12357 26503
rect 12391 26500 12403 26503
rect 12897 26503 12955 26509
rect 12897 26500 12909 26503
rect 12391 26472 12909 26500
rect 12391 26469 12403 26472
rect 12345 26463 12403 26469
rect 12897 26469 12909 26472
rect 12943 26469 12955 26503
rect 13648 26500 13676 26528
rect 12897 26463 12955 26469
rect 13004 26472 13676 26500
rect 10919 26404 11468 26432
rect 10919 26401 10931 26404
rect 10873 26395 10931 26401
rect 11698 26392 11704 26444
rect 11756 26392 11762 26444
rect 12434 26432 12440 26444
rect 12406 26392 12440 26432
rect 12492 26392 12498 26444
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 13004 26441 13032 26472
rect 12805 26435 12863 26441
rect 12805 26432 12817 26435
rect 12676 26404 12817 26432
rect 12676 26392 12682 26404
rect 12805 26401 12817 26404
rect 12851 26401 12863 26435
rect 12805 26395 12863 26401
rect 12989 26435 13047 26441
rect 12989 26401 13001 26435
rect 13035 26401 13047 26435
rect 12989 26395 13047 26401
rect 13633 26435 13691 26441
rect 13633 26401 13645 26435
rect 13679 26432 13691 26435
rect 13740 26432 13768 26528
rect 14108 26441 14136 26528
rect 20901 26503 20959 26509
rect 20901 26500 20913 26503
rect 20470 26472 20913 26500
rect 20901 26469 20913 26472
rect 20947 26469 20959 26503
rect 20901 26463 20959 26469
rect 21634 26460 21640 26512
rect 21692 26500 21698 26512
rect 22940 26500 22968 26531
rect 24578 26528 24584 26540
rect 24636 26528 24642 26580
rect 26878 26528 26884 26580
rect 26936 26528 26942 26580
rect 27154 26528 27160 26580
rect 27212 26528 27218 26580
rect 29549 26571 29607 26577
rect 29549 26537 29561 26571
rect 29595 26568 29607 26571
rect 30098 26568 30104 26580
rect 29595 26540 30104 26568
rect 29595 26537 29607 26540
rect 29549 26531 29607 26537
rect 30098 26528 30104 26540
rect 30156 26528 30162 26580
rect 31478 26528 31484 26580
rect 31536 26528 31542 26580
rect 32030 26528 32036 26580
rect 32088 26528 32094 26580
rect 21692 26472 22968 26500
rect 21692 26460 21698 26472
rect 23842 26460 23848 26512
rect 23900 26500 23906 26512
rect 24121 26503 24179 26509
rect 24121 26500 24133 26503
rect 23900 26472 24133 26500
rect 23900 26460 23906 26472
rect 24121 26469 24133 26472
rect 24167 26469 24179 26503
rect 24121 26463 24179 26469
rect 24765 26503 24823 26509
rect 24765 26469 24777 26503
rect 24811 26500 24823 26503
rect 25866 26500 25872 26512
rect 24811 26472 25872 26500
rect 24811 26469 24823 26472
rect 24765 26463 24823 26469
rect 25866 26460 25872 26472
rect 25924 26500 25930 26512
rect 25924 26472 31754 26500
rect 25924 26460 25930 26472
rect 13679 26404 13768 26432
rect 14093 26435 14151 26441
rect 13679 26401 13691 26404
rect 13633 26395 13691 26401
rect 14093 26401 14105 26435
rect 14139 26401 14151 26435
rect 14093 26395 14151 26401
rect 3234 26324 3240 26376
rect 3292 26324 3298 26376
rect 6914 26324 6920 26376
rect 6972 26324 6978 26376
rect 7650 26324 7656 26376
rect 7708 26324 7714 26376
rect 9858 26324 9864 26376
rect 9916 26324 9922 26376
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26364 11391 26367
rect 11716 26364 11744 26392
rect 11379 26336 11744 26364
rect 11379 26333 11391 26336
rect 11333 26327 11391 26333
rect 11882 26256 11888 26308
rect 11940 26256 11946 26308
rect 11977 26299 12035 26305
rect 11977 26265 11989 26299
rect 12023 26296 12035 26299
rect 12406 26296 12434 26392
rect 12529 26367 12587 26373
rect 12529 26333 12541 26367
rect 12575 26333 12587 26367
rect 12820 26364 12848 26395
rect 14182 26392 14188 26444
rect 14240 26432 14246 26444
rect 14553 26435 14611 26441
rect 14553 26432 14565 26435
rect 14240 26404 14565 26432
rect 14240 26392 14246 26404
rect 14553 26401 14565 26404
rect 14599 26401 14611 26435
rect 14553 26395 14611 26401
rect 14734 26392 14740 26444
rect 14792 26392 14798 26444
rect 15562 26392 15568 26444
rect 15620 26392 15626 26444
rect 16574 26392 16580 26444
rect 16632 26432 16638 26444
rect 17862 26432 17868 26444
rect 16632 26404 17868 26432
rect 16632 26392 16638 26404
rect 17862 26392 17868 26404
rect 17920 26392 17926 26444
rect 18966 26392 18972 26444
rect 19024 26392 19030 26444
rect 20993 26435 21051 26441
rect 20993 26401 21005 26435
rect 21039 26401 21051 26435
rect 20993 26395 21051 26401
rect 12820 26336 14228 26364
rect 12529 26327 12587 26333
rect 12023 26268 12434 26296
rect 12544 26296 12572 26327
rect 13906 26296 13912 26308
rect 12544 26268 13912 26296
rect 12023 26265 12035 26268
rect 11977 26259 12035 26265
rect 13906 26256 13912 26268
rect 13964 26256 13970 26308
rect 6362 26188 6368 26240
rect 6420 26188 6426 26240
rect 14200 26237 14228 26336
rect 18138 26324 18144 26376
rect 18196 26324 18202 26376
rect 19242 26324 19248 26376
rect 19300 26324 19306 26376
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 21008 26364 21036 26395
rect 22186 26392 22192 26444
rect 22244 26392 22250 26444
rect 23382 26392 23388 26444
rect 23440 26432 23446 26444
rect 24854 26432 24860 26444
rect 23440 26404 24860 26432
rect 23440 26392 23446 26404
rect 24854 26392 24860 26404
rect 24912 26392 24918 26444
rect 26786 26392 26792 26444
rect 26844 26392 26850 26444
rect 27065 26435 27123 26441
rect 27065 26401 27077 26435
rect 27111 26401 27123 26435
rect 27065 26395 27123 26401
rect 20956 26336 21036 26364
rect 20956 26324 20962 26336
rect 23474 26324 23480 26376
rect 23532 26324 23538 26376
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26364 24639 26367
rect 24946 26364 24952 26376
rect 24627 26336 24952 26364
rect 24627 26333 24639 26336
rect 24581 26327 24639 26333
rect 17402 26256 17408 26308
rect 17460 26296 17466 26308
rect 18046 26296 18052 26308
rect 17460 26268 18052 26296
rect 17460 26256 17466 26268
rect 18046 26256 18052 26268
rect 18104 26256 18110 26308
rect 20717 26299 20775 26305
rect 20717 26265 20729 26299
rect 20763 26296 20775 26299
rect 23293 26299 23351 26305
rect 20763 26268 22508 26296
rect 20763 26265 20775 26268
rect 20717 26259 20775 26265
rect 14185 26231 14243 26237
rect 14185 26197 14197 26231
rect 14231 26197 14243 26231
rect 14185 26191 14243 26197
rect 14737 26231 14795 26237
rect 14737 26197 14749 26231
rect 14783 26228 14795 26231
rect 14826 26228 14832 26240
rect 14783 26200 14832 26228
rect 14783 26197 14795 26200
rect 14737 26191 14795 26197
rect 14826 26188 14832 26200
rect 14884 26188 14890 26240
rect 15838 26188 15844 26240
rect 15896 26188 15902 26240
rect 17037 26231 17095 26237
rect 17037 26197 17049 26231
rect 17083 26228 17095 26231
rect 17126 26228 17132 26240
rect 17083 26200 17132 26228
rect 17083 26197 17095 26200
rect 17037 26191 17095 26197
rect 17126 26188 17132 26200
rect 17184 26188 17190 26240
rect 21542 26188 21548 26240
rect 21600 26188 21606 26240
rect 22480 26228 22508 26268
rect 23293 26265 23305 26299
rect 23339 26296 23351 26299
rect 24596 26296 24624 26327
rect 24946 26324 24952 26336
rect 25004 26324 25010 26376
rect 25869 26367 25927 26373
rect 25869 26333 25881 26367
rect 25915 26333 25927 26367
rect 25869 26327 25927 26333
rect 23339 26268 24624 26296
rect 25225 26299 25283 26305
rect 23339 26265 23351 26268
rect 23293 26259 23351 26265
rect 25225 26265 25237 26299
rect 25271 26296 25283 26299
rect 25884 26296 25912 26327
rect 25958 26324 25964 26376
rect 26016 26364 26022 26376
rect 26605 26367 26663 26373
rect 26605 26364 26617 26367
rect 26016 26336 26617 26364
rect 26016 26324 26022 26336
rect 26605 26333 26617 26336
rect 26651 26333 26663 26367
rect 27080 26364 27108 26395
rect 27154 26392 27160 26444
rect 27212 26432 27218 26444
rect 27249 26435 27307 26441
rect 27249 26432 27261 26435
rect 27212 26404 27261 26432
rect 27212 26392 27218 26404
rect 27249 26401 27261 26404
rect 27295 26401 27307 26435
rect 27249 26395 27307 26401
rect 28074 26392 28080 26444
rect 28132 26392 28138 26444
rect 28166 26392 28172 26444
rect 28224 26432 28230 26444
rect 28353 26435 28411 26441
rect 28353 26432 28365 26435
rect 28224 26404 28365 26432
rect 28224 26392 28230 26404
rect 28353 26401 28365 26404
rect 28399 26401 28411 26435
rect 28353 26395 28411 26401
rect 28445 26435 28503 26441
rect 28445 26401 28457 26435
rect 28491 26432 28503 26435
rect 29917 26435 29975 26441
rect 29917 26432 29929 26435
rect 28491 26404 29929 26432
rect 28491 26401 28503 26404
rect 28445 26395 28503 26401
rect 29917 26401 29929 26404
rect 29963 26432 29975 26435
rect 30377 26435 30435 26441
rect 30377 26432 30389 26435
rect 29963 26404 30389 26432
rect 29963 26401 29975 26404
rect 29917 26395 29975 26401
rect 30377 26401 30389 26404
rect 30423 26401 30435 26435
rect 30377 26395 30435 26401
rect 27985 26367 28043 26373
rect 27985 26364 27997 26367
rect 26605 26327 26663 26333
rect 26804 26336 27997 26364
rect 26804 26308 26832 26336
rect 27985 26333 27997 26336
rect 28031 26333 28043 26367
rect 27985 26327 28043 26333
rect 29181 26367 29239 26373
rect 29181 26333 29193 26367
rect 29227 26333 29239 26367
rect 29181 26327 29239 26333
rect 30009 26367 30067 26373
rect 30009 26333 30021 26367
rect 30055 26333 30067 26367
rect 30009 26327 30067 26333
rect 30193 26367 30251 26373
rect 30193 26333 30205 26367
rect 30239 26364 30251 26367
rect 30558 26364 30564 26376
rect 30239 26336 30564 26364
rect 30239 26333 30251 26336
rect 30193 26327 30251 26333
rect 25271 26268 25912 26296
rect 25271 26265 25283 26268
rect 25225 26259 25283 26265
rect 26786 26256 26792 26308
rect 26844 26256 26850 26308
rect 27801 26299 27859 26305
rect 27801 26265 27813 26299
rect 27847 26296 27859 26299
rect 29196 26296 29224 26327
rect 27847 26268 29224 26296
rect 30024 26296 30052 26327
rect 30558 26324 30564 26336
rect 30616 26324 30622 26376
rect 30926 26324 30932 26376
rect 30984 26324 30990 26376
rect 31726 26364 31754 26472
rect 32048 26441 32076 26528
rect 32033 26435 32091 26441
rect 32033 26401 32045 26435
rect 32079 26401 32091 26435
rect 32033 26395 32091 26401
rect 32217 26435 32275 26441
rect 32217 26401 32229 26435
rect 32263 26401 32275 26435
rect 32217 26395 32275 26401
rect 32232 26364 32260 26395
rect 31726 26336 32260 26364
rect 33042 26324 33048 26376
rect 33100 26324 33106 26376
rect 31846 26296 31852 26308
rect 30024 26268 31852 26296
rect 27847 26265 27859 26268
rect 27801 26259 27859 26265
rect 31846 26256 31852 26268
rect 31904 26256 31910 26308
rect 24302 26228 24308 26240
rect 22480 26200 24308 26228
rect 24302 26188 24308 26200
rect 24360 26188 24366 26240
rect 24854 26188 24860 26240
rect 24912 26228 24918 26240
rect 25317 26231 25375 26237
rect 25317 26228 25329 26231
rect 24912 26200 25329 26228
rect 24912 26188 24918 26200
rect 25317 26197 25329 26200
rect 25363 26197 25375 26231
rect 25317 26191 25375 26197
rect 25406 26188 25412 26240
rect 25464 26228 25470 26240
rect 26050 26228 26056 26240
rect 25464 26200 26056 26228
rect 25464 26188 25470 26200
rect 26050 26188 26056 26200
rect 26108 26188 26114 26240
rect 26234 26188 26240 26240
rect 26292 26228 26298 26240
rect 27525 26231 27583 26237
rect 27525 26228 27537 26231
rect 26292 26200 27537 26228
rect 26292 26188 26298 26200
rect 27525 26197 27537 26200
rect 27571 26197 27583 26231
rect 27525 26191 27583 26197
rect 28166 26188 28172 26240
rect 28224 26228 28230 26240
rect 28629 26231 28687 26237
rect 28629 26228 28641 26231
rect 28224 26200 28641 26228
rect 28224 26188 28230 26200
rect 28629 26197 28641 26200
rect 28675 26197 28687 26231
rect 28629 26191 28687 26197
rect 2760 26138 34316 26160
rect 2760 26086 6550 26138
rect 6602 26086 6614 26138
rect 6666 26086 6678 26138
rect 6730 26086 6742 26138
rect 6794 26086 6806 26138
rect 6858 26086 14439 26138
rect 14491 26086 14503 26138
rect 14555 26086 14567 26138
rect 14619 26086 14631 26138
rect 14683 26086 14695 26138
rect 14747 26086 22328 26138
rect 22380 26086 22392 26138
rect 22444 26086 22456 26138
rect 22508 26086 22520 26138
rect 22572 26086 22584 26138
rect 22636 26086 30217 26138
rect 30269 26086 30281 26138
rect 30333 26086 30345 26138
rect 30397 26086 30409 26138
rect 30461 26086 30473 26138
rect 30525 26086 34316 26138
rect 2760 26064 34316 26086
rect 7469 26027 7527 26033
rect 7469 25993 7481 26027
rect 7515 26024 7527 26027
rect 7650 26024 7656 26036
rect 7515 25996 7656 26024
rect 7515 25993 7527 25996
rect 7469 25987 7527 25993
rect 7650 25984 7656 25996
rect 7708 25984 7714 26036
rect 9585 26027 9643 26033
rect 9585 25993 9597 26027
rect 9631 26024 9643 26027
rect 9858 26024 9864 26036
rect 9631 25996 9864 26024
rect 9631 25993 9643 25996
rect 9585 25987 9643 25993
rect 9858 25984 9864 25996
rect 9916 25984 9922 26036
rect 10686 25984 10692 26036
rect 10744 25984 10750 26036
rect 12618 25984 12624 26036
rect 12676 26024 12682 26036
rect 13633 26027 13691 26033
rect 13633 26024 13645 26027
rect 12676 25996 13645 26024
rect 12676 25984 12682 25996
rect 13633 25993 13645 25996
rect 13679 25993 13691 26027
rect 13633 25987 13691 25993
rect 19242 25984 19248 26036
rect 19300 25984 19306 26036
rect 22830 25984 22836 26036
rect 22888 26024 22894 26036
rect 23290 26024 23296 26036
rect 22888 25996 23296 26024
rect 22888 25984 22894 25996
rect 23290 25984 23296 25996
rect 23348 25984 23354 26036
rect 23952 25996 25452 26024
rect 4982 25888 4988 25900
rect 3988 25860 4988 25888
rect 3988 25829 4016 25860
rect 4982 25848 4988 25860
rect 5040 25848 5046 25900
rect 5997 25891 6055 25897
rect 5997 25857 6009 25891
rect 6043 25888 6055 25891
rect 6362 25888 6368 25900
rect 6043 25860 6368 25888
rect 6043 25857 6055 25860
rect 5997 25851 6055 25857
rect 6362 25848 6368 25860
rect 6420 25848 6426 25900
rect 7650 25848 7656 25900
rect 7708 25888 7714 25900
rect 10318 25888 10324 25900
rect 7708 25860 7788 25888
rect 7708 25848 7714 25860
rect 3973 25823 4031 25829
rect 3973 25789 3985 25823
rect 4019 25789 4031 25823
rect 3973 25783 4031 25789
rect 4798 25780 4804 25832
rect 4856 25820 4862 25832
rect 7760 25829 7788 25860
rect 9876 25860 10324 25888
rect 9876 25829 9904 25860
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 10704 25888 10732 25984
rect 13538 25916 13544 25968
rect 13596 25956 13602 25968
rect 13596 25928 13860 25956
rect 13596 25916 13602 25928
rect 10520 25860 10732 25888
rect 11701 25891 11759 25897
rect 5721 25823 5779 25829
rect 5721 25820 5733 25823
rect 4856 25792 5733 25820
rect 4856 25780 4862 25792
rect 5721 25789 5733 25792
rect 5767 25789 5779 25823
rect 5721 25783 5779 25789
rect 7745 25823 7803 25829
rect 7745 25789 7757 25823
rect 7791 25789 7803 25823
rect 7745 25783 7803 25789
rect 9861 25823 9919 25829
rect 9861 25789 9873 25823
rect 9907 25789 9919 25823
rect 9861 25783 9919 25789
rect 10137 25823 10195 25829
rect 10137 25789 10149 25823
rect 10183 25820 10195 25823
rect 10520 25820 10548 25860
rect 11701 25857 11713 25891
rect 11747 25888 11759 25891
rect 13446 25888 13452 25900
rect 11747 25860 13452 25888
rect 11747 25857 11759 25860
rect 11701 25851 11759 25857
rect 13446 25848 13452 25860
rect 13504 25848 13510 25900
rect 10183 25792 10548 25820
rect 10183 25789 10195 25792
rect 10137 25783 10195 25789
rect 10594 25780 10600 25832
rect 10652 25780 10658 25832
rect 10686 25780 10692 25832
rect 10744 25780 10750 25832
rect 10965 25823 11023 25829
rect 10965 25789 10977 25823
rect 11011 25820 11023 25823
rect 11054 25820 11060 25832
rect 11011 25792 11060 25820
rect 11011 25789 11023 25792
rect 10965 25783 11023 25789
rect 11054 25780 11060 25792
rect 11112 25780 11118 25832
rect 13541 25823 13599 25829
rect 13541 25789 13553 25823
rect 13587 25820 13599 25823
rect 13630 25820 13636 25832
rect 13587 25792 13636 25820
rect 13587 25789 13599 25792
rect 13541 25783 13599 25789
rect 13630 25780 13636 25792
rect 13688 25780 13694 25832
rect 13722 25780 13728 25832
rect 13780 25780 13786 25832
rect 13832 25829 13860 25928
rect 17402 25916 17408 25968
rect 17460 25956 17466 25968
rect 18325 25959 18383 25965
rect 18325 25956 18337 25959
rect 17460 25928 18337 25956
rect 17460 25916 17466 25928
rect 18325 25925 18337 25928
rect 18371 25925 18383 25959
rect 18325 25919 18383 25925
rect 14826 25888 14832 25900
rect 13924 25860 14832 25888
rect 13924 25829 13952 25860
rect 14826 25848 14832 25860
rect 14884 25848 14890 25900
rect 17497 25891 17555 25897
rect 17497 25857 17509 25891
rect 17543 25888 17555 25891
rect 17678 25888 17684 25900
rect 17543 25860 17684 25888
rect 17543 25857 17555 25860
rect 17497 25851 17555 25857
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 17862 25848 17868 25900
rect 17920 25888 17926 25900
rect 17920 25860 18460 25888
rect 17920 25848 17926 25860
rect 13817 25823 13875 25829
rect 13817 25789 13829 25823
rect 13863 25789 13875 25823
rect 13817 25783 13875 25789
rect 13909 25823 13967 25829
rect 13909 25789 13921 25823
rect 13955 25789 13967 25823
rect 13909 25783 13967 25789
rect 14093 25823 14151 25829
rect 14093 25789 14105 25823
rect 14139 25820 14151 25823
rect 14737 25823 14795 25829
rect 14737 25820 14749 25823
rect 14139 25792 14749 25820
rect 14139 25789 14151 25792
rect 14093 25783 14151 25789
rect 14737 25789 14749 25792
rect 14783 25789 14795 25823
rect 14737 25783 14795 25789
rect 15565 25823 15623 25829
rect 15565 25789 15577 25823
rect 15611 25820 15623 25823
rect 16390 25820 16396 25832
rect 15611 25792 16396 25820
rect 15611 25789 15623 25792
rect 15565 25783 15623 25789
rect 16390 25780 16396 25792
rect 16448 25780 16454 25832
rect 17126 25780 17132 25832
rect 17184 25820 17190 25832
rect 17773 25823 17831 25829
rect 17773 25820 17785 25823
rect 17184 25792 17785 25820
rect 17184 25780 17190 25792
rect 17773 25789 17785 25792
rect 17819 25789 17831 25823
rect 17773 25783 17831 25789
rect 18046 25780 18052 25832
rect 18104 25820 18110 25832
rect 18432 25829 18460 25860
rect 21542 25848 21548 25900
rect 21600 25848 21606 25900
rect 23017 25891 23075 25897
rect 23017 25857 23029 25891
rect 23063 25888 23075 25891
rect 23845 25891 23903 25897
rect 23845 25888 23857 25891
rect 23063 25860 23857 25888
rect 23063 25857 23075 25860
rect 23017 25851 23075 25857
rect 23845 25857 23857 25860
rect 23891 25888 23903 25891
rect 23952 25888 23980 25996
rect 25424 25956 25452 25996
rect 25866 25984 25872 26036
rect 25924 25984 25930 26036
rect 26053 26027 26111 26033
rect 26053 25993 26065 26027
rect 26099 26024 26111 26027
rect 26326 26024 26332 26036
rect 26099 25996 26332 26024
rect 26099 25993 26111 25996
rect 26053 25987 26111 25993
rect 26326 25984 26332 25996
rect 26384 25984 26390 26036
rect 26418 25984 26424 26036
rect 26476 25984 26482 26036
rect 27065 26027 27123 26033
rect 27065 25993 27077 26027
rect 27111 26024 27123 26027
rect 27890 26024 27896 26036
rect 27111 25996 27896 26024
rect 27111 25993 27123 25996
rect 27065 25987 27123 25993
rect 27890 25984 27896 25996
rect 27948 25984 27954 26036
rect 29365 26027 29423 26033
rect 29365 25993 29377 26027
rect 29411 26024 29423 26027
rect 30926 26024 30932 26036
rect 29411 25996 30932 26024
rect 29411 25993 29423 25996
rect 29365 25987 29423 25993
rect 30926 25984 30932 25996
rect 30984 25984 30990 26036
rect 26436 25956 26464 25984
rect 25424 25928 26464 25956
rect 26510 25916 26516 25968
rect 26568 25956 26574 25968
rect 27338 25956 27344 25968
rect 26568 25928 27344 25956
rect 26568 25916 26574 25928
rect 27338 25916 27344 25928
rect 27396 25916 27402 25968
rect 28994 25916 29000 25968
rect 29052 25916 29058 25968
rect 23891 25860 23980 25888
rect 23891 25857 23903 25860
rect 23845 25851 23903 25857
rect 24026 25848 24032 25900
rect 24084 25888 24090 25900
rect 24121 25891 24179 25897
rect 24121 25888 24133 25891
rect 24084 25860 24133 25888
rect 24084 25848 24090 25860
rect 24121 25857 24133 25860
rect 24167 25857 24179 25891
rect 24121 25851 24179 25857
rect 24397 25891 24455 25897
rect 24397 25857 24409 25891
rect 24443 25888 24455 25891
rect 24854 25888 24860 25900
rect 24443 25860 24860 25888
rect 24443 25857 24455 25860
rect 24397 25851 24455 25857
rect 24854 25848 24860 25860
rect 24912 25848 24918 25900
rect 27617 25891 27675 25897
rect 26344 25860 27568 25888
rect 18141 25823 18199 25829
rect 18141 25820 18153 25823
rect 18104 25792 18153 25820
rect 18104 25780 18110 25792
rect 18141 25789 18153 25792
rect 18187 25789 18199 25823
rect 18141 25783 18199 25789
rect 18417 25823 18475 25829
rect 18417 25789 18429 25823
rect 18463 25789 18475 25823
rect 18417 25783 18475 25789
rect 18693 25823 18751 25829
rect 18693 25789 18705 25823
rect 18739 25789 18751 25823
rect 18693 25783 18751 25789
rect 19061 25823 19119 25829
rect 19061 25789 19073 25823
rect 19107 25820 19119 25823
rect 19150 25820 19156 25832
rect 19107 25792 19156 25820
rect 19107 25789 19119 25792
rect 19061 25783 19119 25789
rect 7653 25755 7711 25761
rect 7653 25752 7665 25755
rect 7222 25724 7665 25752
rect 7653 25721 7665 25724
rect 7699 25721 7711 25755
rect 7653 25715 7711 25721
rect 9585 25755 9643 25761
rect 9585 25721 9597 25755
rect 9631 25752 9643 25755
rect 10612 25752 10640 25780
rect 9631 25724 10640 25752
rect 9631 25721 9643 25724
rect 9585 25715 9643 25721
rect 3878 25644 3884 25696
rect 3936 25644 3942 25696
rect 9769 25687 9827 25693
rect 9769 25653 9781 25687
rect 9815 25684 9827 25687
rect 10045 25687 10103 25693
rect 10045 25684 10057 25687
rect 9815 25656 10057 25684
rect 9815 25653 9827 25656
rect 9769 25647 9827 25653
rect 10045 25653 10057 25656
rect 10091 25653 10103 25687
rect 10045 25647 10103 25653
rect 10410 25644 10416 25696
rect 10468 25684 10474 25696
rect 10689 25687 10747 25693
rect 10689 25684 10701 25687
rect 10468 25656 10701 25684
rect 10468 25644 10474 25656
rect 10689 25653 10701 25656
rect 10735 25653 10747 25687
rect 11072 25684 11100 25780
rect 11974 25712 11980 25764
rect 12032 25712 12038 25764
rect 13262 25752 13268 25764
rect 13202 25724 13268 25752
rect 13262 25712 13268 25724
rect 13320 25712 13326 25764
rect 12066 25684 12072 25696
rect 11072 25656 12072 25684
rect 10689 25647 10747 25653
rect 12066 25644 12072 25656
rect 12124 25644 12130 25696
rect 13449 25687 13507 25693
rect 13449 25653 13461 25687
rect 13495 25684 13507 25687
rect 13740 25684 13768 25780
rect 15470 25712 15476 25764
rect 15528 25752 15534 25764
rect 15749 25755 15807 25761
rect 15749 25752 15761 25755
rect 15528 25724 15761 25752
rect 15528 25712 15534 25724
rect 15749 25721 15761 25724
rect 15795 25752 15807 25755
rect 15838 25752 15844 25764
rect 15795 25724 15844 25752
rect 15795 25721 15807 25724
rect 15749 25715 15807 25721
rect 15838 25712 15844 25724
rect 15896 25712 15902 25764
rect 16666 25712 16672 25764
rect 16724 25752 16730 25764
rect 17865 25755 17923 25761
rect 17865 25752 17877 25755
rect 16724 25724 17877 25752
rect 16724 25712 16730 25724
rect 17865 25721 17877 25724
rect 17911 25721 17923 25755
rect 17865 25715 17923 25721
rect 17957 25755 18015 25761
rect 17957 25721 17969 25755
rect 18003 25752 18015 25755
rect 18003 25724 18552 25752
rect 18003 25721 18015 25724
rect 17957 25715 18015 25721
rect 18524 25696 18552 25724
rect 13495 25656 13768 25684
rect 13495 25653 13507 25656
rect 13449 25647 13507 25653
rect 14182 25644 14188 25696
rect 14240 25644 14246 25696
rect 14458 25644 14464 25696
rect 14516 25684 14522 25696
rect 14921 25687 14979 25693
rect 14921 25684 14933 25687
rect 14516 25656 14933 25684
rect 14516 25644 14522 25656
rect 14921 25653 14933 25656
rect 14967 25653 14979 25687
rect 14921 25647 14979 25653
rect 17589 25687 17647 25693
rect 17589 25653 17601 25687
rect 17635 25684 17647 25687
rect 17770 25684 17776 25696
rect 17635 25656 17776 25684
rect 17635 25653 17647 25656
rect 17589 25647 17647 25653
rect 17770 25644 17776 25656
rect 17828 25644 17834 25696
rect 18506 25644 18512 25696
rect 18564 25644 18570 25696
rect 18708 25684 18736 25783
rect 19150 25780 19156 25792
rect 19208 25780 19214 25832
rect 20717 25823 20775 25829
rect 20717 25789 20729 25823
rect 20763 25789 20775 25823
rect 20717 25783 20775 25789
rect 21085 25823 21143 25829
rect 21085 25789 21097 25823
rect 21131 25820 21143 25823
rect 21174 25820 21180 25832
rect 21131 25792 21180 25820
rect 21131 25789 21143 25792
rect 21085 25783 21143 25789
rect 18874 25712 18880 25764
rect 18932 25712 18938 25764
rect 18966 25712 18972 25764
rect 19024 25712 19030 25764
rect 20732 25752 20760 25783
rect 21174 25780 21180 25792
rect 21232 25780 21238 25832
rect 21266 25780 21272 25832
rect 21324 25780 21330 25832
rect 26142 25780 26148 25832
rect 26200 25820 26206 25832
rect 26344 25829 26372 25860
rect 26237 25823 26295 25829
rect 26237 25820 26249 25823
rect 26200 25792 26249 25820
rect 26200 25780 26206 25792
rect 26237 25789 26249 25792
rect 26283 25789 26295 25823
rect 26237 25783 26295 25789
rect 26329 25823 26387 25829
rect 26329 25789 26341 25823
rect 26375 25789 26387 25823
rect 26329 25783 26387 25789
rect 26510 25780 26516 25832
rect 26568 25820 26574 25832
rect 26605 25823 26663 25829
rect 26605 25820 26617 25823
rect 26568 25792 26617 25820
rect 26568 25780 26574 25792
rect 26605 25789 26617 25792
rect 26651 25789 26663 25823
rect 26605 25783 26663 25789
rect 26881 25823 26939 25829
rect 26881 25789 26893 25823
rect 26927 25789 26939 25823
rect 26881 25783 26939 25789
rect 27065 25823 27123 25829
rect 27065 25789 27077 25823
rect 27111 25820 27123 25823
rect 27154 25820 27160 25832
rect 27111 25792 27160 25820
rect 27111 25789 27123 25792
rect 27065 25783 27123 25789
rect 21450 25752 21456 25764
rect 20732 25724 21456 25752
rect 21450 25712 21456 25724
rect 21508 25712 21514 25764
rect 22554 25712 22560 25764
rect 22612 25712 22618 25764
rect 22848 25724 23244 25752
rect 19518 25684 19524 25696
rect 18708 25656 19524 25684
rect 19518 25644 19524 25656
rect 19576 25644 19582 25696
rect 19610 25644 19616 25696
rect 19668 25684 19674 25696
rect 20073 25687 20131 25693
rect 20073 25684 20085 25687
rect 19668 25656 20085 25684
rect 19668 25644 19674 25656
rect 20073 25653 20085 25656
rect 20119 25684 20131 25687
rect 20622 25684 20628 25696
rect 20119 25656 20628 25684
rect 20119 25653 20131 25656
rect 20073 25647 20131 25653
rect 20622 25644 20628 25656
rect 20680 25644 20686 25696
rect 20990 25644 20996 25696
rect 21048 25644 21054 25696
rect 22370 25644 22376 25696
rect 22428 25684 22434 25696
rect 22848 25684 22876 25724
rect 23216 25693 23244 25724
rect 25406 25712 25412 25764
rect 25464 25712 25470 25764
rect 26421 25755 26479 25761
rect 26421 25721 26433 25755
rect 26467 25721 26479 25755
rect 26896 25752 26924 25783
rect 26421 25715 26479 25721
rect 26620 25724 26924 25752
rect 22428 25656 22876 25684
rect 23201 25687 23259 25693
rect 22428 25644 22434 25656
rect 23201 25653 23213 25687
rect 23247 25653 23259 25687
rect 23201 25647 23259 25653
rect 26234 25644 26240 25696
rect 26292 25684 26298 25696
rect 26436 25684 26464 25715
rect 26620 25696 26648 25724
rect 26292 25656 26464 25684
rect 26292 25644 26298 25656
rect 26602 25644 26608 25696
rect 26660 25644 26666 25696
rect 26878 25644 26884 25696
rect 26936 25684 26942 25696
rect 27080 25684 27108 25783
rect 27154 25780 27160 25792
rect 27212 25780 27218 25832
rect 26936 25656 27108 25684
rect 27540 25684 27568 25860
rect 27617 25857 27629 25891
rect 27663 25888 27675 25891
rect 29012 25888 29040 25916
rect 29178 25888 29184 25900
rect 27663 25860 29184 25888
rect 27663 25857 27675 25860
rect 27617 25851 27675 25857
rect 29178 25848 29184 25860
rect 29236 25848 29242 25900
rect 29362 25848 29368 25900
rect 29420 25888 29426 25900
rect 29641 25891 29699 25897
rect 29641 25888 29653 25891
rect 29420 25860 29653 25888
rect 29420 25848 29426 25860
rect 29641 25857 29653 25860
rect 29687 25857 29699 25891
rect 29641 25851 29699 25857
rect 27893 25755 27951 25761
rect 27893 25721 27905 25755
rect 27939 25752 27951 25755
rect 28166 25752 28172 25764
rect 27939 25724 28172 25752
rect 27939 25721 27951 25724
rect 27893 25715 27951 25721
rect 28166 25712 28172 25724
rect 28224 25712 28230 25764
rect 29270 25752 29276 25764
rect 29118 25724 29276 25752
rect 29270 25712 29276 25724
rect 29328 25712 29334 25764
rect 30742 25752 30748 25764
rect 30392 25724 30748 25752
rect 30392 25684 30420 25724
rect 30742 25712 30748 25724
rect 30800 25712 30806 25764
rect 27540 25656 30420 25684
rect 30469 25687 30527 25693
rect 26936 25644 26942 25656
rect 30469 25653 30481 25687
rect 30515 25684 30527 25687
rect 30558 25684 30564 25696
rect 30515 25656 30564 25684
rect 30515 25653 30527 25656
rect 30469 25647 30527 25653
rect 30558 25644 30564 25656
rect 30616 25684 30622 25696
rect 32125 25687 32183 25693
rect 32125 25684 32137 25687
rect 30616 25656 32137 25684
rect 30616 25644 30622 25656
rect 32125 25653 32137 25656
rect 32171 25684 32183 25687
rect 32490 25684 32496 25696
rect 32171 25656 32496 25684
rect 32171 25653 32183 25656
rect 32125 25647 32183 25653
rect 32490 25644 32496 25656
rect 32548 25684 32554 25696
rect 33042 25684 33048 25696
rect 32548 25656 33048 25684
rect 32548 25644 32554 25656
rect 33042 25644 33048 25656
rect 33100 25644 33106 25696
rect 2760 25594 34316 25616
rect 2760 25542 7210 25594
rect 7262 25542 7274 25594
rect 7326 25542 7338 25594
rect 7390 25542 7402 25594
rect 7454 25542 7466 25594
rect 7518 25542 15099 25594
rect 15151 25542 15163 25594
rect 15215 25542 15227 25594
rect 15279 25542 15291 25594
rect 15343 25542 15355 25594
rect 15407 25542 22988 25594
rect 23040 25542 23052 25594
rect 23104 25542 23116 25594
rect 23168 25542 23180 25594
rect 23232 25542 23244 25594
rect 23296 25542 30877 25594
rect 30929 25542 30941 25594
rect 30993 25542 31005 25594
rect 31057 25542 31069 25594
rect 31121 25542 31133 25594
rect 31185 25542 34316 25594
rect 2760 25520 34316 25542
rect 3053 25483 3111 25489
rect 3053 25449 3065 25483
rect 3099 25480 3111 25483
rect 6089 25483 6147 25489
rect 3099 25452 4292 25480
rect 3099 25449 3111 25452
rect 3053 25443 3111 25449
rect 4264 25424 4292 25452
rect 6089 25449 6101 25483
rect 6135 25480 6147 25483
rect 6914 25480 6920 25492
rect 6135 25452 6920 25480
rect 6135 25449 6147 25452
rect 6089 25443 6147 25449
rect 6914 25440 6920 25452
rect 6972 25440 6978 25492
rect 9674 25440 9680 25492
rect 9732 25480 9738 25492
rect 10686 25480 10692 25492
rect 9732 25452 10692 25480
rect 9732 25440 9738 25452
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 11330 25440 11336 25492
rect 11388 25480 11394 25492
rect 12069 25483 12127 25489
rect 12069 25480 12081 25483
rect 11388 25452 12081 25480
rect 11388 25440 11394 25452
rect 12069 25449 12081 25452
rect 12115 25480 12127 25483
rect 12158 25480 12164 25492
rect 12115 25452 12164 25480
rect 12115 25449 12127 25452
rect 12069 25443 12127 25449
rect 12158 25440 12164 25452
rect 12216 25440 12222 25492
rect 13262 25440 13268 25492
rect 13320 25440 13326 25492
rect 13446 25440 13452 25492
rect 13504 25480 13510 25492
rect 14918 25480 14924 25492
rect 13504 25452 14924 25480
rect 13504 25440 13510 25452
rect 3878 25372 3884 25424
rect 3936 25372 3942 25424
rect 4246 25372 4252 25424
rect 4304 25372 4310 25424
rect 6178 25372 6184 25424
rect 6236 25412 6242 25424
rect 6365 25415 6423 25421
rect 6365 25412 6377 25415
rect 6236 25384 6377 25412
rect 6236 25372 6242 25384
rect 6365 25381 6377 25384
rect 6411 25381 6423 25415
rect 6365 25375 6423 25381
rect 6457 25415 6515 25421
rect 6457 25381 6469 25415
rect 6503 25412 6515 25415
rect 7377 25415 7435 25421
rect 7377 25412 7389 25415
rect 6503 25384 7389 25412
rect 6503 25381 6515 25384
rect 6457 25375 6515 25381
rect 7377 25381 7389 25384
rect 7423 25412 7435 25415
rect 8202 25412 8208 25424
rect 7423 25384 8208 25412
rect 7423 25381 7435 25384
rect 7377 25375 7435 25381
rect 8202 25372 8208 25384
rect 8260 25372 8266 25424
rect 8754 25372 8760 25424
rect 8812 25372 8818 25424
rect 11422 25372 11428 25424
rect 11480 25412 11486 25424
rect 12250 25412 12256 25424
rect 11480 25384 12256 25412
rect 11480 25372 11486 25384
rect 4798 25304 4804 25356
rect 4856 25304 4862 25356
rect 6273 25347 6331 25353
rect 6273 25313 6285 25347
rect 6319 25344 6331 25347
rect 6546 25344 6552 25356
rect 6319 25316 6552 25344
rect 6319 25313 6331 25316
rect 6273 25307 6331 25313
rect 6546 25304 6552 25316
rect 6604 25304 6610 25356
rect 6641 25347 6699 25353
rect 6641 25313 6653 25347
rect 6687 25344 6699 25347
rect 6687 25316 6868 25344
rect 6687 25313 6699 25316
rect 6641 25307 6699 25313
rect 4525 25279 4583 25285
rect 4525 25245 4537 25279
rect 4571 25276 4583 25279
rect 4893 25279 4951 25285
rect 4893 25276 4905 25279
rect 4571 25248 4905 25276
rect 4571 25245 4583 25248
rect 4525 25239 4583 25245
rect 4893 25245 4905 25248
rect 4939 25245 4951 25279
rect 4893 25239 4951 25245
rect 5537 25279 5595 25285
rect 5537 25245 5549 25279
rect 5583 25276 5595 25279
rect 5626 25276 5632 25288
rect 5583 25248 5632 25276
rect 5583 25245 5595 25248
rect 5537 25239 5595 25245
rect 5626 25236 5632 25248
rect 5684 25236 5690 25288
rect 6733 25279 6791 25285
rect 6733 25276 6745 25279
rect 6472 25248 6745 25276
rect 6472 25220 6500 25248
rect 6733 25245 6745 25248
rect 6779 25245 6791 25279
rect 6733 25239 6791 25245
rect 6454 25168 6460 25220
rect 6512 25168 6518 25220
rect 5902 25100 5908 25152
rect 5960 25140 5966 25152
rect 6840 25140 6868 25316
rect 8018 25304 8024 25356
rect 8076 25304 8082 25356
rect 11900 25353 11928 25384
rect 12250 25372 12256 25384
rect 12308 25372 12314 25424
rect 13280 25412 13308 25440
rect 13633 25415 13691 25421
rect 13633 25412 13645 25415
rect 13280 25384 13645 25412
rect 13633 25381 13645 25384
rect 13679 25381 13691 25415
rect 13633 25375 13691 25381
rect 11793 25347 11851 25353
rect 11793 25313 11805 25347
rect 11839 25313 11851 25347
rect 11793 25307 11851 25313
rect 11885 25347 11943 25353
rect 11885 25313 11897 25347
rect 11931 25313 11943 25347
rect 11885 25307 11943 25313
rect 8297 25279 8355 25285
rect 8297 25245 8309 25279
rect 8343 25276 8355 25279
rect 8846 25276 8852 25288
rect 8343 25248 8852 25276
rect 8343 25245 8355 25248
rect 8297 25239 8355 25245
rect 8846 25236 8852 25248
rect 8904 25236 8910 25288
rect 11808 25276 11836 25307
rect 12066 25304 12072 25356
rect 12124 25304 12130 25356
rect 13722 25304 13728 25356
rect 13780 25304 13786 25356
rect 13832 25353 13860 25452
rect 14918 25440 14924 25452
rect 14976 25480 14982 25492
rect 17678 25480 17684 25492
rect 14976 25452 17684 25480
rect 14976 25440 14982 25452
rect 17678 25440 17684 25452
rect 17736 25440 17742 25492
rect 19610 25440 19616 25492
rect 19668 25440 19674 25492
rect 19978 25480 19984 25492
rect 19720 25452 19984 25480
rect 14093 25415 14151 25421
rect 14093 25381 14105 25415
rect 14139 25412 14151 25415
rect 14182 25412 14188 25424
rect 14139 25384 14188 25412
rect 14139 25381 14151 25384
rect 14093 25375 14151 25381
rect 14182 25372 14188 25384
rect 14240 25372 14246 25424
rect 15749 25415 15807 25421
rect 15749 25412 15761 25415
rect 15318 25384 15761 25412
rect 15749 25381 15761 25384
rect 15795 25381 15807 25415
rect 15749 25375 15807 25381
rect 16390 25372 16396 25424
rect 16448 25372 16454 25424
rect 17402 25372 17408 25424
rect 17460 25372 17466 25424
rect 17696 25412 17724 25440
rect 19245 25415 19303 25421
rect 19245 25412 19257 25415
rect 17696 25384 18184 25412
rect 13817 25347 13875 25353
rect 13817 25313 13829 25347
rect 13863 25313 13875 25347
rect 13817 25307 13875 25313
rect 15841 25347 15899 25353
rect 15841 25313 15853 25347
rect 15887 25313 15899 25347
rect 15841 25307 15899 25313
rect 14458 25276 14464 25288
rect 11808 25248 14464 25276
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 15856 25220 15884 25307
rect 16408 25285 16436 25372
rect 18156 25353 18184 25384
rect 18800 25384 19257 25412
rect 18800 25353 18828 25384
rect 19245 25381 19257 25384
rect 19291 25381 19303 25415
rect 19245 25375 19303 25381
rect 19337 25415 19395 25421
rect 19337 25381 19349 25415
rect 19383 25412 19395 25415
rect 19628 25412 19656 25440
rect 19383 25384 19656 25412
rect 19383 25381 19395 25384
rect 19337 25375 19395 25381
rect 18141 25347 18199 25353
rect 18141 25313 18153 25347
rect 18187 25313 18199 25347
rect 18785 25347 18843 25353
rect 18785 25344 18797 25347
rect 18141 25307 18199 25313
rect 18616 25316 18797 25344
rect 18616 25288 18644 25316
rect 18785 25313 18797 25316
rect 18831 25313 18843 25347
rect 18785 25307 18843 25313
rect 19061 25347 19119 25353
rect 19061 25313 19073 25347
rect 19107 25313 19119 25347
rect 19061 25307 19119 25313
rect 16393 25279 16451 25285
rect 16393 25245 16405 25279
rect 16439 25245 16451 25279
rect 16393 25239 16451 25245
rect 16666 25236 16672 25288
rect 16724 25236 16730 25288
rect 17770 25236 17776 25288
rect 17828 25276 17834 25288
rect 17865 25279 17923 25285
rect 17865 25276 17877 25279
rect 17828 25248 17877 25276
rect 17828 25236 17834 25248
rect 17865 25245 17877 25248
rect 17911 25245 17923 25279
rect 17865 25239 17923 25245
rect 18598 25236 18604 25288
rect 18656 25236 18662 25288
rect 18690 25236 18696 25288
rect 18748 25276 18754 25288
rect 18969 25279 19027 25285
rect 18969 25276 18981 25279
rect 18748 25248 18981 25276
rect 18748 25236 18754 25248
rect 18969 25245 18981 25248
rect 19015 25245 19027 25279
rect 19076 25276 19104 25307
rect 19150 25304 19156 25356
rect 19208 25344 19214 25356
rect 19429 25347 19487 25353
rect 19429 25344 19441 25347
rect 19208 25316 19441 25344
rect 19208 25304 19214 25316
rect 19429 25313 19441 25316
rect 19475 25313 19487 25347
rect 19429 25307 19487 25313
rect 19518 25304 19524 25356
rect 19576 25304 19582 25356
rect 19720 25353 19748 25452
rect 19978 25440 19984 25452
rect 20036 25480 20042 25492
rect 21266 25480 21272 25492
rect 20036 25452 21272 25480
rect 20036 25440 20042 25452
rect 21266 25440 21272 25452
rect 21324 25440 21330 25492
rect 21450 25440 21456 25492
rect 21508 25440 21514 25492
rect 21545 25483 21603 25489
rect 21545 25449 21557 25483
rect 21591 25449 21603 25483
rect 21545 25443 21603 25449
rect 22005 25483 22063 25489
rect 22005 25449 22017 25483
rect 22051 25480 22063 25483
rect 22370 25480 22376 25492
rect 22051 25452 22376 25480
rect 22051 25449 22063 25452
rect 22005 25443 22063 25449
rect 20990 25372 20996 25424
rect 21048 25372 21054 25424
rect 21560 25412 21588 25443
rect 22370 25440 22376 25452
rect 22428 25440 22434 25492
rect 22465 25483 22523 25489
rect 22465 25449 22477 25483
rect 22511 25480 22523 25483
rect 22554 25480 22560 25492
rect 22511 25452 22560 25480
rect 22511 25449 22523 25452
rect 22465 25443 22523 25449
rect 22554 25440 22560 25452
rect 22612 25440 22618 25492
rect 23106 25480 23112 25492
rect 22664 25452 23112 25480
rect 22186 25412 22192 25424
rect 21560 25384 22192 25412
rect 22186 25372 22192 25384
rect 22244 25372 22250 25424
rect 19705 25347 19763 25353
rect 19705 25313 19717 25347
rect 19751 25313 19763 25347
rect 19705 25307 19763 25313
rect 21913 25347 21971 25353
rect 21913 25313 21925 25347
rect 21959 25313 21971 25347
rect 21913 25307 21971 25313
rect 22557 25347 22615 25353
rect 22557 25313 22569 25347
rect 22603 25344 22615 25347
rect 22664 25344 22692 25452
rect 23106 25440 23112 25452
rect 23164 25440 23170 25492
rect 24762 25480 24768 25492
rect 23492 25452 24768 25480
rect 23017 25415 23075 25421
rect 23017 25381 23029 25415
rect 23063 25412 23075 25415
rect 23382 25412 23388 25424
rect 23063 25384 23388 25412
rect 23063 25381 23075 25384
rect 23017 25375 23075 25381
rect 23382 25372 23388 25384
rect 23440 25372 23446 25424
rect 22603 25316 22692 25344
rect 22741 25347 22799 25353
rect 22603 25313 22615 25316
rect 22557 25307 22615 25313
rect 22741 25313 22753 25347
rect 22787 25313 22799 25347
rect 22741 25307 22799 25313
rect 19536 25276 19564 25304
rect 19076 25248 19564 25276
rect 19981 25279 20039 25285
rect 18969 25239 19027 25245
rect 19981 25245 19993 25279
rect 20027 25276 20039 25279
rect 20530 25276 20536 25288
rect 20027 25248 20536 25276
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 20622 25236 20628 25288
rect 20680 25276 20686 25288
rect 21928 25276 21956 25307
rect 20680 25248 21956 25276
rect 20680 25236 20686 25248
rect 22094 25236 22100 25288
rect 22152 25236 22158 25288
rect 11624 25180 12112 25208
rect 11624 25152 11652 25180
rect 5960 25112 6868 25140
rect 5960 25100 5966 25112
rect 6914 25100 6920 25152
rect 6972 25140 6978 25152
rect 7653 25143 7711 25149
rect 7653 25140 7665 25143
rect 6972 25112 7665 25140
rect 6972 25100 6978 25112
rect 7653 25109 7665 25112
rect 7699 25140 7711 25143
rect 7742 25140 7748 25152
rect 7699 25112 7748 25140
rect 7699 25109 7711 25112
rect 7653 25103 7711 25109
rect 7742 25100 7748 25112
rect 7800 25100 7806 25152
rect 9769 25143 9827 25149
rect 9769 25109 9781 25143
rect 9815 25140 9827 25143
rect 10410 25140 10416 25152
rect 9815 25112 10416 25140
rect 9815 25109 9827 25112
rect 9769 25103 9827 25109
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 11606 25100 11612 25152
rect 11664 25100 11670 25152
rect 12084 25140 12112 25180
rect 12250 25168 12256 25220
rect 12308 25208 12314 25220
rect 12434 25208 12440 25220
rect 12308 25180 12440 25208
rect 12308 25168 12314 25180
rect 12434 25168 12440 25180
rect 12492 25208 12498 25220
rect 13630 25208 13636 25220
rect 12492 25180 13636 25208
rect 12492 25168 12498 25180
rect 13630 25168 13636 25180
rect 13688 25168 13694 25220
rect 15562 25168 15568 25220
rect 15620 25168 15626 25220
rect 15838 25168 15844 25220
rect 15896 25208 15902 25220
rect 16574 25208 16580 25220
rect 15896 25180 16580 25208
rect 15896 25168 15902 25180
rect 16574 25168 16580 25180
rect 16632 25168 16638 25220
rect 16684 25140 16712 25236
rect 18506 25168 18512 25220
rect 18564 25208 18570 25220
rect 18564 25180 19748 25208
rect 18564 25168 18570 25180
rect 18616 25149 18644 25180
rect 12084 25112 16712 25140
rect 18601 25143 18659 25149
rect 18601 25109 18613 25143
rect 18647 25109 18659 25143
rect 18601 25103 18659 25109
rect 19610 25100 19616 25152
rect 19668 25100 19674 25152
rect 19720 25140 19748 25180
rect 22756 25140 22784 25307
rect 22922 25304 22928 25356
rect 22980 25304 22986 25356
rect 23109 25347 23167 25353
rect 23109 25313 23121 25347
rect 23155 25344 23167 25347
rect 23492 25344 23520 25452
rect 24762 25440 24768 25452
rect 24820 25440 24826 25492
rect 25225 25483 25283 25489
rect 25225 25449 25237 25483
rect 25271 25480 25283 25483
rect 25682 25480 25688 25492
rect 25271 25452 25688 25480
rect 25271 25449 25283 25452
rect 25225 25443 25283 25449
rect 25682 25440 25688 25452
rect 25740 25440 25746 25492
rect 25961 25483 26019 25489
rect 25961 25449 25973 25483
rect 26007 25480 26019 25483
rect 26970 25480 26976 25492
rect 26007 25452 26976 25480
rect 26007 25449 26019 25452
rect 25961 25443 26019 25449
rect 26970 25440 26976 25452
rect 27028 25440 27034 25492
rect 27338 25440 27344 25492
rect 27396 25480 27402 25492
rect 28902 25480 28908 25492
rect 27396 25452 28908 25480
rect 27396 25440 27402 25452
rect 28902 25440 28908 25452
rect 28960 25480 28966 25492
rect 29089 25483 29147 25489
rect 29089 25480 29101 25483
rect 28960 25452 29101 25480
rect 28960 25440 28966 25452
rect 29089 25449 29101 25452
rect 29135 25449 29147 25483
rect 29089 25443 29147 25449
rect 26436 25384 27752 25412
rect 23155 25316 23520 25344
rect 23155 25313 23167 25316
rect 23109 25307 23167 25313
rect 24854 25304 24860 25356
rect 24912 25304 24918 25356
rect 22940 25208 22968 25304
rect 23474 25236 23480 25288
rect 23532 25236 23538 25288
rect 23750 25236 23756 25288
rect 23808 25236 23814 25288
rect 25314 25236 25320 25288
rect 25372 25236 25378 25288
rect 26436 25285 26464 25384
rect 26605 25347 26663 25353
rect 26605 25313 26617 25347
rect 26651 25344 26663 25347
rect 27522 25344 27528 25356
rect 26651 25316 27528 25344
rect 26651 25313 26663 25316
rect 26605 25307 26663 25313
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 26421 25279 26479 25285
rect 26421 25245 26433 25279
rect 26467 25245 26479 25279
rect 26421 25239 26479 25245
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25276 26571 25279
rect 26694 25276 26700 25288
rect 26559 25248 26700 25276
rect 26559 25245 26571 25248
rect 26513 25239 26571 25245
rect 26694 25236 26700 25248
rect 26752 25236 26758 25288
rect 27062 25236 27068 25288
rect 27120 25236 27126 25288
rect 27617 25279 27675 25285
rect 27617 25245 27629 25279
rect 27663 25245 27675 25279
rect 27617 25239 27675 25245
rect 26973 25211 27031 25217
rect 22940 25180 23612 25208
rect 19720 25112 22784 25140
rect 23290 25100 23296 25152
rect 23348 25100 23354 25152
rect 23584 25140 23612 25180
rect 26973 25177 26985 25211
rect 27019 25208 27031 25211
rect 27632 25208 27660 25239
rect 27019 25180 27660 25208
rect 27724 25208 27752 25384
rect 28626 25304 28632 25356
rect 28684 25344 28690 25356
rect 28813 25347 28871 25353
rect 28813 25344 28825 25347
rect 28684 25316 28825 25344
rect 28684 25304 28690 25316
rect 28813 25313 28825 25316
rect 28859 25344 28871 25347
rect 30098 25344 30104 25356
rect 28859 25316 30104 25344
rect 28859 25313 28871 25316
rect 28813 25307 28871 25313
rect 30098 25304 30104 25316
rect 30156 25344 30162 25356
rect 30285 25347 30343 25353
rect 30285 25344 30297 25347
rect 30156 25316 30297 25344
rect 30156 25304 30162 25316
rect 30285 25313 30297 25316
rect 30331 25313 30343 25347
rect 30285 25307 30343 25313
rect 27798 25236 27804 25288
rect 27856 25236 27862 25288
rect 27890 25236 27896 25288
rect 27948 25276 27954 25288
rect 28721 25279 28779 25285
rect 28721 25276 28733 25279
rect 27948 25248 28733 25276
rect 27948 25236 27954 25248
rect 28721 25245 28733 25248
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 29822 25236 29828 25288
rect 29880 25236 29886 25288
rect 27724 25180 28488 25208
rect 27019 25177 27031 25180
rect 26973 25171 27031 25177
rect 28460 25152 28488 25180
rect 27706 25140 27712 25152
rect 23584 25112 27712 25140
rect 27706 25100 27712 25112
rect 27764 25100 27770 25152
rect 28442 25100 28448 25152
rect 28500 25100 28506 25152
rect 29273 25143 29331 25149
rect 29273 25109 29285 25143
rect 29319 25140 29331 25143
rect 29362 25140 29368 25152
rect 29319 25112 29368 25140
rect 29319 25109 29331 25112
rect 29273 25103 29331 25109
rect 29362 25100 29368 25112
rect 29420 25100 29426 25152
rect 30193 25143 30251 25149
rect 30193 25109 30205 25143
rect 30239 25140 30251 25143
rect 30558 25140 30564 25152
rect 30239 25112 30564 25140
rect 30239 25109 30251 25112
rect 30193 25103 30251 25109
rect 30558 25100 30564 25112
rect 30616 25100 30622 25152
rect 2760 25050 34316 25072
rect 2760 24998 6550 25050
rect 6602 24998 6614 25050
rect 6666 24998 6678 25050
rect 6730 24998 6742 25050
rect 6794 24998 6806 25050
rect 6858 24998 14439 25050
rect 14491 24998 14503 25050
rect 14555 24998 14567 25050
rect 14619 24998 14631 25050
rect 14683 24998 14695 25050
rect 14747 24998 22328 25050
rect 22380 24998 22392 25050
rect 22444 24998 22456 25050
rect 22508 24998 22520 25050
rect 22572 24998 22584 25050
rect 22636 24998 30217 25050
rect 30269 24998 30281 25050
rect 30333 24998 30345 25050
rect 30397 24998 30409 25050
rect 30461 24998 30473 25050
rect 30525 24998 34316 25050
rect 2760 24976 34316 24998
rect 4709 24939 4767 24945
rect 4709 24905 4721 24939
rect 4755 24936 4767 24939
rect 5626 24936 5632 24948
rect 4755 24908 5632 24936
rect 4755 24905 4767 24908
rect 4709 24899 4767 24905
rect 5626 24896 5632 24908
rect 5684 24896 5690 24948
rect 8573 24939 8631 24945
rect 8573 24905 8585 24939
rect 8619 24936 8631 24939
rect 8754 24936 8760 24948
rect 8619 24908 8760 24936
rect 8619 24905 8631 24908
rect 8573 24899 8631 24905
rect 8754 24896 8760 24908
rect 8812 24896 8818 24948
rect 8846 24896 8852 24948
rect 8904 24936 8910 24948
rect 9217 24939 9275 24945
rect 9217 24936 9229 24939
rect 8904 24908 9229 24936
rect 8904 24896 8910 24908
rect 9217 24905 9229 24908
rect 9263 24905 9275 24939
rect 9217 24899 9275 24905
rect 11422 24896 11428 24948
rect 11480 24896 11486 24948
rect 13722 24896 13728 24948
rect 13780 24936 13786 24948
rect 15838 24936 15844 24948
rect 13780 24908 15844 24936
rect 13780 24896 13786 24908
rect 15838 24896 15844 24908
rect 15896 24896 15902 24948
rect 18230 24896 18236 24948
rect 18288 24936 18294 24948
rect 18417 24939 18475 24945
rect 18417 24936 18429 24939
rect 18288 24908 18429 24936
rect 18288 24896 18294 24908
rect 18417 24905 18429 24908
rect 18463 24905 18475 24939
rect 18417 24899 18475 24905
rect 18598 24896 18604 24948
rect 18656 24896 18662 24948
rect 20530 24896 20536 24948
rect 20588 24896 20594 24948
rect 23474 24936 23480 24948
rect 22066 24908 23480 24936
rect 4172 24840 4936 24868
rect 4172 24809 4200 24840
rect 4908 24812 4936 24840
rect 6362 24828 6368 24880
rect 6420 24868 6426 24880
rect 6546 24868 6552 24880
rect 6420 24840 6552 24868
rect 6420 24828 6426 24840
rect 6546 24828 6552 24840
rect 6604 24828 6610 24880
rect 9876 24840 10640 24868
rect 4157 24803 4215 24809
rect 4157 24769 4169 24803
rect 4203 24769 4215 24803
rect 4157 24763 4215 24769
rect 4246 24760 4252 24812
rect 4304 24760 4310 24812
rect 4890 24760 4896 24812
rect 4948 24760 4954 24812
rect 5534 24760 5540 24812
rect 5592 24800 5598 24812
rect 6089 24803 6147 24809
rect 6089 24800 6101 24803
rect 5592 24772 6101 24800
rect 5592 24760 5598 24772
rect 6089 24769 6101 24772
rect 6135 24800 6147 24803
rect 7834 24800 7840 24812
rect 6135 24772 7840 24800
rect 6135 24769 6147 24772
rect 6089 24763 6147 24769
rect 7834 24760 7840 24772
rect 7892 24800 7898 24812
rect 9122 24800 9128 24812
rect 7892 24772 9128 24800
rect 7892 24760 7898 24772
rect 9122 24760 9128 24772
rect 9180 24760 9186 24812
rect 9876 24809 9904 24840
rect 10612 24812 10640 24840
rect 9861 24803 9919 24809
rect 9861 24769 9873 24803
rect 9907 24769 9919 24803
rect 9861 24763 9919 24769
rect 10060 24772 10548 24800
rect 1302 24692 1308 24744
rect 1360 24732 1366 24744
rect 3053 24735 3111 24741
rect 3053 24732 3065 24735
rect 1360 24704 3065 24732
rect 1360 24692 1366 24704
rect 3053 24701 3065 24704
rect 3099 24701 3111 24735
rect 3053 24695 3111 24701
rect 3329 24735 3387 24741
rect 3329 24701 3341 24735
rect 3375 24701 3387 24735
rect 3329 24695 3387 24701
rect 3344 24664 3372 24695
rect 4338 24692 4344 24744
rect 4396 24692 4402 24744
rect 6730 24732 6736 24744
rect 4632 24704 6736 24732
rect 4632 24664 4660 24704
rect 6730 24692 6736 24704
rect 6788 24692 6794 24744
rect 7650 24692 7656 24744
rect 7708 24732 7714 24744
rect 10060 24741 10088 24772
rect 10520 24744 10548 24772
rect 10594 24760 10600 24812
rect 10652 24760 10658 24812
rect 11440 24800 11468 24896
rect 21726 24828 21732 24880
rect 21784 24868 21790 24880
rect 22066 24868 22094 24908
rect 23474 24896 23480 24908
rect 23532 24896 23538 24948
rect 23750 24896 23756 24948
rect 23808 24936 23814 24948
rect 24213 24939 24271 24945
rect 24213 24936 24225 24939
rect 23808 24908 24225 24936
rect 23808 24896 23814 24908
rect 24213 24905 24225 24908
rect 24259 24905 24271 24939
rect 24213 24899 24271 24905
rect 25406 24896 25412 24948
rect 25464 24896 25470 24948
rect 26316 24939 26374 24945
rect 26316 24905 26328 24939
rect 26362 24936 26374 24939
rect 27062 24936 27068 24948
rect 26362 24908 27068 24936
rect 26362 24905 26374 24908
rect 26316 24899 26374 24905
rect 27062 24896 27068 24908
rect 27120 24896 27126 24948
rect 27798 24896 27804 24948
rect 27856 24896 27862 24948
rect 21784 24840 22094 24868
rect 21784 24828 21790 24840
rect 10980 24772 11468 24800
rect 8481 24735 8539 24741
rect 8481 24732 8493 24735
rect 7708 24704 8493 24732
rect 7708 24692 7714 24704
rect 8481 24701 8493 24704
rect 8527 24701 8539 24735
rect 8481 24695 8539 24701
rect 10045 24735 10103 24741
rect 10045 24701 10057 24735
rect 10091 24701 10103 24735
rect 10045 24695 10103 24701
rect 10226 24692 10232 24744
rect 10284 24692 10290 24744
rect 10502 24692 10508 24744
rect 10560 24692 10566 24744
rect 10980 24741 11008 24772
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24701 11023 24735
rect 10965 24695 11023 24701
rect 11057 24735 11115 24741
rect 11057 24701 11069 24735
rect 11103 24701 11115 24735
rect 11057 24695 11115 24701
rect 11149 24735 11207 24741
rect 11149 24701 11161 24735
rect 11195 24701 11207 24735
rect 11149 24695 11207 24701
rect 11241 24735 11299 24741
rect 11241 24701 11253 24735
rect 11287 24732 11299 24735
rect 11330 24732 11336 24744
rect 11287 24704 11336 24732
rect 11287 24701 11299 24704
rect 11241 24695 11299 24701
rect 7837 24667 7895 24673
rect 7837 24664 7849 24667
rect 3344 24636 4660 24664
rect 6196 24636 7849 24664
rect 6196 24608 6224 24636
rect 7837 24633 7849 24636
rect 7883 24633 7895 24667
rect 7837 24627 7895 24633
rect 9585 24667 9643 24673
rect 9585 24633 9597 24667
rect 9631 24664 9643 24667
rect 10137 24667 10195 24673
rect 10137 24664 10149 24667
rect 9631 24636 10149 24664
rect 9631 24633 9643 24636
rect 9585 24627 9643 24633
rect 10137 24633 10149 24636
rect 10183 24633 10195 24667
rect 10244 24664 10272 24692
rect 11072 24664 11100 24695
rect 10244 24636 11100 24664
rect 10137 24627 10195 24633
rect 4890 24556 4896 24608
rect 4948 24596 4954 24608
rect 4985 24599 5043 24605
rect 4985 24596 4997 24599
rect 4948 24568 4997 24596
rect 4948 24556 4954 24568
rect 4985 24565 4997 24568
rect 5031 24565 5043 24599
rect 4985 24559 5043 24565
rect 5442 24556 5448 24608
rect 5500 24596 5506 24608
rect 5626 24596 5632 24608
rect 5500 24568 5632 24596
rect 5500 24556 5506 24568
rect 5626 24556 5632 24568
rect 5684 24556 5690 24608
rect 6178 24556 6184 24608
rect 6236 24556 6242 24608
rect 6362 24556 6368 24608
rect 6420 24556 6426 24608
rect 6914 24556 6920 24608
rect 6972 24556 6978 24608
rect 7006 24556 7012 24608
rect 7064 24596 7070 24608
rect 7469 24599 7527 24605
rect 7469 24596 7481 24599
rect 7064 24568 7481 24596
rect 7064 24556 7070 24568
rect 7469 24565 7481 24568
rect 7515 24565 7527 24599
rect 7469 24559 7527 24565
rect 8570 24556 8576 24608
rect 8628 24596 8634 24608
rect 9677 24599 9735 24605
rect 9677 24596 9689 24599
rect 8628 24568 9689 24596
rect 8628 24556 8634 24568
rect 9677 24565 9689 24568
rect 9723 24596 9735 24599
rect 10781 24599 10839 24605
rect 10781 24596 10793 24599
rect 9723 24568 10793 24596
rect 9723 24565 9735 24568
rect 9677 24559 9735 24565
rect 10781 24565 10793 24568
rect 10827 24565 10839 24599
rect 11164 24596 11192 24695
rect 11330 24692 11336 24704
rect 11388 24692 11394 24744
rect 11440 24732 11468 24772
rect 13630 24760 13636 24812
rect 13688 24800 13694 24812
rect 15654 24800 15660 24812
rect 13688 24772 15660 24800
rect 13688 24760 13694 24772
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 16390 24760 16396 24812
rect 16448 24760 16454 24812
rect 16666 24760 16672 24812
rect 16724 24760 16730 24812
rect 16850 24809 16856 24812
rect 16807 24803 16856 24809
rect 16807 24769 16819 24803
rect 16853 24769 16856 24803
rect 16807 24763 16856 24769
rect 16850 24760 16856 24763
rect 16908 24760 16914 24812
rect 18049 24803 18107 24809
rect 18049 24769 18061 24803
rect 18095 24800 18107 24803
rect 18506 24800 18512 24812
rect 18095 24772 18512 24800
rect 18095 24769 18107 24772
rect 18049 24763 18107 24769
rect 18506 24760 18512 24772
rect 18564 24800 18570 24812
rect 19337 24803 19395 24809
rect 19337 24800 19349 24803
rect 18564 24772 19349 24800
rect 18564 24760 18570 24772
rect 19337 24769 19349 24772
rect 19383 24769 19395 24803
rect 19337 24763 19395 24769
rect 19610 24760 19616 24812
rect 19668 24800 19674 24812
rect 19889 24803 19947 24809
rect 19889 24800 19901 24803
rect 19668 24772 19901 24800
rect 19668 24760 19674 24772
rect 19889 24769 19901 24772
rect 19935 24769 19947 24803
rect 19889 24763 19947 24769
rect 20898 24760 20904 24812
rect 20956 24800 20962 24812
rect 21450 24800 21456 24812
rect 20956 24772 21456 24800
rect 20956 24760 20962 24772
rect 11514 24732 11520 24744
rect 11440 24704 11520 24732
rect 11514 24692 11520 24704
rect 11572 24732 11578 24744
rect 11609 24735 11667 24741
rect 11609 24732 11621 24735
rect 11572 24704 11621 24732
rect 11572 24692 11578 24704
rect 11609 24701 11621 24704
rect 11655 24701 11667 24735
rect 11609 24695 11667 24701
rect 11698 24692 11704 24744
rect 11756 24732 11762 24744
rect 11793 24735 11851 24741
rect 11793 24732 11805 24735
rect 11756 24704 11805 24732
rect 11756 24692 11762 24704
rect 11793 24701 11805 24704
rect 11839 24701 11851 24735
rect 11793 24695 11851 24701
rect 15746 24692 15752 24744
rect 15804 24692 15810 24744
rect 15933 24735 15991 24741
rect 15933 24701 15945 24735
rect 15979 24701 15991 24735
rect 15933 24695 15991 24701
rect 11422 24624 11428 24676
rect 11480 24624 11486 24676
rect 15948 24664 15976 24695
rect 16942 24692 16948 24744
rect 17000 24692 17006 24744
rect 18690 24732 18696 24744
rect 18340 24704 18696 24732
rect 15580 24636 15976 24664
rect 15580 24608 15608 24636
rect 18340 24608 18368 24704
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 18874 24692 18880 24744
rect 18932 24692 18938 24744
rect 19061 24735 19119 24741
rect 19061 24701 19073 24735
rect 19107 24732 19119 24735
rect 19426 24732 19432 24744
rect 19107 24704 19432 24732
rect 19107 24701 19119 24704
rect 19061 24695 19119 24701
rect 19426 24692 19432 24704
rect 19484 24692 19490 24744
rect 19702 24692 19708 24744
rect 19760 24692 19766 24744
rect 21008 24741 21036 24772
rect 21450 24760 21456 24772
rect 21508 24760 21514 24812
rect 22094 24760 22100 24812
rect 22152 24800 22158 24812
rect 22830 24800 22836 24812
rect 22152 24772 22836 24800
rect 22152 24760 22158 24772
rect 22830 24760 22836 24772
rect 22888 24760 22894 24812
rect 23290 24760 23296 24812
rect 23348 24800 23354 24812
rect 23569 24803 23627 24809
rect 23569 24800 23581 24803
rect 23348 24772 23581 24800
rect 23348 24760 23354 24772
rect 23569 24769 23581 24772
rect 23615 24769 23627 24803
rect 28626 24800 28632 24812
rect 23569 24763 23627 24769
rect 25884 24772 28632 24800
rect 20993 24735 21051 24741
rect 20993 24701 21005 24735
rect 21039 24701 21051 24735
rect 20993 24695 21051 24701
rect 21174 24692 21180 24744
rect 21232 24732 21238 24744
rect 21545 24735 21603 24741
rect 21545 24732 21557 24735
rect 21232 24704 21557 24732
rect 21232 24692 21238 24704
rect 21545 24701 21557 24704
rect 21591 24732 21603 24735
rect 23106 24732 23112 24744
rect 21591 24704 23112 24732
rect 21591 24701 21603 24704
rect 21545 24695 21603 24701
rect 23106 24692 23112 24704
rect 23164 24732 23170 24744
rect 24305 24735 24363 24741
rect 24305 24732 24317 24735
rect 23164 24704 24317 24732
rect 23164 24692 23170 24704
rect 18598 24624 18604 24676
rect 18656 24664 18662 24676
rect 18892 24664 18920 24692
rect 18656 24636 18920 24664
rect 19720 24664 19748 24692
rect 22922 24664 22928 24676
rect 19720 24636 20024 24664
rect 18656 24624 18662 24636
rect 12710 24596 12716 24608
rect 11164 24568 12716 24596
rect 10781 24559 10839 24565
rect 12710 24556 12716 24568
rect 12768 24556 12774 24608
rect 15562 24556 15568 24608
rect 15620 24556 15626 24608
rect 17586 24556 17592 24608
rect 17644 24556 17650 24608
rect 17957 24599 18015 24605
rect 17957 24565 17969 24599
rect 18003 24596 18015 24599
rect 18322 24596 18328 24608
rect 18003 24568 18328 24596
rect 18003 24565 18015 24568
rect 17957 24559 18015 24565
rect 18322 24556 18328 24568
rect 18380 24556 18386 24608
rect 18414 24556 18420 24608
rect 18472 24556 18478 24608
rect 19610 24556 19616 24608
rect 19668 24596 19674 24608
rect 19705 24599 19763 24605
rect 19705 24596 19717 24599
rect 19668 24568 19717 24596
rect 19668 24556 19674 24568
rect 19705 24565 19717 24568
rect 19751 24565 19763 24599
rect 19996 24596 20024 24636
rect 22066 24636 22928 24664
rect 22066 24596 22094 24636
rect 22922 24624 22928 24636
rect 22980 24664 22986 24676
rect 23201 24667 23259 24673
rect 23201 24664 23213 24667
rect 22980 24636 23213 24664
rect 22980 24624 22986 24636
rect 23201 24633 23213 24636
rect 23247 24633 23259 24667
rect 23201 24627 23259 24633
rect 23768 24608 23796 24704
rect 24305 24701 24317 24704
rect 24351 24701 24363 24735
rect 24305 24695 24363 24701
rect 24397 24735 24455 24741
rect 24397 24701 24409 24735
rect 24443 24732 24455 24735
rect 24854 24732 24860 24744
rect 24443 24704 24860 24732
rect 24443 24701 24455 24704
rect 24397 24695 24455 24701
rect 24320 24664 24348 24695
rect 24854 24692 24860 24704
rect 24912 24692 24918 24744
rect 25884 24741 25912 24772
rect 28626 24760 28632 24772
rect 28684 24760 28690 24812
rect 28994 24760 29000 24812
rect 29052 24760 29058 24812
rect 29273 24803 29331 24809
rect 29273 24769 29285 24803
rect 29319 24800 29331 24803
rect 29362 24800 29368 24812
rect 29319 24772 29368 24800
rect 29319 24769 29331 24772
rect 29273 24763 29331 24769
rect 29362 24760 29368 24772
rect 29420 24760 29426 24812
rect 25501 24735 25559 24741
rect 25501 24701 25513 24735
rect 25547 24701 25559 24735
rect 25501 24695 25559 24701
rect 25869 24735 25927 24741
rect 25869 24701 25881 24735
rect 25915 24701 25927 24735
rect 25869 24695 25927 24701
rect 26053 24735 26111 24741
rect 26053 24701 26065 24735
rect 26099 24701 26111 24735
rect 26053 24695 26111 24701
rect 25516 24664 25544 24695
rect 24320 24636 25544 24664
rect 25590 24624 25596 24676
rect 25648 24664 25654 24676
rect 26068 24664 26096 24695
rect 28810 24692 28816 24744
rect 28868 24692 28874 24744
rect 30558 24732 30564 24744
rect 30406 24704 30564 24732
rect 30558 24692 30564 24704
rect 30616 24692 30622 24744
rect 25648 24636 26096 24664
rect 26436 24636 26818 24664
rect 25648 24624 25654 24636
rect 19996 24568 22094 24596
rect 19705 24559 19763 24565
rect 22554 24556 22560 24608
rect 22612 24556 22618 24608
rect 23750 24556 23756 24608
rect 23808 24556 23814 24608
rect 25777 24599 25835 24605
rect 25777 24565 25789 24599
rect 25823 24596 25835 24599
rect 26436 24596 26464 24636
rect 27706 24624 27712 24676
rect 27764 24664 27770 24676
rect 28534 24664 28540 24676
rect 27764 24636 28540 24664
rect 27764 24624 27770 24636
rect 28534 24624 28540 24636
rect 28592 24624 28598 24676
rect 25823 24568 26464 24596
rect 25823 24565 25835 24568
rect 25777 24559 25835 24565
rect 27154 24556 27160 24608
rect 27212 24596 27218 24608
rect 27982 24596 27988 24608
rect 27212 24568 27988 24596
rect 27212 24556 27218 24568
rect 27982 24556 27988 24568
rect 28040 24556 28046 24608
rect 28258 24556 28264 24608
rect 28316 24556 28322 24608
rect 30558 24556 30564 24608
rect 30616 24596 30622 24608
rect 30745 24599 30803 24605
rect 30745 24596 30757 24599
rect 30616 24568 30757 24596
rect 30616 24556 30622 24568
rect 30745 24565 30757 24568
rect 30791 24565 30803 24599
rect 30745 24559 30803 24565
rect 2760 24506 34316 24528
rect 2760 24454 7210 24506
rect 7262 24454 7274 24506
rect 7326 24454 7338 24506
rect 7390 24454 7402 24506
rect 7454 24454 7466 24506
rect 7518 24454 15099 24506
rect 15151 24454 15163 24506
rect 15215 24454 15227 24506
rect 15279 24454 15291 24506
rect 15343 24454 15355 24506
rect 15407 24454 22988 24506
rect 23040 24454 23052 24506
rect 23104 24454 23116 24506
rect 23168 24454 23180 24506
rect 23232 24454 23244 24506
rect 23296 24454 30877 24506
rect 30929 24454 30941 24506
rect 30993 24454 31005 24506
rect 31057 24454 31069 24506
rect 31121 24454 31133 24506
rect 31185 24454 34316 24506
rect 2760 24432 34316 24454
rect 5813 24395 5871 24401
rect 5813 24361 5825 24395
rect 5859 24392 5871 24395
rect 6270 24392 6276 24404
rect 5859 24364 6276 24392
rect 5859 24361 5871 24364
rect 5813 24355 5871 24361
rect 6270 24352 6276 24364
rect 6328 24352 6334 24404
rect 6454 24352 6460 24404
rect 6512 24392 6518 24404
rect 6641 24395 6699 24401
rect 6641 24392 6653 24395
rect 6512 24364 6653 24392
rect 6512 24352 6518 24364
rect 6641 24361 6653 24364
rect 6687 24361 6699 24395
rect 6641 24355 6699 24361
rect 6730 24352 6736 24404
rect 6788 24392 6794 24404
rect 11054 24392 11060 24404
rect 6788 24364 11060 24392
rect 6788 24352 6794 24364
rect 11054 24352 11060 24364
rect 11112 24352 11118 24404
rect 12621 24395 12679 24401
rect 12621 24392 12633 24395
rect 11348 24364 12633 24392
rect 5074 24284 5080 24336
rect 5132 24284 5138 24336
rect 6825 24327 6883 24333
rect 6825 24293 6837 24327
rect 6871 24324 6883 24327
rect 7745 24327 7803 24333
rect 6871 24296 7604 24324
rect 6871 24293 6883 24296
rect 6825 24287 6883 24293
rect 5810 24216 5816 24268
rect 5868 24256 5874 24268
rect 6089 24259 6147 24265
rect 6089 24256 6101 24259
rect 5868 24228 6101 24256
rect 5868 24216 5874 24228
rect 6089 24225 6101 24228
rect 6135 24225 6147 24259
rect 6089 24219 6147 24225
rect 6178 24216 6184 24268
rect 6236 24216 6242 24268
rect 6457 24259 6515 24265
rect 6457 24225 6469 24259
rect 6503 24256 6515 24259
rect 6503 24228 6960 24256
rect 6503 24225 6515 24228
rect 6457 24219 6515 24225
rect 6932 24200 6960 24228
rect 4065 24191 4123 24197
rect 4065 24157 4077 24191
rect 4111 24157 4123 24191
rect 4065 24151 4123 24157
rect 4341 24191 4399 24197
rect 4341 24157 4353 24191
rect 4387 24188 4399 24191
rect 6549 24191 6607 24197
rect 4387 24160 5948 24188
rect 4387 24157 4399 24160
rect 4341 24151 4399 24157
rect 4080 24052 4108 24151
rect 5920 24129 5948 24160
rect 6549 24157 6561 24191
rect 6595 24157 6607 24191
rect 6549 24151 6607 24157
rect 5905 24123 5963 24129
rect 5905 24089 5917 24123
rect 5951 24089 5963 24123
rect 5905 24083 5963 24089
rect 6086 24080 6092 24132
rect 6144 24120 6150 24132
rect 6564 24120 6592 24151
rect 6914 24148 6920 24200
rect 6972 24148 6978 24200
rect 6144 24092 6592 24120
rect 7193 24123 7251 24129
rect 6144 24080 6150 24092
rect 7193 24089 7205 24123
rect 7239 24120 7251 24123
rect 7466 24120 7472 24132
rect 7239 24092 7472 24120
rect 7239 24089 7251 24092
rect 7193 24083 7251 24089
rect 7466 24080 7472 24092
rect 7524 24080 7530 24132
rect 4798 24052 4804 24064
rect 4080 24024 4804 24052
rect 4798 24012 4804 24024
rect 4856 24012 4862 24064
rect 6270 24012 6276 24064
rect 6328 24052 6334 24064
rect 6825 24055 6883 24061
rect 6825 24052 6837 24055
rect 6328 24024 6837 24052
rect 6328 24012 6334 24024
rect 6825 24021 6837 24024
rect 6871 24052 6883 24055
rect 7006 24052 7012 24064
rect 6871 24024 7012 24052
rect 6871 24021 6883 24024
rect 6825 24015 6883 24021
rect 7006 24012 7012 24024
rect 7064 24012 7070 24064
rect 7576 24061 7604 24296
rect 7745 24293 7757 24327
rect 7791 24324 7803 24327
rect 7791 24296 8786 24324
rect 7791 24293 7803 24296
rect 7745 24287 7803 24293
rect 9674 24284 9680 24336
rect 9732 24324 9738 24336
rect 11348 24324 11376 24364
rect 12621 24361 12633 24364
rect 12667 24392 12679 24395
rect 18141 24395 18199 24401
rect 12667 24364 15516 24392
rect 12667 24361 12679 24364
rect 12621 24355 12679 24361
rect 9732 24296 11376 24324
rect 9732 24284 9738 24296
rect 11422 24284 11428 24336
rect 11480 24284 11486 24336
rect 11882 24284 11888 24336
rect 11940 24284 11946 24336
rect 13446 24324 13452 24336
rect 13188 24296 13452 24324
rect 7653 24259 7711 24265
rect 7653 24225 7665 24259
rect 7699 24225 7711 24259
rect 7653 24219 7711 24225
rect 7660 24132 7688 24219
rect 10318 24216 10324 24268
rect 10376 24216 10382 24268
rect 10502 24216 10508 24268
rect 10560 24256 10566 24268
rect 10873 24259 10931 24265
rect 10873 24256 10885 24259
rect 10560 24228 10885 24256
rect 10560 24216 10566 24228
rect 10873 24225 10885 24228
rect 10919 24256 10931 24259
rect 11440 24256 11468 24284
rect 10919 24228 11468 24256
rect 10919 24225 10931 24228
rect 10873 24219 10931 24225
rect 11514 24216 11520 24268
rect 11572 24265 11578 24268
rect 13188 24265 13216 24296
rect 13446 24284 13452 24296
rect 13504 24284 13510 24336
rect 13998 24284 14004 24336
rect 14056 24284 14062 24336
rect 11572 24259 11604 24265
rect 11592 24225 11604 24259
rect 11572 24219 11604 24225
rect 12529 24259 12587 24265
rect 12529 24225 12541 24259
rect 12575 24256 12587 24259
rect 13173 24259 13231 24265
rect 12575 24228 13124 24256
rect 12575 24225 12587 24228
rect 12529 24219 12587 24225
rect 11572 24216 11578 24219
rect 8018 24148 8024 24200
rect 8076 24148 8082 24200
rect 8294 24148 8300 24200
rect 8352 24148 8358 24200
rect 11057 24191 11115 24197
rect 11057 24157 11069 24191
rect 11103 24188 11115 24191
rect 12342 24188 12348 24200
rect 11103 24160 12348 24188
rect 11103 24157 11115 24160
rect 11057 24151 11115 24157
rect 12342 24148 12348 24160
rect 12400 24148 12406 24200
rect 7650 24080 7656 24132
rect 7708 24080 7714 24132
rect 11241 24123 11299 24129
rect 11241 24089 11253 24123
rect 11287 24120 11299 24123
rect 11287 24092 12204 24120
rect 11287 24089 11299 24092
rect 11241 24083 11299 24089
rect 12176 24064 12204 24092
rect 7561 24055 7619 24061
rect 7561 24021 7573 24055
rect 7607 24052 7619 24055
rect 8478 24052 8484 24064
rect 7607 24024 8484 24052
rect 7607 24021 7619 24024
rect 7561 24015 7619 24021
rect 8478 24012 8484 24024
rect 8536 24012 8542 24064
rect 9769 24055 9827 24061
rect 9769 24021 9781 24055
rect 9815 24052 9827 24055
rect 10870 24052 10876 24064
rect 9815 24024 10876 24052
rect 9815 24021 9827 24024
rect 9769 24015 9827 24021
rect 10870 24012 10876 24024
rect 10928 24012 10934 24064
rect 11606 24012 11612 24064
rect 11664 24012 11670 24064
rect 11698 24012 11704 24064
rect 11756 24061 11762 24064
rect 11756 24055 11778 24061
rect 11766 24021 11778 24055
rect 11756 24015 11778 24021
rect 11756 24012 11762 24015
rect 12158 24012 12164 24064
rect 12216 24012 12222 24064
rect 13096 24052 13124 24228
rect 13173 24225 13185 24259
rect 13219 24225 13231 24259
rect 13173 24219 13231 24225
rect 14458 24216 14464 24268
rect 14516 24216 14522 24268
rect 15488 24265 15516 24364
rect 18141 24361 18153 24395
rect 18187 24392 18199 24395
rect 18598 24392 18604 24404
rect 18187 24364 18604 24392
rect 18187 24361 18199 24364
rect 18141 24355 18199 24361
rect 18598 24352 18604 24364
rect 18656 24352 18662 24404
rect 22002 24352 22008 24404
rect 22060 24392 22066 24404
rect 22094 24392 22100 24404
rect 22060 24364 22100 24392
rect 22060 24352 22066 24364
rect 22094 24352 22100 24364
rect 22152 24352 22158 24404
rect 28258 24392 28264 24404
rect 28177 24364 28264 24392
rect 17310 24284 17316 24336
rect 17368 24324 17374 24336
rect 17957 24327 18015 24333
rect 17957 24324 17969 24327
rect 17368 24296 17969 24324
rect 17368 24284 17374 24296
rect 17957 24293 17969 24296
rect 18003 24293 18015 24327
rect 17957 24287 18015 24293
rect 20625 24327 20683 24333
rect 20625 24293 20637 24327
rect 20671 24324 20683 24327
rect 22554 24324 22560 24336
rect 20671 24296 22560 24324
rect 20671 24293 20683 24296
rect 20625 24287 20683 24293
rect 22554 24284 22560 24296
rect 22612 24324 22618 24336
rect 23382 24324 23388 24336
rect 22612 24296 23388 24324
rect 22612 24284 22618 24296
rect 23382 24284 23388 24296
rect 23440 24284 23446 24336
rect 26234 24324 26240 24336
rect 23492 24296 26240 24324
rect 15473 24259 15531 24265
rect 15473 24225 15485 24259
rect 15519 24225 15531 24259
rect 19337 24259 19395 24265
rect 19337 24256 19349 24259
rect 15473 24219 15531 24225
rect 16960 24228 19349 24256
rect 13446 24148 13452 24200
rect 13504 24148 13510 24200
rect 14476 24188 14504 24216
rect 16960 24200 16988 24228
rect 19337 24225 19349 24228
rect 19383 24225 19395 24259
rect 19337 24219 19395 24225
rect 19518 24216 19524 24268
rect 19576 24256 19582 24268
rect 23492 24256 23520 24296
rect 26234 24284 26240 24296
rect 26292 24284 26298 24336
rect 27890 24324 27896 24336
rect 27738 24296 27896 24324
rect 27890 24284 27896 24296
rect 27948 24284 27954 24336
rect 28177 24333 28205 24364
rect 28258 24352 28264 24364
rect 28316 24352 28322 24404
rect 29365 24395 29423 24401
rect 29365 24361 29377 24395
rect 29411 24392 29423 24395
rect 29822 24392 29828 24404
rect 29411 24364 29828 24392
rect 29411 24361 29423 24364
rect 29365 24355 29423 24361
rect 29822 24352 29828 24364
rect 29880 24352 29886 24404
rect 28169 24327 28227 24333
rect 28169 24293 28181 24327
rect 28215 24293 28227 24327
rect 28169 24287 28227 24293
rect 28718 24284 28724 24336
rect 28776 24324 28782 24336
rect 28776 24296 31754 24324
rect 28776 24284 28782 24296
rect 19576 24228 23520 24256
rect 23661 24259 23719 24265
rect 19576 24216 19582 24228
rect 23661 24225 23673 24259
rect 23707 24225 23719 24259
rect 23661 24219 23719 24225
rect 14921 24191 14979 24197
rect 14921 24188 14933 24191
rect 14476 24160 14933 24188
rect 14476 24052 14504 24160
rect 14921 24157 14933 24160
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 15381 24191 15439 24197
rect 15381 24157 15393 24191
rect 15427 24188 15439 24191
rect 15654 24188 15660 24200
rect 15427 24160 15660 24188
rect 15427 24157 15439 24160
rect 15381 24151 15439 24157
rect 15654 24148 15660 24160
rect 15712 24148 15718 24200
rect 16942 24148 16948 24200
rect 17000 24148 17006 24200
rect 18230 24188 18236 24200
rect 17972 24160 18236 24188
rect 17586 24080 17592 24132
rect 17644 24080 17650 24132
rect 17972 24061 18000 24160
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 22646 24148 22652 24200
rect 22704 24188 22710 24200
rect 23017 24191 23075 24197
rect 23017 24188 23029 24191
rect 22704 24160 23029 24188
rect 22704 24148 22710 24160
rect 23017 24157 23029 24160
rect 23063 24157 23075 24191
rect 23676 24188 23704 24219
rect 28534 24216 28540 24268
rect 28592 24256 28598 24268
rect 28629 24259 28687 24265
rect 28629 24256 28641 24259
rect 28592 24228 28641 24256
rect 28592 24216 28598 24228
rect 28629 24225 28641 24228
rect 28675 24225 28687 24259
rect 28629 24219 28687 24225
rect 29546 24216 29552 24268
rect 29604 24216 29610 24268
rect 29638 24216 29644 24268
rect 29696 24216 29702 24268
rect 29733 24259 29791 24265
rect 29733 24225 29745 24259
rect 29779 24225 29791 24259
rect 29733 24219 29791 24225
rect 23750 24188 23756 24200
rect 23676 24160 23756 24188
rect 23017 24151 23075 24157
rect 23750 24148 23756 24160
rect 23808 24148 23814 24200
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24188 26755 24191
rect 27706 24188 27712 24200
rect 26743 24160 27712 24188
rect 26743 24157 26755 24160
rect 26697 24151 26755 24157
rect 27706 24148 27712 24160
rect 27764 24148 27770 24200
rect 28445 24191 28503 24197
rect 28445 24157 28457 24191
rect 28491 24188 28503 24191
rect 29178 24188 29184 24200
rect 28491 24160 29184 24188
rect 28491 24157 28503 24160
rect 28445 24151 28503 24157
rect 29178 24148 29184 24160
rect 29236 24148 29242 24200
rect 18414 24120 18420 24132
rect 18064 24092 18420 24120
rect 18064 24064 18092 24092
rect 18414 24080 18420 24092
rect 18472 24120 18478 24132
rect 18877 24123 18935 24129
rect 18877 24120 18889 24123
rect 18472 24092 18889 24120
rect 18472 24080 18478 24092
rect 18877 24089 18889 24092
rect 18923 24089 18935 24123
rect 27154 24120 27160 24132
rect 18877 24083 18935 24089
rect 19904 24092 27160 24120
rect 19904 24064 19932 24092
rect 27154 24080 27160 24092
rect 27212 24080 27218 24132
rect 29748 24120 29776 24219
rect 29822 24216 29828 24268
rect 29880 24265 29886 24268
rect 29880 24259 29929 24265
rect 29880 24225 29883 24259
rect 29917 24225 29929 24259
rect 29880 24219 29929 24225
rect 29880 24216 29886 24219
rect 30558 24216 30564 24268
rect 30616 24256 30622 24268
rect 30837 24259 30895 24265
rect 30837 24256 30849 24259
rect 30616 24228 30849 24256
rect 30616 24216 30622 24228
rect 30837 24225 30849 24228
rect 30883 24225 30895 24259
rect 30837 24219 30895 24225
rect 30009 24191 30067 24197
rect 30009 24188 30021 24191
rect 28644 24092 29776 24120
rect 29932 24160 30021 24188
rect 13096 24024 14504 24052
rect 17129 24055 17187 24061
rect 17129 24021 17141 24055
rect 17175 24052 17187 24055
rect 17497 24055 17555 24061
rect 17497 24052 17509 24055
rect 17175 24024 17509 24052
rect 17175 24021 17187 24024
rect 17129 24015 17187 24021
rect 17497 24021 17509 24024
rect 17543 24052 17555 24055
rect 17957 24055 18015 24061
rect 17957 24052 17969 24055
rect 17543 24024 17969 24052
rect 17543 24021 17555 24024
rect 17497 24015 17555 24021
rect 17957 24021 17969 24024
rect 18003 24021 18015 24055
rect 17957 24015 18015 24021
rect 18046 24012 18052 24064
rect 18104 24012 18110 24064
rect 18322 24012 18328 24064
rect 18380 24052 18386 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 18380 24024 18613 24052
rect 18380 24012 18386 24024
rect 18601 24021 18613 24024
rect 18647 24052 18659 24055
rect 18966 24052 18972 24064
rect 18647 24024 18972 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 18966 24012 18972 24024
rect 19024 24012 19030 24064
rect 19886 24012 19892 24064
rect 19944 24012 19950 24064
rect 21726 24012 21732 24064
rect 21784 24052 21790 24064
rect 21913 24055 21971 24061
rect 21913 24052 21925 24055
rect 21784 24024 21925 24052
rect 21784 24012 21790 24024
rect 21913 24021 21925 24024
rect 21959 24021 21971 24055
rect 21913 24015 21971 24021
rect 22186 24012 22192 24064
rect 22244 24052 22250 24064
rect 22465 24055 22523 24061
rect 22465 24052 22477 24055
rect 22244 24024 22477 24052
rect 22244 24012 22250 24024
rect 22465 24021 22477 24024
rect 22511 24021 22523 24055
rect 22465 24015 22523 24021
rect 23566 24012 23572 24064
rect 23624 24012 23630 24064
rect 26602 24012 26608 24064
rect 26660 24012 26666 24064
rect 27614 24012 27620 24064
rect 27672 24052 27678 24064
rect 28644 24052 28672 24092
rect 29932 24064 29960 24160
rect 30009 24157 30021 24160
rect 30055 24188 30067 24191
rect 30653 24191 30711 24197
rect 30653 24188 30665 24191
rect 30055 24160 30665 24188
rect 30055 24157 30067 24160
rect 30009 24151 30067 24157
rect 30653 24157 30665 24160
rect 30699 24157 30711 24191
rect 30653 24151 30711 24157
rect 31726 24120 31754 24296
rect 32217 24259 32275 24265
rect 32217 24225 32229 24259
rect 32263 24225 32275 24259
rect 32217 24219 32275 24225
rect 32232 24120 32260 24219
rect 33413 24191 33471 24197
rect 33413 24157 33425 24191
rect 33459 24188 33471 24191
rect 34698 24188 34704 24200
rect 33459 24160 34704 24188
rect 33459 24157 33471 24160
rect 33413 24151 33471 24157
rect 34698 24148 34704 24160
rect 34756 24148 34762 24200
rect 31726 24092 32260 24120
rect 27672 24024 28672 24052
rect 27672 24012 27678 24024
rect 28718 24012 28724 24064
rect 28776 24052 28782 24064
rect 28813 24055 28871 24061
rect 28813 24052 28825 24055
rect 28776 24024 28825 24052
rect 28776 24012 28782 24024
rect 28813 24021 28825 24024
rect 28859 24021 28871 24055
rect 28813 24015 28871 24021
rect 29914 24012 29920 24064
rect 29972 24012 29978 24064
rect 2760 23962 34316 23984
rect 2760 23910 6550 23962
rect 6602 23910 6614 23962
rect 6666 23910 6678 23962
rect 6730 23910 6742 23962
rect 6794 23910 6806 23962
rect 6858 23910 14439 23962
rect 14491 23910 14503 23962
rect 14555 23910 14567 23962
rect 14619 23910 14631 23962
rect 14683 23910 14695 23962
rect 14747 23910 22328 23962
rect 22380 23910 22392 23962
rect 22444 23910 22456 23962
rect 22508 23910 22520 23962
rect 22572 23910 22584 23962
rect 22636 23910 30217 23962
rect 30269 23910 30281 23962
rect 30333 23910 30345 23962
rect 30397 23910 30409 23962
rect 30461 23910 30473 23962
rect 30525 23910 34316 23962
rect 2760 23888 34316 23910
rect 5074 23808 5080 23860
rect 5132 23848 5138 23860
rect 5169 23851 5227 23857
rect 5169 23848 5181 23851
rect 5132 23820 5181 23848
rect 5132 23808 5138 23820
rect 5169 23817 5181 23820
rect 5215 23817 5227 23851
rect 5169 23811 5227 23817
rect 5994 23808 6000 23860
rect 6052 23848 6058 23860
rect 6089 23851 6147 23857
rect 6089 23848 6101 23851
rect 6052 23820 6101 23848
rect 6052 23808 6058 23820
rect 6089 23817 6101 23820
rect 6135 23848 6147 23851
rect 6270 23848 6276 23860
rect 6135 23820 6276 23848
rect 6135 23817 6147 23820
rect 6089 23811 6147 23817
rect 6270 23808 6276 23820
rect 6328 23808 6334 23860
rect 6454 23808 6460 23860
rect 6512 23848 6518 23860
rect 6733 23851 6791 23857
rect 6733 23848 6745 23851
rect 6512 23820 6745 23848
rect 6512 23808 6518 23820
rect 6733 23817 6745 23820
rect 6779 23848 6791 23851
rect 6822 23848 6828 23860
rect 6779 23820 6828 23848
rect 6779 23817 6791 23820
rect 6733 23811 6791 23817
rect 6822 23808 6828 23820
rect 6880 23808 6886 23860
rect 8205 23851 8263 23857
rect 8205 23817 8217 23851
rect 8251 23848 8263 23851
rect 8294 23848 8300 23860
rect 8251 23820 8300 23848
rect 8251 23817 8263 23820
rect 8205 23811 8263 23817
rect 8294 23808 8300 23820
rect 8352 23808 8358 23860
rect 9950 23808 9956 23860
rect 10008 23808 10014 23860
rect 10318 23808 10324 23860
rect 10376 23808 10382 23860
rect 11054 23808 11060 23860
rect 11112 23848 11118 23860
rect 11606 23848 11612 23860
rect 11112 23820 11612 23848
rect 11112 23808 11118 23820
rect 11606 23808 11612 23820
rect 11664 23808 11670 23860
rect 12897 23851 12955 23857
rect 12897 23817 12909 23851
rect 12943 23848 12955 23851
rect 13446 23848 13452 23860
rect 12943 23820 13452 23848
rect 12943 23817 12955 23820
rect 12897 23811 12955 23817
rect 13446 23808 13452 23820
rect 13504 23808 13510 23860
rect 13722 23808 13728 23860
rect 13780 23808 13786 23860
rect 13998 23808 14004 23860
rect 14056 23808 14062 23860
rect 15746 23808 15752 23860
rect 15804 23848 15810 23860
rect 15804 23820 25360 23848
rect 15804 23808 15810 23820
rect 6472 23780 6500 23808
rect 10226 23780 10232 23792
rect 5736 23752 6500 23780
rect 7944 23752 10232 23780
rect 3510 23672 3516 23724
rect 3568 23672 3574 23724
rect 4982 23672 4988 23724
rect 5040 23712 5046 23724
rect 5736 23721 5764 23752
rect 5721 23715 5779 23721
rect 5040 23684 5120 23712
rect 5040 23672 5046 23684
rect 3050 23604 3056 23656
rect 3108 23604 3114 23656
rect 5092 23653 5120 23684
rect 5721 23681 5733 23715
rect 5767 23681 5779 23715
rect 5721 23675 5779 23681
rect 5902 23672 5908 23724
rect 5960 23712 5966 23724
rect 6089 23715 6147 23721
rect 6089 23712 6101 23715
rect 5960 23684 6101 23712
rect 5960 23672 5966 23684
rect 6089 23681 6101 23684
rect 6135 23712 6147 23715
rect 6362 23712 6368 23724
rect 6135 23684 6368 23712
rect 6135 23681 6147 23684
rect 6089 23675 6147 23681
rect 6362 23672 6368 23684
rect 6420 23672 6426 23724
rect 7944 23721 7972 23752
rect 10226 23740 10232 23752
rect 10284 23740 10290 23792
rect 11146 23740 11152 23792
rect 11204 23780 11210 23792
rect 11425 23783 11483 23789
rect 11425 23780 11437 23783
rect 11204 23752 11437 23780
rect 11204 23740 11210 23752
rect 11425 23749 11437 23752
rect 11471 23749 11483 23783
rect 11425 23743 11483 23749
rect 7929 23715 7987 23721
rect 7929 23681 7941 23715
rect 7975 23681 7987 23715
rect 7929 23675 7987 23681
rect 8021 23715 8079 23721
rect 8021 23681 8033 23715
rect 8067 23712 8079 23715
rect 8570 23712 8576 23724
rect 8067 23684 8576 23712
rect 8067 23681 8079 23684
rect 8021 23675 8079 23681
rect 5077 23647 5135 23653
rect 5077 23613 5089 23647
rect 5123 23613 5135 23647
rect 5077 23607 5135 23613
rect 6917 23647 6975 23653
rect 6917 23613 6929 23647
rect 6963 23644 6975 23647
rect 7650 23644 7656 23656
rect 6963 23616 7656 23644
rect 6963 23613 6975 23616
rect 6917 23607 6975 23613
rect 5092 23576 5120 23607
rect 6932 23576 6960 23607
rect 7650 23604 7656 23616
rect 7708 23604 7714 23656
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 8036 23644 8064 23675
rect 8570 23672 8576 23684
rect 8628 23672 8634 23724
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23712 9827 23715
rect 10502 23712 10508 23724
rect 9815 23684 10508 23712
rect 9815 23681 9827 23684
rect 9769 23675 9827 23681
rect 10502 23672 10508 23684
rect 10560 23672 10566 23724
rect 12434 23712 12440 23724
rect 11624 23684 12440 23712
rect 7892 23616 8064 23644
rect 7892 23604 7898 23616
rect 8294 23604 8300 23656
rect 8352 23604 8358 23656
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23644 8999 23647
rect 9033 23647 9091 23653
rect 9033 23644 9045 23647
rect 8987 23616 9045 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 9033 23613 9045 23616
rect 9079 23613 9091 23647
rect 9033 23607 9091 23613
rect 9214 23604 9220 23656
rect 9272 23644 9278 23656
rect 9585 23647 9643 23653
rect 9585 23644 9597 23647
rect 9272 23616 9597 23644
rect 9272 23604 9278 23616
rect 9585 23613 9597 23616
rect 9631 23613 9643 23647
rect 9585 23607 9643 23613
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 10042 23644 10048 23656
rect 9916 23616 10048 23644
rect 9916 23604 9922 23616
rect 10042 23604 10048 23616
rect 10100 23604 10106 23656
rect 10229 23647 10287 23653
rect 10229 23644 10241 23647
rect 10152 23616 10241 23644
rect 10152 23588 10180 23616
rect 10229 23613 10241 23616
rect 10275 23613 10287 23647
rect 10229 23607 10287 23613
rect 10410 23604 10416 23656
rect 10468 23644 10474 23656
rect 11624 23653 11652 23684
rect 12434 23672 12440 23684
rect 12492 23712 12498 23724
rect 12492 23684 12756 23712
rect 12492 23672 12498 23684
rect 10689 23647 10747 23653
rect 10689 23644 10701 23647
rect 10468 23616 10701 23644
rect 10468 23604 10474 23616
rect 10689 23613 10701 23616
rect 10735 23613 10747 23647
rect 10689 23607 10747 23613
rect 11609 23647 11667 23653
rect 11609 23613 11621 23647
rect 11655 23613 11667 23647
rect 11609 23607 11667 23613
rect 11698 23604 11704 23656
rect 11756 23604 11762 23656
rect 11790 23604 11796 23656
rect 11848 23644 11854 23656
rect 11885 23647 11943 23653
rect 11885 23644 11897 23647
rect 11848 23616 11897 23644
rect 11848 23604 11854 23616
rect 11885 23613 11897 23616
rect 11931 23613 11943 23647
rect 11885 23607 11943 23613
rect 11974 23604 11980 23656
rect 12032 23604 12038 23656
rect 12066 23604 12072 23656
rect 12124 23644 12130 23656
rect 12728 23653 12756 23684
rect 12345 23647 12403 23653
rect 12124 23616 12169 23644
rect 12124 23604 12130 23616
rect 12345 23613 12357 23647
rect 12391 23644 12403 23647
rect 12621 23647 12679 23653
rect 12621 23644 12633 23647
rect 12391 23616 12633 23644
rect 12391 23613 12403 23616
rect 12345 23607 12403 23613
rect 12621 23613 12633 23616
rect 12667 23613 12679 23647
rect 12621 23607 12679 23613
rect 12713 23647 12771 23653
rect 12713 23613 12725 23647
rect 12759 23613 12771 23647
rect 12713 23607 12771 23613
rect 13633 23647 13691 23653
rect 13633 23613 13645 23647
rect 13679 23644 13691 23647
rect 13740 23644 13768 23808
rect 16390 23740 16396 23792
rect 16448 23780 16454 23792
rect 18325 23783 18383 23789
rect 18325 23780 18337 23783
rect 16448 23752 18337 23780
rect 16448 23740 16454 23752
rect 18325 23749 18337 23752
rect 18371 23780 18383 23783
rect 18598 23780 18604 23792
rect 18371 23752 18604 23780
rect 18371 23749 18383 23752
rect 18325 23743 18383 23749
rect 18598 23740 18604 23752
rect 18656 23740 18662 23792
rect 19334 23740 19340 23792
rect 19392 23780 19398 23792
rect 19392 23752 20024 23780
rect 19392 23740 19398 23752
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23712 15623 23715
rect 18414 23712 18420 23724
rect 15611 23684 18420 23712
rect 15611 23681 15623 23684
rect 15565 23675 15623 23681
rect 18414 23672 18420 23684
rect 18472 23672 18478 23724
rect 19076 23684 19748 23712
rect 13909 23647 13967 23653
rect 13909 23644 13921 23647
rect 13679 23616 13921 23644
rect 13679 23613 13691 23616
rect 13633 23607 13691 23613
rect 13909 23613 13921 23616
rect 13955 23613 13967 23647
rect 13909 23607 13967 23613
rect 14826 23604 14832 23656
rect 14884 23604 14890 23656
rect 16393 23647 16451 23653
rect 16393 23613 16405 23647
rect 16439 23644 16451 23647
rect 16850 23644 16856 23656
rect 16439 23616 16856 23644
rect 16439 23613 16451 23616
rect 16393 23607 16451 23613
rect 16850 23604 16856 23616
rect 16908 23604 16914 23656
rect 19076 23653 19104 23684
rect 19061 23647 19119 23653
rect 19061 23613 19073 23647
rect 19107 23613 19119 23647
rect 19610 23644 19616 23656
rect 19061 23607 19119 23613
rect 19444 23616 19616 23644
rect 5092 23548 6960 23576
rect 7561 23579 7619 23585
rect 7561 23545 7573 23579
rect 7607 23576 7619 23579
rect 7607 23548 9444 23576
rect 7607 23545 7619 23548
rect 7561 23539 7619 23545
rect 5810 23468 5816 23520
rect 5868 23508 5874 23520
rect 5905 23511 5963 23517
rect 5905 23508 5917 23511
rect 5868 23480 5917 23508
rect 5868 23468 5874 23480
rect 5905 23477 5917 23480
rect 5951 23477 5963 23511
rect 5905 23471 5963 23477
rect 7006 23468 7012 23520
rect 7064 23468 7070 23520
rect 7466 23468 7472 23520
rect 7524 23508 7530 23520
rect 7650 23508 7656 23520
rect 7524 23480 7656 23508
rect 7524 23468 7530 23480
rect 7650 23468 7656 23480
rect 7708 23468 7714 23520
rect 8938 23468 8944 23520
rect 8996 23508 9002 23520
rect 9214 23508 9220 23520
rect 8996 23480 9220 23508
rect 8996 23468 9002 23480
rect 9214 23468 9220 23480
rect 9272 23468 9278 23520
rect 9416 23517 9444 23548
rect 10134 23536 10140 23588
rect 10192 23576 10198 23588
rect 11716 23576 11744 23604
rect 10192 23548 11744 23576
rect 10192 23536 10198 23548
rect 12894 23536 12900 23588
rect 12952 23536 12958 23588
rect 13725 23579 13783 23585
rect 13725 23545 13737 23579
rect 13771 23576 13783 23579
rect 13771 23548 14136 23576
rect 13771 23545 13783 23548
rect 13725 23539 13783 23545
rect 14108 23520 14136 23548
rect 15672 23548 17448 23576
rect 15672 23520 15700 23548
rect 9401 23511 9459 23517
rect 9401 23477 9413 23511
rect 9447 23477 9459 23511
rect 9401 23471 9459 23477
rect 10594 23468 10600 23520
rect 10652 23508 10658 23520
rect 10873 23511 10931 23517
rect 10873 23508 10885 23511
rect 10652 23480 10885 23508
rect 10652 23468 10658 23480
rect 10873 23477 10885 23480
rect 10919 23508 10931 23511
rect 11790 23508 11796 23520
rect 10919 23480 11796 23508
rect 10919 23477 10931 23480
rect 10873 23471 10931 23477
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 12342 23468 12348 23520
rect 12400 23508 12406 23520
rect 13814 23508 13820 23520
rect 12400 23480 13820 23508
rect 12400 23468 12406 23480
rect 13814 23468 13820 23480
rect 13872 23468 13878 23520
rect 14090 23468 14096 23520
rect 14148 23468 14154 23520
rect 14182 23468 14188 23520
rect 14240 23468 14246 23520
rect 14274 23468 14280 23520
rect 14332 23508 14338 23520
rect 14921 23511 14979 23517
rect 14921 23508 14933 23511
rect 14332 23480 14933 23508
rect 14332 23468 14338 23480
rect 14921 23477 14933 23480
rect 14967 23477 14979 23511
rect 14921 23471 14979 23477
rect 15654 23468 15660 23520
rect 15712 23468 15718 23520
rect 15746 23468 15752 23520
rect 15804 23468 15810 23520
rect 17310 23468 17316 23520
rect 17368 23468 17374 23520
rect 17420 23508 17448 23548
rect 17862 23536 17868 23588
rect 17920 23536 17926 23588
rect 17957 23511 18015 23517
rect 17957 23508 17969 23511
rect 17420 23480 17969 23508
rect 17957 23477 17969 23480
rect 18003 23508 18015 23511
rect 18046 23508 18052 23520
rect 18003 23480 18052 23508
rect 18003 23477 18015 23480
rect 17957 23471 18015 23477
rect 18046 23468 18052 23480
rect 18104 23468 18110 23520
rect 18969 23511 19027 23517
rect 18969 23477 18981 23511
rect 19015 23508 19027 23511
rect 19058 23508 19064 23520
rect 19015 23480 19064 23508
rect 19015 23477 19027 23480
rect 18969 23471 19027 23477
rect 19058 23468 19064 23480
rect 19116 23468 19122 23520
rect 19334 23468 19340 23520
rect 19392 23508 19398 23520
rect 19444 23517 19472 23616
rect 19610 23604 19616 23616
rect 19668 23604 19674 23656
rect 19429 23511 19487 23517
rect 19429 23508 19441 23511
rect 19392 23480 19441 23508
rect 19392 23468 19398 23480
rect 19429 23477 19441 23480
rect 19475 23477 19487 23511
rect 19720 23508 19748 23684
rect 19886 23604 19892 23656
rect 19944 23604 19950 23656
rect 19996 23653 20024 23752
rect 23566 23740 23572 23792
rect 23624 23740 23630 23792
rect 23658 23740 23664 23792
rect 23716 23740 23722 23792
rect 25332 23780 25360 23820
rect 25406 23808 25412 23860
rect 25464 23848 25470 23860
rect 28074 23848 28080 23860
rect 25464 23820 28080 23848
rect 25464 23808 25470 23820
rect 28074 23808 28080 23820
rect 28132 23808 28138 23860
rect 28261 23851 28319 23857
rect 28261 23817 28273 23851
rect 28307 23848 28319 23851
rect 28810 23848 28816 23860
rect 28307 23820 28816 23848
rect 28307 23817 28319 23820
rect 28261 23811 28319 23817
rect 28810 23808 28816 23820
rect 28868 23808 28874 23860
rect 28902 23808 28908 23860
rect 28960 23808 28966 23860
rect 29546 23808 29552 23860
rect 29604 23848 29610 23860
rect 29917 23851 29975 23857
rect 29917 23848 29929 23851
rect 29604 23820 29929 23848
rect 29604 23808 29610 23820
rect 29917 23817 29929 23820
rect 29963 23817 29975 23851
rect 29917 23811 29975 23817
rect 28920 23780 28948 23808
rect 25332 23752 28948 23780
rect 29638 23740 29644 23792
rect 29696 23780 29702 23792
rect 29733 23783 29791 23789
rect 29733 23780 29745 23783
rect 29696 23752 29745 23780
rect 29696 23740 29702 23752
rect 29733 23749 29745 23752
rect 29779 23749 29791 23783
rect 29733 23743 29791 23749
rect 22186 23672 22192 23724
rect 22244 23672 22250 23724
rect 19981 23647 20039 23653
rect 19981 23613 19993 23647
rect 20027 23644 20039 23647
rect 20530 23644 20536 23656
rect 20027 23616 20536 23644
rect 20027 23613 20039 23616
rect 19981 23607 20039 23613
rect 20530 23604 20536 23616
rect 20588 23604 20594 23656
rect 20993 23647 21051 23653
rect 20993 23613 21005 23647
rect 21039 23644 21051 23647
rect 21082 23644 21088 23656
rect 21039 23616 21088 23644
rect 21039 23613 21051 23616
rect 20993 23607 21051 23613
rect 19794 23536 19800 23588
rect 19852 23536 19858 23588
rect 21008 23576 21036 23607
rect 21082 23604 21088 23616
rect 21140 23604 21146 23656
rect 21726 23604 21732 23656
rect 21784 23644 21790 23656
rect 21913 23647 21971 23653
rect 21913 23644 21925 23647
rect 21784 23616 21925 23644
rect 21784 23604 21790 23616
rect 21913 23613 21925 23616
rect 21959 23613 21971 23647
rect 23584 23644 23612 23740
rect 24026 23672 24032 23724
rect 24084 23712 24090 23724
rect 25590 23712 25596 23724
rect 24084 23684 25596 23712
rect 24084 23672 24090 23684
rect 25590 23672 25596 23684
rect 25648 23672 25654 23724
rect 25777 23715 25835 23721
rect 25777 23681 25789 23715
rect 25823 23712 25835 23715
rect 27617 23715 27675 23721
rect 25823 23684 27476 23712
rect 25823 23681 25835 23684
rect 25777 23675 25835 23681
rect 27448 23656 27476 23684
rect 27617 23681 27629 23715
rect 27663 23712 27675 23715
rect 27663 23684 28396 23712
rect 27663 23681 27675 23684
rect 27617 23675 27675 23681
rect 28368 23656 28396 23684
rect 29564 23684 29868 23712
rect 23322 23616 23612 23644
rect 21913 23607 21971 23613
rect 26326 23604 26332 23656
rect 26384 23644 26390 23656
rect 26605 23647 26663 23653
rect 26605 23644 26617 23647
rect 26384 23616 26617 23644
rect 26384 23604 26390 23616
rect 26605 23613 26617 23616
rect 26651 23613 26663 23647
rect 26605 23607 26663 23613
rect 26694 23604 26700 23656
rect 26752 23604 26758 23656
rect 27430 23604 27436 23656
rect 27488 23604 27494 23656
rect 27706 23644 27712 23656
rect 27540 23616 27712 23644
rect 19904 23548 21036 23576
rect 24305 23579 24363 23585
rect 19904 23508 19932 23548
rect 24305 23545 24317 23579
rect 24351 23545 24363 23579
rect 24305 23539 24363 23545
rect 19720 23480 19932 23508
rect 19429 23471 19487 23477
rect 20162 23468 20168 23520
rect 20220 23468 20226 23520
rect 20990 23468 20996 23520
rect 21048 23508 21054 23520
rect 21085 23511 21143 23517
rect 21085 23508 21097 23511
rect 21048 23480 21097 23508
rect 21048 23468 21054 23480
rect 21085 23477 21097 23480
rect 21131 23477 21143 23511
rect 24320 23508 24348 23539
rect 25038 23536 25044 23588
rect 25096 23536 25102 23588
rect 26053 23579 26111 23585
rect 26053 23576 26065 23579
rect 25608 23548 26065 23576
rect 25608 23508 25636 23548
rect 26053 23545 26065 23548
rect 26099 23545 26111 23579
rect 26712 23576 26740 23604
rect 27540 23576 27568 23616
rect 27706 23604 27712 23616
rect 27764 23653 27770 23656
rect 27764 23647 27813 23653
rect 27764 23613 27767 23647
rect 27801 23613 27813 23647
rect 27764 23607 27813 23613
rect 27893 23647 27951 23653
rect 27893 23613 27905 23647
rect 27939 23613 27951 23647
rect 27893 23607 27951 23613
rect 27764 23604 27770 23607
rect 26712 23548 27568 23576
rect 26053 23539 26111 23545
rect 27614 23536 27620 23588
rect 27672 23536 27678 23588
rect 24320 23480 25636 23508
rect 27249 23511 27307 23517
rect 21085 23471 21143 23477
rect 27249 23477 27261 23511
rect 27295 23508 27307 23511
rect 27338 23508 27344 23520
rect 27295 23480 27344 23508
rect 27295 23477 27307 23480
rect 27249 23471 27307 23477
rect 27338 23468 27344 23480
rect 27396 23468 27402 23520
rect 27632 23508 27660 23536
rect 27908 23508 27936 23607
rect 28074 23604 28080 23656
rect 28132 23604 28138 23656
rect 28350 23604 28356 23656
rect 28408 23604 28414 23656
rect 28537 23647 28595 23653
rect 28537 23613 28549 23647
rect 28583 23613 28595 23647
rect 29564 23644 29592 23684
rect 29840 23653 29868 23684
rect 28537 23607 28595 23613
rect 28966 23616 29592 23644
rect 29641 23647 29699 23653
rect 27985 23579 28043 23585
rect 27985 23545 27997 23579
rect 28031 23576 28043 23579
rect 28445 23579 28503 23585
rect 28445 23576 28457 23579
rect 28031 23548 28457 23576
rect 28031 23545 28043 23548
rect 27985 23539 28043 23545
rect 28445 23545 28457 23548
rect 28491 23545 28503 23579
rect 28445 23539 28503 23545
rect 28552 23576 28580 23607
rect 28966 23576 28994 23616
rect 29641 23613 29653 23647
rect 29687 23613 29699 23647
rect 29641 23607 29699 23613
rect 29825 23647 29883 23653
rect 29825 23613 29837 23647
rect 29871 23644 29883 23647
rect 30285 23647 30343 23653
rect 30285 23644 30297 23647
rect 29871 23616 30297 23644
rect 29871 23613 29883 23616
rect 29825 23607 29883 23613
rect 30285 23613 30297 23616
rect 30331 23613 30343 23647
rect 30285 23607 30343 23613
rect 28552 23548 28994 23576
rect 29656 23576 29684 23607
rect 33778 23604 33784 23656
rect 33836 23604 33842 23656
rect 29914 23576 29920 23588
rect 29656 23548 29920 23576
rect 28552 23520 28580 23548
rect 29914 23536 29920 23548
rect 29972 23576 29978 23588
rect 30101 23579 30159 23585
rect 30101 23576 30113 23579
rect 29972 23548 30113 23576
rect 29972 23536 29978 23548
rect 30101 23545 30113 23548
rect 30147 23545 30159 23579
rect 30101 23539 30159 23545
rect 27632 23480 27936 23508
rect 28534 23468 28540 23520
rect 28592 23468 28598 23520
rect 28902 23468 28908 23520
rect 28960 23508 28966 23520
rect 33796 23508 33824 23604
rect 28960 23480 33824 23508
rect 28960 23468 28966 23480
rect 2760 23418 34316 23440
rect 2760 23366 7210 23418
rect 7262 23366 7274 23418
rect 7326 23366 7338 23418
rect 7390 23366 7402 23418
rect 7454 23366 7466 23418
rect 7518 23366 15099 23418
rect 15151 23366 15163 23418
rect 15215 23366 15227 23418
rect 15279 23366 15291 23418
rect 15343 23366 15355 23418
rect 15407 23366 22988 23418
rect 23040 23366 23052 23418
rect 23104 23366 23116 23418
rect 23168 23366 23180 23418
rect 23232 23366 23244 23418
rect 23296 23366 30877 23418
rect 30929 23366 30941 23418
rect 30993 23366 31005 23418
rect 31057 23366 31069 23418
rect 31121 23366 31133 23418
rect 31185 23366 34316 23418
rect 2760 23344 34316 23366
rect 7745 23307 7803 23313
rect 7745 23273 7757 23307
rect 7791 23304 7803 23307
rect 8294 23304 8300 23316
rect 7791 23276 8300 23304
rect 7791 23273 7803 23276
rect 7745 23267 7803 23273
rect 8294 23264 8300 23276
rect 8352 23264 8358 23316
rect 9858 23304 9864 23316
rect 8404 23276 9864 23304
rect 4157 23239 4215 23245
rect 4157 23205 4169 23239
rect 4203 23236 4215 23239
rect 5534 23236 5540 23248
rect 4203 23208 5540 23236
rect 4203 23205 4215 23208
rect 4157 23199 4215 23205
rect 5534 23196 5540 23208
rect 5592 23196 5598 23248
rect 7006 23196 7012 23248
rect 7064 23196 7070 23248
rect 7834 23196 7840 23248
rect 7892 23196 7898 23248
rect 5442 23128 5448 23180
rect 5500 23168 5506 23180
rect 5997 23171 6055 23177
rect 5997 23168 6009 23171
rect 5500 23140 6009 23168
rect 5500 23128 5506 23140
rect 5997 23137 6009 23140
rect 6043 23137 6055 23171
rect 7852 23168 7880 23196
rect 8021 23171 8079 23177
rect 8021 23168 8033 23171
rect 7852 23140 8033 23168
rect 5997 23131 6055 23137
rect 8021 23137 8033 23140
rect 8067 23137 8079 23171
rect 8021 23131 8079 23137
rect 8205 23171 8263 23177
rect 8205 23137 8217 23171
rect 8251 23168 8263 23171
rect 8404 23168 8432 23276
rect 9858 23264 9864 23276
rect 9916 23264 9922 23316
rect 9950 23264 9956 23316
rect 10008 23304 10014 23316
rect 10689 23307 10747 23313
rect 10689 23304 10701 23307
rect 10008 23276 10701 23304
rect 10008 23264 10014 23276
rect 10689 23273 10701 23276
rect 10735 23273 10747 23307
rect 14274 23304 14280 23316
rect 10689 23267 10747 23273
rect 11808 23276 14280 23304
rect 9030 23236 9036 23248
rect 8680 23208 9036 23236
rect 8251 23140 8432 23168
rect 8481 23171 8539 23177
rect 8251 23137 8263 23140
rect 8205 23131 8263 23137
rect 8481 23137 8493 23171
rect 8527 23168 8539 23171
rect 8570 23168 8576 23180
rect 8527 23140 8576 23168
rect 8527 23137 8539 23140
rect 8481 23131 8539 23137
rect 8570 23128 8576 23140
rect 8628 23128 8634 23180
rect 8680 23177 8708 23208
rect 9030 23196 9036 23208
rect 9088 23196 9094 23248
rect 9214 23196 9220 23248
rect 9272 23236 9278 23248
rect 9272 23208 9996 23236
rect 9272 23196 9278 23208
rect 8665 23171 8723 23177
rect 8665 23137 8677 23171
rect 8711 23137 8723 23171
rect 8665 23131 8723 23137
rect 8757 23171 8815 23177
rect 8757 23137 8769 23171
rect 8803 23168 8815 23171
rect 9858 23168 9864 23180
rect 8803 23140 9864 23168
rect 8803 23137 8815 23140
rect 8757 23131 8815 23137
rect 9858 23128 9864 23140
rect 9916 23128 9922 23180
rect 9968 23177 9996 23208
rect 10134 23196 10140 23248
rect 10192 23196 10198 23248
rect 10226 23196 10232 23248
rect 10284 23236 10290 23248
rect 10284 23208 11376 23236
rect 10284 23196 10290 23208
rect 9953 23171 10011 23177
rect 9953 23137 9965 23171
rect 9999 23137 10011 23171
rect 9953 23131 10011 23137
rect 10594 23128 10600 23180
rect 10652 23128 10658 23180
rect 10796 23177 10824 23208
rect 11348 23180 11376 23208
rect 10757 23171 10824 23177
rect 10757 23137 10769 23171
rect 10803 23140 10824 23171
rect 10879 23171 10937 23177
rect 10803 23137 10815 23140
rect 10757 23131 10815 23137
rect 10879 23137 10891 23171
rect 10925 23137 10937 23171
rect 11057 23171 11115 23177
rect 11057 23168 11069 23171
rect 10879 23131 10937 23137
rect 10980 23140 11069 23168
rect 3418 23060 3424 23112
rect 3476 23060 3482 23112
rect 6273 23103 6331 23109
rect 6273 23069 6285 23103
rect 6319 23100 6331 23103
rect 7834 23100 7840 23112
rect 6319 23072 7840 23100
rect 6319 23069 6331 23072
rect 6273 23063 6331 23069
rect 7834 23060 7840 23072
rect 7892 23060 7898 23112
rect 8297 23103 8355 23109
rect 8297 23069 8309 23103
rect 8343 23100 8355 23103
rect 8849 23103 8907 23109
rect 8849 23100 8861 23103
rect 8343 23072 8861 23100
rect 8343 23069 8355 23072
rect 8297 23063 8355 23069
rect 8849 23069 8861 23072
rect 8895 23069 8907 23103
rect 8849 23063 8907 23069
rect 9030 23060 9036 23112
rect 9088 23100 9094 23112
rect 9490 23100 9496 23112
rect 9088 23072 9496 23100
rect 9088 23060 9094 23072
rect 9490 23060 9496 23072
rect 9548 23060 9554 23112
rect 9582 23060 9588 23112
rect 9640 23100 9646 23112
rect 9677 23103 9735 23109
rect 9677 23100 9689 23103
rect 9640 23072 9689 23100
rect 9640 23060 9646 23072
rect 9677 23069 9689 23072
rect 9723 23069 9735 23103
rect 10888 23100 10916 23131
rect 9677 23063 9735 23069
rect 9784 23072 10916 23100
rect 10980 23100 11008 23140
rect 11057 23137 11069 23140
rect 11103 23137 11115 23171
rect 11057 23131 11115 23137
rect 11330 23128 11336 23180
rect 11388 23128 11394 23180
rect 11808 23177 11836 23276
rect 14274 23264 14280 23276
rect 14332 23264 14338 23316
rect 14461 23307 14519 23313
rect 14461 23273 14473 23307
rect 14507 23304 14519 23307
rect 15286 23304 15292 23316
rect 14507 23276 15292 23304
rect 14507 23273 14519 23276
rect 14461 23267 14519 23273
rect 15286 23264 15292 23276
rect 15344 23264 15350 23316
rect 19702 23264 19708 23316
rect 19760 23304 19766 23316
rect 19797 23307 19855 23313
rect 19797 23304 19809 23307
rect 19760 23276 19809 23304
rect 19760 23264 19766 23276
rect 19797 23273 19809 23276
rect 19843 23304 19855 23307
rect 20346 23304 20352 23316
rect 19843 23276 20352 23304
rect 19843 23273 19855 23276
rect 19797 23267 19855 23273
rect 20346 23264 20352 23276
rect 20404 23264 20410 23316
rect 22189 23307 22247 23313
rect 22189 23273 22201 23307
rect 22235 23304 22247 23307
rect 22646 23304 22652 23316
rect 22235 23276 22652 23304
rect 22235 23273 22247 23276
rect 22189 23267 22247 23273
rect 22646 23264 22652 23276
rect 22704 23264 22710 23316
rect 25038 23264 25044 23316
rect 25096 23264 25102 23316
rect 26145 23307 26203 23313
rect 26145 23273 26157 23307
rect 26191 23304 26203 23307
rect 26326 23304 26332 23316
rect 26191 23276 26332 23304
rect 26191 23273 26203 23276
rect 26145 23267 26203 23273
rect 26326 23264 26332 23276
rect 26384 23264 26390 23316
rect 26602 23264 26608 23316
rect 26660 23264 26666 23316
rect 27430 23264 27436 23316
rect 27488 23304 27494 23316
rect 27801 23307 27859 23313
rect 27488 23276 27752 23304
rect 27488 23264 27494 23276
rect 14182 23236 14188 23248
rect 12360 23208 14188 23236
rect 11793 23171 11851 23177
rect 11793 23137 11805 23171
rect 11839 23137 11851 23171
rect 11793 23131 11851 23137
rect 11882 23128 11888 23180
rect 11940 23128 11946 23180
rect 12360 23177 12388 23208
rect 14182 23196 14188 23208
rect 14240 23236 14246 23248
rect 14369 23239 14427 23245
rect 14369 23236 14381 23239
rect 14240 23208 14381 23236
rect 14240 23196 14246 23208
rect 14369 23205 14381 23208
rect 14415 23205 14427 23239
rect 14369 23199 14427 23205
rect 16482 23196 16488 23248
rect 16540 23236 16546 23248
rect 18601 23239 18659 23245
rect 18601 23236 18613 23239
rect 16540 23208 18613 23236
rect 16540 23196 16546 23208
rect 18601 23205 18613 23208
rect 18647 23205 18659 23239
rect 18601 23199 18659 23205
rect 18800 23208 19288 23236
rect 12069 23171 12127 23177
rect 12069 23137 12081 23171
rect 12115 23137 12127 23171
rect 12069 23131 12127 23137
rect 12345 23171 12403 23177
rect 12345 23137 12357 23171
rect 12391 23137 12403 23171
rect 12345 23131 12403 23137
rect 12084 23100 12112 23131
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 12529 23171 12587 23177
rect 12529 23168 12541 23171
rect 12492 23140 12541 23168
rect 12492 23128 12498 23140
rect 12529 23137 12541 23140
rect 12575 23137 12587 23171
rect 12529 23131 12587 23137
rect 12710 23128 12716 23180
rect 12768 23128 12774 23180
rect 14918 23128 14924 23180
rect 14976 23128 14982 23180
rect 16574 23168 16580 23180
rect 16330 23140 16580 23168
rect 16574 23128 16580 23140
rect 16632 23128 16638 23180
rect 18509 23171 18567 23177
rect 18509 23137 18521 23171
rect 18555 23137 18567 23171
rect 18509 23131 18567 23137
rect 10980 23072 12112 23100
rect 12253 23103 12311 23109
rect 9784 23044 9812 23072
rect 10980 23044 11008 23072
rect 12253 23069 12265 23103
rect 12299 23100 12311 23103
rect 12299 23072 12572 23100
rect 12299 23069 12311 23072
rect 12253 23063 12311 23069
rect 3804 23004 6132 23032
rect 3804 22976 3832 23004
rect 3786 22924 3792 22976
rect 3844 22924 3850 22976
rect 4062 22924 4068 22976
rect 4120 22924 4126 22976
rect 4798 22924 4804 22976
rect 4856 22964 4862 22976
rect 5442 22964 5448 22976
rect 4856 22936 5448 22964
rect 4856 22924 4862 22936
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 6104 22964 6132 23004
rect 7944 23004 9628 23032
rect 7944 22964 7972 23004
rect 6104 22936 7972 22964
rect 8021 22967 8079 22973
rect 8021 22933 8033 22967
rect 8067 22964 8079 22967
rect 9214 22964 9220 22976
rect 8067 22936 9220 22964
rect 8067 22933 8079 22936
rect 8021 22927 8079 22933
rect 9214 22924 9220 22936
rect 9272 22924 9278 22976
rect 9490 22924 9496 22976
rect 9548 22924 9554 22976
rect 9600 22964 9628 23004
rect 9766 22992 9772 23044
rect 9824 22992 9830 23044
rect 10962 22992 10968 23044
rect 11020 22992 11026 23044
rect 11054 22992 11060 23044
rect 11112 22992 11118 23044
rect 12158 22992 12164 23044
rect 12216 22992 12222 23044
rect 11606 22964 11612 22976
rect 9600 22936 11612 22964
rect 11606 22924 11612 22936
rect 11664 22924 11670 22976
rect 12544 22964 12572 23072
rect 13722 23060 13728 23112
rect 13780 23060 13786 23112
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 14182 23100 14188 23112
rect 13872 23072 14188 23100
rect 13872 23060 13878 23072
rect 14182 23060 14188 23072
rect 14240 23060 14246 23112
rect 15194 23060 15200 23112
rect 15252 23060 15258 23112
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 15746 23100 15752 23112
rect 15344 23072 15752 23100
rect 15344 23060 15350 23072
rect 15746 23060 15752 23072
rect 15804 23060 15810 23112
rect 17129 23103 17187 23109
rect 17129 23100 17141 23103
rect 16868 23072 17141 23100
rect 16868 22976 16896 23072
rect 17129 23069 17141 23072
rect 17175 23069 17187 23103
rect 17129 23063 17187 23069
rect 17402 23060 17408 23112
rect 17460 23100 17466 23112
rect 18524 23100 18552 23131
rect 18690 23128 18696 23180
rect 18748 23128 18754 23180
rect 18800 23100 18828 23208
rect 19260 23180 19288 23208
rect 20162 23196 20168 23248
rect 20220 23236 20226 23248
rect 20257 23239 20315 23245
rect 20257 23236 20269 23239
rect 20220 23208 20269 23236
rect 20220 23196 20226 23208
rect 20257 23205 20269 23208
rect 20303 23205 20315 23239
rect 20257 23199 20315 23205
rect 20990 23196 20996 23248
rect 21048 23196 21054 23248
rect 26513 23239 26571 23245
rect 26513 23205 26525 23239
rect 26559 23205 26571 23239
rect 26513 23199 26571 23205
rect 18877 23171 18935 23177
rect 18877 23137 18889 23171
rect 18923 23168 18935 23171
rect 18923 23140 19104 23168
rect 18923 23137 18935 23140
rect 18877 23131 18935 23137
rect 17460 23072 18828 23100
rect 17460 23060 17466 23072
rect 19076 23032 19104 23140
rect 19242 23128 19248 23180
rect 19300 23128 19306 23180
rect 19978 23128 19984 23180
rect 20036 23128 20042 23180
rect 21818 23128 21824 23180
rect 21876 23168 21882 23180
rect 22557 23171 22615 23177
rect 22557 23168 22569 23171
rect 21876 23140 22569 23168
rect 21876 23128 21882 23140
rect 22557 23137 22569 23140
rect 22603 23137 22615 23171
rect 22557 23131 22615 23137
rect 22649 23171 22707 23177
rect 22649 23137 22661 23171
rect 22695 23168 22707 23171
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 22695 23140 23489 23168
rect 22695 23137 22707 23140
rect 22649 23131 22707 23137
rect 23477 23137 23489 23140
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 23658 23128 23664 23180
rect 23716 23168 23722 23180
rect 24029 23171 24087 23177
rect 24029 23168 24041 23171
rect 23716 23140 24041 23168
rect 23716 23128 23722 23140
rect 24029 23137 24041 23140
rect 24075 23137 24087 23171
rect 24029 23131 24087 23137
rect 24949 23171 25007 23177
rect 24949 23137 24961 23171
rect 24995 23168 25007 23171
rect 26329 23171 26387 23177
rect 24995 23140 25728 23168
rect 24995 23137 25007 23140
rect 24949 23131 25007 23137
rect 19150 23060 19156 23112
rect 19208 23100 19214 23112
rect 22741 23103 22799 23109
rect 22741 23100 22753 23103
rect 19208 23072 22753 23100
rect 19208 23060 19214 23072
rect 19076 23004 19288 23032
rect 12618 22964 12624 22976
rect 12544 22936 12624 22964
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 13078 22924 13084 22976
rect 13136 22964 13142 22976
rect 13173 22967 13231 22973
rect 13173 22964 13185 22967
rect 13136 22936 13185 22964
rect 13136 22924 13142 22936
rect 13173 22933 13185 22936
rect 13219 22933 13231 22967
rect 13173 22927 13231 22933
rect 14829 22967 14887 22973
rect 14829 22933 14841 22967
rect 14875 22964 14887 22967
rect 16298 22964 16304 22976
rect 14875 22936 16304 22964
rect 14875 22933 14887 22936
rect 14829 22927 14887 22933
rect 16298 22924 16304 22936
rect 16356 22924 16362 22976
rect 16669 22967 16727 22973
rect 16669 22933 16681 22967
rect 16715 22964 16727 22967
rect 16850 22964 16856 22976
rect 16715 22936 16856 22964
rect 16715 22933 16727 22936
rect 16669 22927 16727 22933
rect 16850 22924 16856 22936
rect 16908 22924 16914 22976
rect 17770 22924 17776 22976
rect 17828 22924 17834 22976
rect 18322 22924 18328 22976
rect 18380 22924 18386 22976
rect 19260 22973 19288 23004
rect 19245 22967 19303 22973
rect 19245 22933 19257 22967
rect 19291 22964 19303 22967
rect 19334 22964 19340 22976
rect 19291 22936 19340 22964
rect 19291 22933 19303 22936
rect 19245 22927 19303 22933
rect 19334 22924 19340 22936
rect 19392 22924 19398 22976
rect 21652 22964 21680 23072
rect 22741 23069 22753 23072
rect 22787 23069 22799 23103
rect 22741 23063 22799 23069
rect 23566 23060 23572 23112
rect 23624 23100 23630 23112
rect 25406 23100 25412 23112
rect 23624 23072 25412 23100
rect 23624 23060 23630 23072
rect 25406 23060 25412 23072
rect 25464 23060 25470 23112
rect 25700 23044 25728 23140
rect 26329 23137 26341 23171
rect 26375 23137 26387 23171
rect 26329 23131 26387 23137
rect 26421 23171 26479 23177
rect 26421 23137 26433 23171
rect 26467 23137 26479 23171
rect 26421 23131 26479 23137
rect 25866 23060 25872 23112
rect 25924 23060 25930 23112
rect 21729 23035 21787 23041
rect 21729 23001 21741 23035
rect 21775 23032 21787 23035
rect 25314 23032 25320 23044
rect 21775 23004 22324 23032
rect 21775 23001 21787 23004
rect 21729 22995 21787 23001
rect 22097 22967 22155 22973
rect 22097 22964 22109 22967
rect 21652 22936 22109 22964
rect 22097 22933 22109 22936
rect 22143 22933 22155 22967
rect 22296 22964 22324 23004
rect 22848 23004 25320 23032
rect 22848 22964 22876 23004
rect 25314 22992 25320 23004
rect 25372 22992 25378 23044
rect 25682 22992 25688 23044
rect 25740 22992 25746 23044
rect 22296 22936 22876 22964
rect 22097 22927 22155 22933
rect 24762 22924 24768 22976
rect 24820 22964 24826 22976
rect 25225 22967 25283 22973
rect 25225 22964 25237 22967
rect 24820 22936 25237 22964
rect 24820 22924 24826 22936
rect 25225 22933 25237 22936
rect 25271 22933 25283 22967
rect 26344 22964 26372 23131
rect 26436 23032 26464 23131
rect 26528 23112 26556 23199
rect 26620 23177 26648 23264
rect 27249 23239 27307 23245
rect 27249 23205 27261 23239
rect 27295 23236 27307 23239
rect 27724 23236 27752 23276
rect 27801 23273 27813 23307
rect 27847 23304 27859 23307
rect 28074 23304 28080 23316
rect 27847 23276 28080 23304
rect 27847 23273 27859 23276
rect 27801 23267 27859 23273
rect 28074 23264 28080 23276
rect 28132 23264 28138 23316
rect 30098 23264 30104 23316
rect 30156 23264 30162 23316
rect 27295 23208 27568 23236
rect 27724 23208 28120 23236
rect 27295 23205 27307 23208
rect 27249 23199 27307 23205
rect 26620 23171 26689 23177
rect 26620 23140 26643 23171
rect 26631 23137 26643 23140
rect 26677 23137 26689 23171
rect 26631 23131 26689 23137
rect 26789 23171 26847 23177
rect 26789 23137 26801 23171
rect 26835 23168 26847 23171
rect 27065 23171 27123 23177
rect 27065 23168 27077 23171
rect 26835 23140 27077 23168
rect 26835 23137 26847 23140
rect 26789 23131 26847 23137
rect 27065 23137 27077 23140
rect 27111 23168 27123 23171
rect 27338 23168 27344 23180
rect 27111 23140 27344 23168
rect 27111 23137 27123 23140
rect 27065 23131 27123 23137
rect 27338 23128 27344 23140
rect 27396 23128 27402 23180
rect 27540 23177 27568 23208
rect 27525 23171 27583 23177
rect 27525 23137 27537 23171
rect 27571 23168 27583 23171
rect 27614 23168 27620 23180
rect 27571 23140 27620 23168
rect 27571 23137 27583 23140
rect 27525 23131 27583 23137
rect 27614 23128 27620 23140
rect 27672 23168 27678 23180
rect 27798 23168 27804 23180
rect 27672 23140 27804 23168
rect 27672 23128 27678 23140
rect 27798 23128 27804 23140
rect 27856 23168 27862 23180
rect 28092 23177 28120 23208
rect 29288 23208 29960 23236
rect 27985 23171 28043 23177
rect 27985 23168 27997 23171
rect 27856 23140 27997 23168
rect 27856 23128 27862 23140
rect 27985 23137 27997 23140
rect 28031 23137 28043 23171
rect 27985 23131 28043 23137
rect 28077 23171 28135 23177
rect 28077 23137 28089 23171
rect 28123 23137 28135 23171
rect 28077 23131 28135 23137
rect 28261 23171 28319 23177
rect 28261 23137 28273 23171
rect 28307 23168 28319 23171
rect 28350 23168 28356 23180
rect 28307 23140 28356 23168
rect 28307 23137 28319 23140
rect 28261 23131 28319 23137
rect 28350 23128 28356 23140
rect 28408 23168 28414 23180
rect 28718 23168 28724 23180
rect 28408 23140 28724 23168
rect 28408 23128 28414 23140
rect 28718 23128 28724 23140
rect 28776 23128 28782 23180
rect 29086 23128 29092 23180
rect 29144 23168 29150 23180
rect 29288 23177 29316 23208
rect 29273 23171 29331 23177
rect 29273 23168 29285 23171
rect 29144 23140 29285 23168
rect 29144 23128 29150 23140
rect 29273 23137 29285 23140
rect 29319 23137 29331 23171
rect 29273 23131 29331 23137
rect 29641 23171 29699 23177
rect 29641 23137 29653 23171
rect 29687 23168 29699 23171
rect 29822 23168 29828 23180
rect 29687 23140 29828 23168
rect 29687 23137 29699 23140
rect 29641 23131 29699 23137
rect 26510 23060 26516 23112
rect 26568 23060 26574 23112
rect 27356 23100 27384 23128
rect 27356 23072 28028 23100
rect 28000 23044 28028 23072
rect 28166 23060 28172 23112
rect 28224 23060 28230 23112
rect 29656 23100 29684 23131
rect 29822 23128 29828 23140
rect 29880 23128 29886 23180
rect 28966 23072 29684 23100
rect 27433 23035 27491 23041
rect 27433 23032 27445 23035
rect 26436 23004 27445 23032
rect 27433 23001 27445 23004
rect 27479 23001 27491 23035
rect 27433 22995 27491 23001
rect 27706 22992 27712 23044
rect 27764 22992 27770 23044
rect 27982 22992 27988 23044
rect 28040 22992 28046 23044
rect 26881 22967 26939 22973
rect 26881 22964 26893 22967
rect 26344 22936 26893 22964
rect 25225 22927 25283 22933
rect 26881 22933 26893 22936
rect 26927 22933 26939 22967
rect 27724 22964 27752 22992
rect 28966 22964 28994 23072
rect 29932 23032 29960 23208
rect 30116 23168 30144 23264
rect 30193 23171 30251 23177
rect 30193 23168 30205 23171
rect 30116 23140 30205 23168
rect 30193 23137 30205 23140
rect 30239 23137 30251 23171
rect 30193 23131 30251 23137
rect 31110 23128 31116 23180
rect 31168 23128 31174 23180
rect 31754 23168 31760 23180
rect 31312 23140 31760 23168
rect 30006 23060 30012 23112
rect 30064 23100 30070 23112
rect 31205 23103 31263 23109
rect 31205 23100 31217 23103
rect 30064 23072 31217 23100
rect 30064 23060 30070 23072
rect 31205 23069 31217 23072
rect 31251 23069 31263 23103
rect 31205 23063 31263 23069
rect 31312 23032 31340 23140
rect 31754 23128 31760 23140
rect 31812 23128 31818 23180
rect 29932 23004 31340 23032
rect 27724 22936 28994 22964
rect 26881 22927 26939 22933
rect 29638 22924 29644 22976
rect 29696 22924 29702 22976
rect 29822 22924 29828 22976
rect 29880 22924 29886 22976
rect 30098 22924 30104 22976
rect 30156 22964 30162 22976
rect 30285 22967 30343 22973
rect 30285 22964 30297 22967
rect 30156 22936 30297 22964
rect 30156 22924 30162 22936
rect 30285 22933 30297 22936
rect 30331 22933 30343 22967
rect 30285 22927 30343 22933
rect 30926 22924 30932 22976
rect 30984 22924 30990 22976
rect 2760 22874 34316 22896
rect 2760 22822 6550 22874
rect 6602 22822 6614 22874
rect 6666 22822 6678 22874
rect 6730 22822 6742 22874
rect 6794 22822 6806 22874
rect 6858 22822 14439 22874
rect 14491 22822 14503 22874
rect 14555 22822 14567 22874
rect 14619 22822 14631 22874
rect 14683 22822 14695 22874
rect 14747 22822 22328 22874
rect 22380 22822 22392 22874
rect 22444 22822 22456 22874
rect 22508 22822 22520 22874
rect 22572 22822 22584 22874
rect 22636 22822 30217 22874
rect 30269 22822 30281 22874
rect 30333 22822 30345 22874
rect 30397 22822 30409 22874
rect 30461 22822 30473 22874
rect 30525 22822 34316 22874
rect 2760 22800 34316 22822
rect 3050 22720 3056 22772
rect 3108 22720 3114 22772
rect 5626 22720 5632 22772
rect 5684 22760 5690 22772
rect 6089 22763 6147 22769
rect 6089 22760 6101 22763
rect 5684 22732 6101 22760
rect 5684 22720 5690 22732
rect 6089 22729 6101 22732
rect 6135 22729 6147 22763
rect 6089 22723 6147 22729
rect 9214 22720 9220 22772
rect 9272 22720 9278 22772
rect 9858 22720 9864 22772
rect 9916 22760 9922 22772
rect 10318 22760 10324 22772
rect 9916 22732 10324 22760
rect 9916 22720 9922 22732
rect 10318 22720 10324 22732
rect 10376 22760 10382 22772
rect 10413 22763 10471 22769
rect 10413 22760 10425 22763
rect 10376 22732 10425 22760
rect 10376 22720 10382 22732
rect 10413 22729 10425 22732
rect 10459 22729 10471 22763
rect 10413 22723 10471 22729
rect 12529 22763 12587 22769
rect 12529 22729 12541 22763
rect 12575 22760 12587 22763
rect 13722 22760 13728 22772
rect 12575 22732 13728 22760
rect 12575 22729 12587 22732
rect 12529 22723 12587 22729
rect 13722 22720 13728 22732
rect 13780 22720 13786 22772
rect 14461 22763 14519 22769
rect 14461 22729 14473 22763
rect 14507 22760 14519 22763
rect 14826 22760 14832 22772
rect 14507 22732 14832 22760
rect 14507 22729 14519 22732
rect 14461 22723 14519 22729
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 15194 22720 15200 22772
rect 15252 22760 15258 22772
rect 15749 22763 15807 22769
rect 15749 22760 15761 22763
rect 15252 22732 15761 22760
rect 15252 22720 15258 22732
rect 15749 22729 15761 22732
rect 15795 22729 15807 22763
rect 15749 22723 15807 22729
rect 16298 22720 16304 22772
rect 16356 22720 16362 22772
rect 16574 22720 16580 22772
rect 16632 22720 16638 22772
rect 17773 22763 17831 22769
rect 17773 22729 17785 22763
rect 17819 22760 17831 22763
rect 17862 22760 17868 22772
rect 17819 22732 17868 22760
rect 17819 22729 17831 22732
rect 17773 22723 17831 22729
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 18322 22720 18328 22772
rect 18380 22720 18386 22772
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 19978 22760 19984 22772
rect 19668 22732 19984 22760
rect 19668 22720 19674 22732
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 24292 22763 24350 22769
rect 24292 22729 24304 22763
rect 24338 22760 24350 22763
rect 24762 22760 24768 22772
rect 24338 22732 24768 22760
rect 24338 22729 24350 22732
rect 24292 22723 24350 22729
rect 24762 22720 24768 22732
rect 24820 22720 24826 22772
rect 25866 22720 25872 22772
rect 25924 22760 25930 22772
rect 26145 22763 26203 22769
rect 26145 22760 26157 22763
rect 25924 22732 26157 22760
rect 25924 22720 25930 22732
rect 26145 22729 26157 22732
rect 26191 22729 26203 22763
rect 28166 22760 28172 22772
rect 26145 22723 26203 22729
rect 26331 22732 28172 22760
rect 8938 22652 8944 22704
rect 8996 22692 9002 22704
rect 8996 22664 10824 22692
rect 8996 22652 9002 22664
rect 4062 22584 4068 22636
rect 4120 22624 4126 22636
rect 4525 22627 4583 22633
rect 4525 22624 4537 22627
rect 4120 22596 4537 22624
rect 4120 22584 4126 22596
rect 4525 22593 4537 22596
rect 4571 22593 4583 22627
rect 6733 22627 6791 22633
rect 6733 22624 6745 22627
rect 4525 22587 4583 22593
rect 4816 22596 6745 22624
rect 4816 22568 4844 22596
rect 6733 22593 6745 22596
rect 6779 22593 6791 22627
rect 6733 22587 6791 22593
rect 7009 22627 7067 22633
rect 7009 22593 7021 22627
rect 7055 22624 7067 22627
rect 8849 22627 8907 22633
rect 8849 22624 8861 22627
rect 7055 22596 8861 22624
rect 7055 22593 7067 22596
rect 7009 22587 7067 22593
rect 8849 22593 8861 22596
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 9048 22596 9536 22624
rect 4798 22516 4804 22568
rect 4856 22516 4862 22568
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 5442 22516 5448 22568
rect 5500 22516 5506 22568
rect 9048 22565 9076 22596
rect 9508 22568 9536 22596
rect 9033 22559 9091 22565
rect 9033 22525 9045 22559
rect 9079 22525 9091 22559
rect 9033 22519 9091 22525
rect 9309 22559 9367 22565
rect 9309 22525 9321 22559
rect 9355 22525 9367 22559
rect 9309 22519 9367 22525
rect 4985 22491 5043 22497
rect 4985 22488 4997 22491
rect 4094 22460 4997 22488
rect 4985 22457 4997 22460
rect 5031 22457 5043 22491
rect 4985 22451 5043 22457
rect 4706 22380 4712 22432
rect 4764 22420 4770 22432
rect 5092 22420 5120 22516
rect 7742 22448 7748 22500
rect 7800 22448 7806 22500
rect 9324 22488 9352 22519
rect 9490 22516 9496 22568
rect 9548 22516 9554 22568
rect 9766 22516 9772 22568
rect 9824 22516 9830 22568
rect 10796 22565 10824 22664
rect 10962 22652 10968 22704
rect 11020 22692 11026 22704
rect 11020 22664 11468 22692
rect 11020 22652 11026 22664
rect 11440 22568 11468 22664
rect 11882 22652 11888 22704
rect 11940 22692 11946 22704
rect 11940 22664 12113 22692
rect 11940 22652 11946 22664
rect 11974 22584 11980 22636
rect 12032 22584 12038 22636
rect 12085 22624 12113 22664
rect 12345 22627 12403 22633
rect 12345 22624 12357 22627
rect 12085 22596 12357 22624
rect 12345 22593 12357 22596
rect 12391 22593 12403 22627
rect 12345 22587 12403 22593
rect 12989 22627 13047 22633
rect 12989 22593 13001 22627
rect 13035 22624 13047 22627
rect 13078 22624 13084 22636
rect 13035 22596 13084 22624
rect 13035 22593 13047 22596
rect 12989 22587 13047 22593
rect 13078 22584 13084 22596
rect 13136 22584 13142 22636
rect 16316 22633 16344 22720
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22593 16359 22627
rect 18340 22624 18368 22720
rect 19797 22627 19855 22633
rect 19797 22624 19809 22627
rect 18340 22596 19809 22624
rect 16301 22587 16359 22593
rect 19797 22593 19809 22596
rect 19843 22593 19855 22627
rect 19996 22624 20024 22720
rect 20717 22695 20775 22701
rect 20717 22661 20729 22695
rect 20763 22692 20775 22695
rect 20763 22664 22094 22692
rect 20763 22661 20775 22664
rect 20717 22655 20775 22661
rect 20073 22627 20131 22633
rect 20073 22624 20085 22627
rect 19996 22596 20085 22624
rect 19797 22587 19855 22593
rect 20073 22593 20085 22596
rect 20119 22593 20131 22627
rect 22066 22624 22094 22664
rect 22465 22627 22523 22633
rect 22465 22624 22477 22627
rect 20073 22587 20131 22593
rect 21100 22596 21312 22624
rect 22066 22596 22477 22624
rect 21100 22568 21128 22596
rect 10781 22559 10839 22565
rect 10781 22525 10793 22559
rect 10827 22525 10839 22559
rect 10781 22519 10839 22525
rect 10870 22516 10876 22568
rect 10928 22556 10934 22568
rect 11149 22559 11207 22565
rect 11149 22556 11161 22559
rect 10928 22528 11161 22556
rect 10928 22516 10934 22528
rect 11149 22525 11161 22528
rect 11195 22556 11207 22559
rect 11238 22556 11244 22568
rect 11195 22528 11244 22556
rect 11195 22525 11207 22528
rect 11149 22519 11207 22525
rect 11238 22516 11244 22528
rect 11296 22516 11302 22568
rect 11422 22516 11428 22568
rect 11480 22516 11486 22568
rect 11606 22516 11612 22568
rect 11664 22556 11670 22568
rect 11885 22559 11943 22565
rect 11885 22556 11897 22559
rect 11664 22528 11897 22556
rect 11664 22516 11670 22528
rect 11885 22525 11897 22528
rect 11931 22525 11943 22559
rect 11885 22519 11943 22525
rect 12253 22559 12311 22565
rect 12253 22525 12265 22559
rect 12299 22556 12311 22559
rect 12618 22556 12624 22568
rect 12299 22528 12624 22556
rect 12299 22525 12311 22528
rect 12253 22519 12311 22525
rect 9582 22488 9588 22500
rect 9324 22460 9588 22488
rect 9582 22448 9588 22460
rect 9640 22488 9646 22500
rect 10597 22491 10655 22497
rect 10597 22488 10609 22491
rect 9640 22460 10609 22488
rect 9640 22448 9646 22460
rect 9968 22432 9996 22460
rect 10597 22457 10609 22460
rect 10643 22457 10655 22491
rect 12268 22488 12296 22519
rect 12618 22516 12624 22528
rect 12676 22516 12682 22568
rect 12710 22516 12716 22568
rect 12768 22516 12774 22568
rect 14090 22516 14096 22568
rect 14148 22516 14154 22568
rect 15010 22516 15016 22568
rect 15068 22556 15074 22568
rect 15473 22559 15531 22565
rect 15473 22556 15485 22559
rect 15068 22528 15485 22556
rect 15068 22516 15074 22528
rect 15473 22525 15485 22528
rect 15519 22525 15531 22559
rect 15473 22519 15531 22525
rect 16666 22516 16672 22568
rect 16724 22516 16730 22568
rect 17218 22516 17224 22568
rect 17276 22556 17282 22568
rect 17862 22556 17868 22568
rect 17276 22528 17868 22556
rect 17276 22516 17282 22528
rect 17862 22516 17868 22528
rect 17920 22516 17926 22568
rect 18230 22556 18236 22568
rect 18064 22528 18236 22556
rect 10597 22451 10655 22457
rect 11348 22460 12296 22488
rect 11348 22432 11376 22460
rect 4764 22392 5120 22420
rect 4764 22380 4770 22392
rect 5994 22380 6000 22432
rect 6052 22420 6058 22432
rect 6454 22420 6460 22432
rect 6052 22392 6460 22420
rect 6052 22380 6058 22392
rect 6454 22380 6460 22392
rect 6512 22420 6518 22432
rect 6549 22423 6607 22429
rect 6549 22420 6561 22423
rect 6512 22392 6561 22420
rect 6512 22380 6518 22392
rect 6549 22389 6561 22392
rect 6595 22389 6607 22423
rect 6549 22383 6607 22389
rect 8481 22423 8539 22429
rect 8481 22389 8493 22423
rect 8527 22420 8539 22423
rect 9030 22420 9036 22432
rect 8527 22392 9036 22420
rect 8527 22389 8539 22392
rect 8481 22383 8539 22389
rect 9030 22380 9036 22392
rect 9088 22380 9094 22432
rect 9950 22380 9956 22432
rect 10008 22380 10014 22432
rect 11330 22380 11336 22432
rect 11388 22380 11394 22432
rect 11790 22380 11796 22432
rect 11848 22420 11854 22432
rect 12069 22423 12127 22429
rect 12069 22420 12081 22423
rect 11848 22392 12081 22420
rect 11848 22380 11854 22392
rect 12069 22389 12081 22392
rect 12115 22420 12127 22423
rect 12434 22420 12440 22432
rect 12115 22392 12440 22420
rect 12115 22389 12127 22392
rect 12069 22383 12127 22389
rect 12434 22380 12440 22392
rect 12492 22380 12498 22432
rect 14826 22380 14832 22432
rect 14884 22420 14890 22432
rect 14921 22423 14979 22429
rect 14921 22420 14933 22423
rect 14884 22392 14933 22420
rect 14884 22380 14890 22392
rect 14921 22389 14933 22392
rect 14967 22389 14979 22423
rect 14921 22383 14979 22389
rect 17954 22380 17960 22432
rect 18012 22420 18018 22432
rect 18064 22429 18092 22528
rect 18230 22516 18236 22528
rect 18288 22516 18294 22568
rect 18414 22516 18420 22568
rect 18472 22516 18478 22568
rect 20165 22559 20223 22565
rect 20165 22525 20177 22559
rect 20211 22525 20223 22559
rect 20165 22519 20223 22525
rect 18049 22423 18107 22429
rect 18049 22420 18061 22423
rect 18012 22392 18061 22420
rect 18012 22380 18018 22392
rect 18049 22389 18061 22392
rect 18095 22389 18107 22423
rect 18049 22383 18107 22389
rect 18325 22423 18383 22429
rect 18325 22389 18337 22423
rect 18371 22420 18383 22423
rect 18432 22420 18460 22516
rect 19058 22448 19064 22500
rect 19116 22448 19122 22500
rect 19702 22448 19708 22500
rect 19760 22488 19766 22500
rect 20180 22488 20208 22519
rect 20346 22516 20352 22568
rect 20404 22516 20410 22568
rect 20530 22516 20536 22568
rect 20588 22516 20594 22568
rect 21082 22516 21088 22568
rect 21140 22516 21146 22568
rect 21174 22516 21180 22568
rect 21232 22516 21238 22568
rect 21284 22556 21312 22596
rect 22465 22593 22477 22596
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 24026 22584 24032 22636
rect 24084 22584 24090 22636
rect 25777 22627 25835 22633
rect 25777 22593 25789 22627
rect 25823 22624 25835 22627
rect 26331 22624 26359 22732
rect 26694 22652 26700 22704
rect 26752 22652 26758 22704
rect 26712 22624 26740 22652
rect 25823 22596 26359 22624
rect 26666 22596 26740 22624
rect 26789 22627 26847 22633
rect 25823 22593 25835 22596
rect 25777 22587 25835 22593
rect 22646 22556 22652 22568
rect 21284 22528 22652 22556
rect 22646 22516 22652 22528
rect 22704 22556 22710 22568
rect 23750 22556 23756 22568
rect 22704 22528 23756 22556
rect 22704 22516 22710 22528
rect 23750 22516 23756 22528
rect 23808 22556 23814 22568
rect 23808 22528 23980 22556
rect 23808 22516 23814 22528
rect 19760 22460 20208 22488
rect 20441 22491 20499 22497
rect 19760 22448 19766 22460
rect 20441 22457 20453 22491
rect 20487 22488 20499 22491
rect 21818 22488 21824 22500
rect 20487 22460 21824 22488
rect 20487 22457 20499 22460
rect 20441 22451 20499 22457
rect 21818 22448 21824 22460
rect 21876 22448 21882 22500
rect 18371 22392 18460 22420
rect 18371 22389 18383 22392
rect 18325 22383 18383 22389
rect 20990 22380 20996 22432
rect 21048 22380 21054 22432
rect 21910 22380 21916 22432
rect 21968 22380 21974 22432
rect 22830 22380 22836 22432
rect 22888 22380 22894 22432
rect 23842 22380 23848 22432
rect 23900 22380 23906 22432
rect 23952 22420 23980 22528
rect 25406 22516 25412 22568
rect 25464 22516 25470 22568
rect 26326 22516 26332 22568
rect 26384 22516 26390 22568
rect 26666 22565 26694 22596
rect 26789 22593 26801 22627
rect 26835 22593 26847 22627
rect 26789 22587 26847 22593
rect 26881 22627 26939 22633
rect 26881 22593 26893 22627
rect 26927 22624 26939 22627
rect 26988 22624 27016 22732
rect 28166 22720 28172 22732
rect 28224 22720 28230 22772
rect 31021 22763 31079 22769
rect 31021 22729 31033 22763
rect 31067 22760 31079 22763
rect 31110 22760 31116 22772
rect 31067 22732 31116 22760
rect 31067 22729 31079 22732
rect 31021 22723 31079 22729
rect 31110 22720 31116 22732
rect 31168 22720 31174 22772
rect 31202 22720 31208 22772
rect 31260 22760 31266 22772
rect 31297 22763 31355 22769
rect 31297 22760 31309 22763
rect 31260 22732 31309 22760
rect 31260 22720 31266 22732
rect 31297 22729 31309 22732
rect 31343 22760 31355 22763
rect 31754 22760 31760 22772
rect 31343 22732 31760 22760
rect 31343 22729 31355 22732
rect 31297 22723 31355 22729
rect 31754 22720 31760 22732
rect 31812 22720 31818 22772
rect 27890 22652 27896 22704
rect 27948 22692 27954 22704
rect 28350 22692 28356 22704
rect 27948 22664 28356 22692
rect 27948 22652 27954 22664
rect 28350 22652 28356 22664
rect 28408 22652 28414 22704
rect 26927 22596 27016 22624
rect 27157 22627 27215 22633
rect 26927 22593 26939 22596
rect 26881 22587 26939 22593
rect 27157 22593 27169 22627
rect 27203 22593 27215 22627
rect 27157 22587 27215 22593
rect 26651 22559 26709 22565
rect 26651 22525 26663 22559
rect 26697 22525 26709 22559
rect 26651 22519 26709 22525
rect 26418 22448 26424 22500
rect 26476 22448 26482 22500
rect 26510 22448 26516 22500
rect 26568 22448 26574 22500
rect 26804 22488 26832 22587
rect 27172 22556 27200 22587
rect 29178 22584 29184 22636
rect 29236 22624 29242 22636
rect 29273 22627 29331 22633
rect 29273 22624 29285 22627
rect 29236 22596 29285 22624
rect 29236 22584 29242 22596
rect 29273 22593 29285 22596
rect 29319 22624 29331 22627
rect 31570 22624 31576 22636
rect 29319 22596 31576 22624
rect 29319 22593 29331 22596
rect 29273 22587 29331 22593
rect 31570 22584 31576 22596
rect 31628 22624 31634 22636
rect 33045 22627 33103 22633
rect 33045 22624 33057 22627
rect 31628 22596 33057 22624
rect 31628 22584 31634 22596
rect 33045 22593 33057 22596
rect 33091 22593 33103 22627
rect 33410 22624 33416 22636
rect 33045 22587 33103 22593
rect 33336 22596 33416 22624
rect 28077 22559 28135 22565
rect 28077 22556 28089 22559
rect 27172 22528 28089 22556
rect 27062 22488 27068 22500
rect 26804 22460 27068 22488
rect 27062 22448 27068 22460
rect 27120 22488 27126 22500
rect 27172 22488 27200 22528
rect 28077 22525 28089 22528
rect 28123 22525 28135 22559
rect 28077 22519 28135 22525
rect 28261 22559 28319 22565
rect 28261 22525 28273 22559
rect 28307 22556 28319 22559
rect 28442 22556 28448 22568
rect 28307 22528 28448 22556
rect 28307 22525 28319 22528
rect 28261 22519 28319 22525
rect 28442 22516 28448 22528
rect 28500 22516 28506 22568
rect 33336 22565 33364 22596
rect 33410 22584 33416 22596
rect 33468 22584 33474 22636
rect 33321 22559 33379 22565
rect 33321 22525 33333 22559
rect 33367 22525 33379 22559
rect 33321 22519 33379 22525
rect 33965 22559 34023 22565
rect 33965 22525 33977 22559
rect 34011 22556 34023 22559
rect 35158 22556 35164 22568
rect 34011 22528 35164 22556
rect 34011 22525 34023 22528
rect 33965 22519 34023 22525
rect 35158 22516 35164 22528
rect 35216 22516 35222 22568
rect 27120 22460 27200 22488
rect 27120 22448 27126 22460
rect 29546 22448 29552 22500
rect 29604 22448 29610 22500
rect 30098 22448 30104 22500
rect 30156 22448 30162 22500
rect 32338 22460 32444 22488
rect 25682 22420 25688 22432
rect 23952 22392 25688 22420
rect 25682 22380 25688 22392
rect 25740 22380 25746 22432
rect 26528 22420 26556 22448
rect 27154 22420 27160 22432
rect 26528 22392 27160 22420
rect 27154 22380 27160 22392
rect 27212 22380 27218 22432
rect 28166 22380 28172 22432
rect 28224 22380 28230 22432
rect 28442 22380 28448 22432
rect 28500 22380 28506 22432
rect 32416 22420 32444 22460
rect 32766 22448 32772 22500
rect 32824 22448 32830 22500
rect 33229 22491 33287 22497
rect 33229 22457 33241 22491
rect 33275 22457 33287 22491
rect 33229 22451 33287 22457
rect 33244 22420 33272 22451
rect 32416 22392 33272 22420
rect 33778 22380 33784 22432
rect 33836 22380 33842 22432
rect 2760 22330 34316 22352
rect 2760 22278 7210 22330
rect 7262 22278 7274 22330
rect 7326 22278 7338 22330
rect 7390 22278 7402 22330
rect 7454 22278 7466 22330
rect 7518 22278 15099 22330
rect 15151 22278 15163 22330
rect 15215 22278 15227 22330
rect 15279 22278 15291 22330
rect 15343 22278 15355 22330
rect 15407 22278 22988 22330
rect 23040 22278 23052 22330
rect 23104 22278 23116 22330
rect 23168 22278 23180 22330
rect 23232 22278 23244 22330
rect 23296 22278 30877 22330
rect 30929 22278 30941 22330
rect 30993 22278 31005 22330
rect 31057 22278 31069 22330
rect 31121 22278 31133 22330
rect 31185 22278 34316 22330
rect 2760 22256 34316 22278
rect 3050 22176 3056 22228
rect 3108 22176 3114 22228
rect 3418 22176 3424 22228
rect 3476 22176 3482 22228
rect 3881 22219 3939 22225
rect 3881 22216 3893 22219
rect 3528 22188 3893 22216
rect 3068 22148 3096 22176
rect 3528 22148 3556 22188
rect 3881 22185 3893 22188
rect 3927 22185 3939 22219
rect 4706 22216 4712 22228
rect 3881 22179 3939 22185
rect 4172 22188 4712 22216
rect 3068 22120 3556 22148
rect 3786 22108 3792 22160
rect 3844 22108 3850 22160
rect 3329 22083 3387 22089
rect 3329 22049 3341 22083
rect 3375 22080 3387 22083
rect 4172 22080 4200 22188
rect 4706 22176 4712 22188
rect 4764 22176 4770 22228
rect 5350 22176 5356 22228
rect 5408 22216 5414 22228
rect 5997 22219 6055 22225
rect 5997 22216 6009 22219
rect 5408 22188 6009 22216
rect 5408 22176 5414 22188
rect 5997 22185 6009 22188
rect 6043 22185 6055 22219
rect 5997 22179 6055 22185
rect 7742 22176 7748 22228
rect 7800 22176 7806 22228
rect 7834 22176 7840 22228
rect 7892 22216 7898 22228
rect 8021 22219 8079 22225
rect 8021 22216 8033 22219
rect 7892 22188 8033 22216
rect 7892 22176 7898 22188
rect 8021 22185 8033 22188
rect 8067 22185 8079 22219
rect 8021 22179 8079 22185
rect 8389 22219 8447 22225
rect 8389 22185 8401 22219
rect 8435 22216 8447 22219
rect 8938 22216 8944 22228
rect 8435 22188 8944 22216
rect 8435 22185 8447 22188
rect 8389 22179 8447 22185
rect 8938 22176 8944 22188
rect 8996 22176 9002 22228
rect 9490 22176 9496 22228
rect 9548 22176 9554 22228
rect 9677 22219 9735 22225
rect 9677 22185 9689 22219
rect 9723 22216 9735 22219
rect 9766 22216 9772 22228
rect 9723 22188 9772 22216
rect 9723 22185 9735 22188
rect 9677 22179 9735 22185
rect 9766 22176 9772 22188
rect 9824 22176 9830 22228
rect 12158 22216 12164 22228
rect 9876 22188 11100 22216
rect 4798 22148 4804 22160
rect 4264 22120 4804 22148
rect 4264 22089 4292 22120
rect 4798 22108 4804 22120
rect 4856 22108 4862 22160
rect 8110 22148 8116 22160
rect 7668 22120 8116 22148
rect 7668 22089 7696 22120
rect 8110 22108 8116 22120
rect 8168 22108 8174 22160
rect 9508 22148 9536 22176
rect 9876 22157 9904 22188
rect 11072 22160 11100 22188
rect 11256 22188 12164 22216
rect 9048 22120 9536 22148
rect 9861 22151 9919 22157
rect 3375 22052 4200 22080
rect 4238 22083 4296 22089
rect 3375 22049 3387 22052
rect 3329 22043 3387 22049
rect 4238 22049 4250 22083
rect 4284 22049 4296 22083
rect 6181 22083 6239 22089
rect 6181 22080 6193 22083
rect 5658 22052 6193 22080
rect 4238 22043 4296 22049
rect 6181 22049 6193 22052
rect 6227 22049 6239 22083
rect 6181 22043 6239 22049
rect 6273 22083 6331 22089
rect 6273 22049 6285 22083
rect 6319 22080 6331 22083
rect 7653 22083 7711 22089
rect 7653 22080 7665 22083
rect 6319 22052 7665 22080
rect 6319 22049 6331 22052
rect 6273 22043 6331 22049
rect 7653 22049 7665 22052
rect 7699 22049 7711 22083
rect 7653 22043 7711 22049
rect 8205 22083 8263 22089
rect 8205 22049 8217 22083
rect 8251 22080 8263 22083
rect 8294 22080 8300 22092
rect 8251 22052 8300 22080
rect 8251 22049 8263 22052
rect 8205 22043 8263 22049
rect 4065 22015 4123 22021
rect 4065 21981 4077 22015
rect 4111 22012 4123 22015
rect 4111 21984 4384 22012
rect 4111 21981 4123 21984
rect 4065 21975 4123 21981
rect 3234 21836 3240 21888
rect 3292 21836 3298 21888
rect 4246 21836 4252 21888
rect 4304 21876 4310 21888
rect 4356 21876 4384 21984
rect 4522 21972 4528 22024
rect 4580 21972 4586 22024
rect 5074 21972 5080 22024
rect 5132 22012 5138 22024
rect 5258 22012 5264 22024
rect 5132 21984 5264 22012
rect 5132 21972 5138 21984
rect 5258 21972 5264 21984
rect 5316 22012 5322 22024
rect 6288 22012 6316 22043
rect 8294 22040 8300 22052
rect 8352 22040 8358 22092
rect 8481 22083 8539 22089
rect 8481 22049 8493 22083
rect 8527 22080 8539 22083
rect 9048 22080 9076 22120
rect 9861 22117 9873 22151
rect 9907 22117 9919 22151
rect 9861 22111 9919 22117
rect 10045 22151 10103 22157
rect 10045 22117 10057 22151
rect 10091 22148 10103 22151
rect 10226 22148 10232 22160
rect 10091 22120 10232 22148
rect 10091 22117 10103 22120
rect 10045 22111 10103 22117
rect 10226 22108 10232 22120
rect 10284 22108 10290 22160
rect 11054 22108 11060 22160
rect 11112 22108 11118 22160
rect 8527 22052 9076 22080
rect 10137 22083 10195 22089
rect 8527 22049 8539 22052
rect 8481 22043 8539 22049
rect 10137 22049 10149 22083
rect 10183 22049 10195 22083
rect 10137 22043 10195 22049
rect 5316 21984 6316 22012
rect 5316 21972 5322 21984
rect 9030 21972 9036 22024
rect 9088 21972 9094 22024
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 10152 22012 10180 22043
rect 10318 22040 10324 22092
rect 10376 22040 10382 22092
rect 11256 22080 11284 22188
rect 12158 22176 12164 22188
rect 12216 22176 12222 22228
rect 16209 22219 16267 22225
rect 16209 22185 16221 22219
rect 16255 22216 16267 22219
rect 17218 22216 17224 22228
rect 16255 22188 17224 22216
rect 16255 22185 16267 22188
rect 16209 22179 16267 22185
rect 17218 22176 17224 22188
rect 17276 22176 17282 22228
rect 17770 22176 17776 22228
rect 17828 22216 17834 22228
rect 19981 22219 20039 22225
rect 17828 22188 18460 22216
rect 17828 22176 17834 22188
rect 11701 22151 11759 22157
rect 11701 22117 11713 22151
rect 11747 22148 11759 22151
rect 13173 22151 13231 22157
rect 13173 22148 13185 22151
rect 11747 22120 13185 22148
rect 11747 22117 11759 22120
rect 11701 22111 11759 22117
rect 13173 22117 13185 22120
rect 13219 22117 13231 22151
rect 13173 22111 13231 22117
rect 14737 22151 14795 22157
rect 14737 22117 14749 22151
rect 14783 22148 14795 22151
rect 14826 22148 14832 22160
rect 14783 22120 14832 22148
rect 14783 22117 14795 22120
rect 14737 22111 14795 22117
rect 14826 22108 14832 22120
rect 14884 22108 14890 22160
rect 17957 22151 18015 22157
rect 17957 22117 17969 22151
rect 18003 22148 18015 22151
rect 18322 22148 18328 22160
rect 18003 22120 18328 22148
rect 18003 22117 18015 22120
rect 17957 22111 18015 22117
rect 18322 22108 18328 22120
rect 18380 22108 18386 22160
rect 18432 22157 18460 22188
rect 19981 22185 19993 22219
rect 20027 22216 20039 22219
rect 21174 22216 21180 22228
rect 20027 22188 21180 22216
rect 20027 22185 20039 22188
rect 19981 22179 20039 22185
rect 21174 22176 21180 22188
rect 21232 22176 21238 22228
rect 21910 22216 21916 22228
rect 21468 22188 21916 22216
rect 18417 22151 18475 22157
rect 18417 22117 18429 22151
rect 18463 22117 18475 22151
rect 18417 22111 18475 22117
rect 20990 22108 20996 22160
rect 21048 22108 21054 22160
rect 21468 22157 21496 22188
rect 21910 22176 21916 22188
rect 21968 22176 21974 22228
rect 22646 22216 22652 22228
rect 22296 22188 22652 22216
rect 21453 22151 21511 22157
rect 21453 22117 21465 22151
rect 21499 22117 21511 22151
rect 21453 22111 21511 22117
rect 10428 22052 11284 22080
rect 10428 22012 10456 22052
rect 11514 22040 11520 22092
rect 11572 22080 11578 22092
rect 12069 22083 12127 22089
rect 12069 22080 12081 22083
rect 11572 22052 12081 22080
rect 11572 22040 11578 22052
rect 12069 22049 12081 22052
rect 12115 22049 12127 22083
rect 12069 22043 12127 22049
rect 12342 22040 12348 22092
rect 12400 22040 12406 22092
rect 13538 22040 13544 22092
rect 13596 22080 13602 22092
rect 14093 22083 14151 22089
rect 14093 22080 14105 22083
rect 13596 22052 14105 22080
rect 13596 22040 13602 22052
rect 14093 22049 14105 22052
rect 14139 22049 14151 22083
rect 14093 22043 14151 22049
rect 15838 22040 15844 22092
rect 15896 22040 15902 22092
rect 16945 22083 17003 22089
rect 16945 22049 16957 22083
rect 16991 22049 17003 22083
rect 16945 22043 17003 22049
rect 17313 22083 17371 22089
rect 17313 22049 17325 22083
rect 17359 22080 17371 22083
rect 17494 22080 17500 22092
rect 17359 22052 17500 22080
rect 17359 22049 17371 22052
rect 17313 22043 17371 22049
rect 9548 21984 10456 22012
rect 9548 21972 9554 21984
rect 10502 21972 10508 22024
rect 10560 22012 10566 22024
rect 12161 22015 12219 22021
rect 12161 22012 12173 22015
rect 10560 21984 12173 22012
rect 10560 21972 10566 21984
rect 12161 21981 12173 21984
rect 12207 21981 12219 22015
rect 12161 21975 12219 21981
rect 12250 21972 12256 22024
rect 12308 21972 12314 22024
rect 12618 21972 12624 22024
rect 12676 21972 12682 22024
rect 13814 21972 13820 22024
rect 13872 21972 13878 22024
rect 13998 21972 14004 22024
rect 14056 21972 14062 22024
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 22012 14519 22015
rect 14826 22012 14832 22024
rect 14507 21984 14832 22012
rect 14507 21981 14519 21984
rect 14461 21975 14519 21981
rect 5994 21904 6000 21956
rect 6052 21944 6058 21956
rect 6641 21947 6699 21953
rect 6641 21944 6653 21947
rect 6052 21916 6653 21944
rect 6052 21904 6058 21916
rect 6641 21913 6653 21916
rect 6687 21944 6699 21947
rect 12636 21944 12664 21972
rect 14476 21944 14504 21975
rect 14826 21972 14832 21984
rect 14884 21972 14890 22024
rect 16853 22015 16911 22021
rect 16853 21981 16865 22015
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 6687 21916 12434 21944
rect 12636 21916 14504 21944
rect 16577 21947 16635 21953
rect 6687 21913 6699 21916
rect 6641 21907 6699 21913
rect 4890 21876 4896 21888
rect 4304 21848 4896 21876
rect 4304 21836 4310 21848
rect 4890 21836 4896 21848
rect 4948 21876 4954 21888
rect 6917 21879 6975 21885
rect 6917 21876 6929 21879
rect 4948 21848 6929 21876
rect 4948 21836 4954 21848
rect 6917 21845 6929 21848
rect 6963 21845 6975 21879
rect 6917 21839 6975 21845
rect 9582 21836 9588 21888
rect 9640 21836 9646 21888
rect 10318 21836 10324 21888
rect 10376 21836 10382 21888
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 11514 21876 11520 21888
rect 11204 21848 11520 21876
rect 11204 21836 11210 21848
rect 11514 21836 11520 21848
rect 11572 21836 11578 21888
rect 11609 21879 11667 21885
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11698 21876 11704 21888
rect 11655 21848 11704 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 11885 21879 11943 21885
rect 11885 21845 11897 21879
rect 11931 21876 11943 21879
rect 12066 21876 12072 21888
rect 11931 21848 12072 21876
rect 11931 21845 11943 21848
rect 11885 21839 11943 21845
rect 12066 21836 12072 21848
rect 12124 21836 12130 21888
rect 12406 21876 12434 21916
rect 16577 21913 16589 21947
rect 16623 21944 16635 21947
rect 16868 21944 16896 21975
rect 16623 21916 16896 21944
rect 16960 21944 16988 22043
rect 17494 22040 17500 22052
rect 17552 22040 17558 22092
rect 18874 22040 18880 22092
rect 18932 22040 18938 22092
rect 19245 22083 19303 22089
rect 19245 22049 19257 22083
rect 19291 22049 19303 22083
rect 19245 22043 19303 22049
rect 21913 22083 21971 22089
rect 21913 22049 21925 22083
rect 21959 22080 21971 22083
rect 22296 22080 22324 22188
rect 22646 22176 22652 22188
rect 22704 22176 22710 22228
rect 25130 22216 25136 22228
rect 23216 22188 25136 22216
rect 23216 22157 23244 22188
rect 25130 22176 25136 22188
rect 25188 22176 25194 22228
rect 25225 22219 25283 22225
rect 25225 22185 25237 22219
rect 25271 22185 25283 22219
rect 25225 22179 25283 22185
rect 23201 22151 23259 22157
rect 23201 22148 23213 22151
rect 21959 22052 22324 22080
rect 22388 22120 23213 22148
rect 21959 22049 21971 22052
rect 21913 22043 21971 22049
rect 17221 22015 17279 22021
rect 17221 21981 17233 22015
rect 17267 22012 17279 22015
rect 17402 22012 17408 22024
rect 17267 21984 17408 22012
rect 17267 21981 17279 21984
rect 17221 21975 17279 21981
rect 17402 21972 17408 21984
rect 17460 21972 17466 22024
rect 18966 22012 18972 22024
rect 17512 21984 18972 22012
rect 17512 21944 17540 21984
rect 18966 21972 18972 21984
rect 19024 21972 19030 22024
rect 19058 21972 19064 22024
rect 19116 21972 19122 22024
rect 16960 21916 17540 21944
rect 16623 21913 16635 21916
rect 16577 21907 16635 21913
rect 16592 21876 16620 21907
rect 12406 21848 16620 21876
rect 16666 21836 16672 21888
rect 16724 21836 16730 21888
rect 16868 21876 16896 21916
rect 17586 21904 17592 21956
rect 17644 21944 17650 21956
rect 18141 21947 18199 21953
rect 17644 21916 18092 21944
rect 17644 21904 17650 21916
rect 17862 21876 17868 21888
rect 16868 21848 17868 21876
rect 17862 21836 17868 21848
rect 17920 21836 17926 21888
rect 17954 21836 17960 21888
rect 18012 21836 18018 21888
rect 18064 21876 18092 21916
rect 18141 21913 18153 21947
rect 18187 21944 18199 21947
rect 18690 21944 18696 21956
rect 18187 21916 18696 21944
rect 18187 21913 18199 21916
rect 18141 21907 18199 21913
rect 18690 21904 18696 21916
rect 18748 21944 18754 21956
rect 19260 21944 19288 22043
rect 19610 21972 19616 22024
rect 19668 22012 19674 22024
rect 21726 22012 21732 22024
rect 19668 21984 21732 22012
rect 19668 21972 19674 21984
rect 21726 21972 21732 21984
rect 21784 21972 21790 22024
rect 18748 21916 19288 21944
rect 19429 21947 19487 21953
rect 18748 21904 18754 21916
rect 19429 21913 19441 21947
rect 19475 21944 19487 21947
rect 19475 21916 20484 21944
rect 19475 21913 19487 21916
rect 19429 21907 19487 21913
rect 18230 21876 18236 21888
rect 18064 21848 18236 21876
rect 18230 21836 18236 21848
rect 18288 21836 18294 21888
rect 18414 21836 18420 21888
rect 18472 21876 18478 21888
rect 18509 21879 18567 21885
rect 18509 21876 18521 21879
rect 18472 21848 18521 21876
rect 18472 21836 18478 21848
rect 18509 21845 18521 21848
rect 18555 21845 18567 21879
rect 18509 21839 18567 21845
rect 18782 21836 18788 21888
rect 18840 21836 18846 21888
rect 19702 21836 19708 21888
rect 19760 21876 19766 21888
rect 19797 21879 19855 21885
rect 19797 21876 19809 21879
rect 19760 21848 19809 21876
rect 19760 21836 19766 21848
rect 19797 21845 19809 21848
rect 19843 21845 19855 21879
rect 20456 21876 20484 21916
rect 21910 21876 21916 21888
rect 20456 21848 21916 21876
rect 19797 21839 19855 21845
rect 21910 21836 21916 21848
rect 21968 21836 21974 21888
rect 22002 21836 22008 21888
rect 22060 21836 22066 21888
rect 22186 21836 22192 21888
rect 22244 21876 22250 21888
rect 22388 21885 22416 22120
rect 23201 22117 23213 22120
rect 23247 22117 23259 22151
rect 23201 22111 23259 22117
rect 23290 22108 23296 22160
rect 23348 22148 23354 22160
rect 23348 22120 23520 22148
rect 23348 22108 23354 22120
rect 22922 22040 22928 22092
rect 22980 22040 22986 22092
rect 23492 22089 23520 22120
rect 23842 22108 23848 22160
rect 23900 22148 23906 22160
rect 25240 22148 25268 22179
rect 25406 22176 25412 22228
rect 25464 22216 25470 22228
rect 25501 22219 25559 22225
rect 25501 22216 25513 22219
rect 25464 22188 25513 22216
rect 25464 22176 25470 22188
rect 25501 22185 25513 22188
rect 25547 22185 25559 22219
rect 25501 22179 25559 22185
rect 25958 22176 25964 22228
rect 26016 22176 26022 22228
rect 26326 22176 26332 22228
rect 26384 22176 26390 22228
rect 26418 22176 26424 22228
rect 26476 22216 26482 22228
rect 26513 22219 26571 22225
rect 26513 22216 26525 22219
rect 26476 22188 26525 22216
rect 26476 22176 26482 22188
rect 26513 22185 26525 22188
rect 26559 22185 26571 22219
rect 26513 22179 26571 22185
rect 26694 22176 26700 22228
rect 26752 22216 26758 22228
rect 27249 22219 27307 22225
rect 27249 22216 27261 22219
rect 26752 22188 27261 22216
rect 26752 22176 26758 22188
rect 27249 22185 27261 22188
rect 27295 22216 27307 22219
rect 27430 22216 27436 22228
rect 27295 22188 27436 22216
rect 27295 22185 27307 22188
rect 27249 22179 27307 22185
rect 27430 22176 27436 22188
rect 27488 22216 27494 22228
rect 27488 22188 28580 22216
rect 27488 22176 27494 22188
rect 25976 22148 26004 22176
rect 23900 22120 24242 22148
rect 25240 22120 26004 22148
rect 26344 22148 26372 22176
rect 26881 22151 26939 22157
rect 26881 22148 26893 22151
rect 26344 22120 26893 22148
rect 23900 22108 23906 22120
rect 26881 22117 26893 22120
rect 26927 22117 26939 22151
rect 27614 22148 27620 22160
rect 26881 22111 26939 22117
rect 26988 22120 27620 22148
rect 23477 22083 23535 22089
rect 23477 22049 23489 22083
rect 23523 22049 23535 22083
rect 23477 22043 23535 22049
rect 25593 22083 25651 22089
rect 25593 22049 25605 22083
rect 25639 22080 25651 22083
rect 26513 22083 26571 22089
rect 25639 22052 25728 22080
rect 25639 22049 25651 22052
rect 25593 22043 25651 22049
rect 25700 22024 25728 22052
rect 26513 22049 26525 22083
rect 26559 22049 26571 22083
rect 26513 22043 26571 22049
rect 26605 22083 26663 22089
rect 26605 22049 26617 22083
rect 26651 22080 26663 22083
rect 26694 22080 26700 22092
rect 26651 22052 26700 22080
rect 26651 22049 26663 22052
rect 26605 22043 26663 22049
rect 22738 21972 22744 22024
rect 22796 22012 22802 22024
rect 22833 22015 22891 22021
rect 22833 22012 22845 22015
rect 22796 21984 22845 22012
rect 22796 21972 22802 21984
rect 22833 21981 22845 21984
rect 22879 21981 22891 22015
rect 22833 21975 22891 21981
rect 23198 21972 23204 22024
rect 23256 22012 23262 22024
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 23256 21984 23305 22012
rect 23256 21972 23262 21984
rect 23293 21981 23305 21984
rect 23339 21981 23351 22015
rect 23753 22015 23811 22021
rect 23753 22012 23765 22015
rect 23293 21975 23351 21981
rect 23584 21984 23765 22012
rect 22649 21947 22707 21953
rect 22649 21913 22661 21947
rect 22695 21944 22707 21947
rect 23584 21944 23612 21984
rect 23753 21981 23765 21984
rect 23799 21981 23811 22015
rect 23753 21975 23811 21981
rect 25682 21972 25688 22024
rect 25740 21972 25746 22024
rect 22695 21916 23612 21944
rect 26528 21944 26556 22043
rect 26694 22040 26700 22052
rect 26752 22040 26758 22092
rect 26789 22083 26847 22089
rect 26789 22049 26801 22083
rect 26835 22080 26847 22083
rect 26988 22080 27016 22120
rect 26835 22052 27016 22080
rect 26835 22049 26847 22052
rect 26789 22043 26847 22049
rect 26988 22012 27016 22052
rect 27062 22040 27068 22092
rect 27120 22080 27126 22092
rect 27356 22089 27384 22120
rect 27614 22108 27620 22120
rect 27672 22108 27678 22160
rect 28552 22148 28580 22188
rect 31570 22176 31576 22228
rect 31628 22216 31634 22228
rect 31849 22219 31907 22225
rect 31849 22216 31861 22219
rect 31628 22188 31861 22216
rect 31628 22176 31634 22188
rect 31849 22185 31861 22188
rect 31895 22185 31907 22219
rect 31849 22179 31907 22185
rect 32217 22219 32275 22225
rect 32217 22185 32229 22219
rect 32263 22216 32275 22219
rect 32766 22216 32772 22228
rect 32263 22188 32772 22216
rect 32263 22185 32275 22188
rect 32217 22179 32275 22185
rect 32766 22176 32772 22188
rect 32824 22176 32830 22228
rect 27908 22120 28304 22148
rect 28552 22120 28672 22148
rect 27908 22092 27936 22120
rect 27341 22083 27399 22089
rect 27120 22052 27292 22080
rect 27120 22040 27126 22052
rect 27264 22012 27292 22052
rect 27341 22049 27353 22083
rect 27387 22049 27399 22083
rect 27341 22043 27399 22049
rect 27801 22083 27859 22089
rect 27801 22049 27813 22083
rect 27847 22080 27859 22083
rect 27890 22080 27896 22092
rect 27847 22052 27896 22080
rect 27847 22049 27859 22052
rect 27801 22043 27859 22049
rect 27890 22040 27896 22052
rect 27948 22040 27954 22092
rect 28169 22083 28227 22089
rect 28169 22080 28181 22083
rect 28000 22052 28181 22080
rect 28000 22012 28028 22052
rect 28169 22049 28181 22052
rect 28215 22049 28227 22083
rect 28276 22080 28304 22120
rect 28644 22089 28672 22120
rect 29270 22108 29276 22160
rect 29328 22148 29334 22160
rect 30377 22151 30435 22157
rect 30377 22148 30389 22151
rect 29328 22120 30389 22148
rect 29328 22108 29334 22120
rect 28629 22083 28687 22089
rect 28276 22052 28396 22080
rect 28169 22043 28227 22049
rect 26988 21984 27108 22012
rect 27264 21984 28028 22012
rect 27080 21956 27108 21984
rect 28074 21972 28080 22024
rect 28132 22012 28138 22024
rect 28261 22015 28319 22021
rect 28261 22012 28273 22015
rect 28132 21984 28273 22012
rect 28132 21972 28138 21984
rect 28261 21981 28273 21984
rect 28307 21981 28319 22015
rect 28368 22012 28396 22052
rect 28629 22049 28641 22083
rect 28675 22049 28687 22083
rect 28629 22043 28687 22049
rect 28905 22083 28963 22089
rect 28905 22049 28917 22083
rect 28951 22080 28963 22083
rect 29086 22080 29092 22092
rect 28951 22052 29092 22080
rect 28951 22049 28963 22052
rect 28905 22043 28963 22049
rect 29086 22040 29092 22052
rect 29144 22040 29150 22092
rect 29380 22080 29408 22120
rect 30377 22117 30389 22120
rect 30423 22117 30435 22151
rect 30377 22111 30435 22117
rect 30650 22108 30656 22160
rect 30708 22148 30714 22160
rect 30708 22120 31892 22148
rect 30708 22108 30714 22120
rect 29457 22083 29515 22089
rect 29457 22080 29469 22083
rect 29380 22052 29469 22080
rect 29457 22049 29469 22052
rect 29503 22049 29515 22083
rect 29457 22043 29515 22049
rect 29546 22040 29552 22092
rect 29604 22040 29610 22092
rect 31864 22080 31892 22120
rect 31938 22108 31944 22160
rect 31996 22148 32002 22160
rect 32369 22151 32427 22157
rect 32369 22148 32381 22151
rect 31996 22120 32381 22148
rect 31996 22108 32002 22120
rect 32369 22117 32381 22120
rect 32415 22117 32427 22151
rect 32585 22151 32643 22157
rect 32585 22148 32597 22151
rect 32369 22111 32427 22117
rect 32508 22120 32597 22148
rect 32508 22080 32536 22120
rect 32585 22117 32597 22120
rect 32631 22117 32643 22151
rect 32585 22111 32643 22117
rect 31864 22052 32536 22080
rect 28721 22015 28779 22021
rect 28721 22012 28733 22015
rect 28368 21984 28733 22012
rect 28261 21975 28319 21981
rect 28721 21981 28733 21984
rect 28767 21981 28779 22015
rect 28721 21975 28779 21981
rect 30098 21972 30104 22024
rect 30156 21972 30162 22024
rect 26970 21944 26976 21956
rect 26528 21916 26976 21944
rect 22695 21913 22707 21916
rect 22649 21907 22707 21913
rect 26970 21904 26976 21916
rect 27028 21904 27034 21956
rect 27062 21904 27068 21956
rect 27120 21904 27126 21956
rect 28920 21916 30604 21944
rect 22373 21879 22431 21885
rect 22373 21876 22385 21879
rect 22244 21848 22385 21876
rect 22244 21836 22250 21848
rect 22373 21845 22385 21848
rect 22419 21845 22431 21879
rect 22373 21839 22431 21845
rect 22554 21836 22560 21888
rect 22612 21876 22618 21888
rect 22738 21876 22744 21888
rect 22612 21848 22744 21876
rect 22612 21836 22618 21848
rect 22738 21836 22744 21848
rect 22796 21836 22802 21888
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 24118 21876 24124 21888
rect 23348 21848 24124 21876
rect 23348 21836 23354 21848
rect 24118 21836 24124 21848
rect 24176 21836 24182 21888
rect 27614 21836 27620 21888
rect 27672 21836 27678 21888
rect 27893 21879 27951 21885
rect 27893 21845 27905 21879
rect 27939 21876 27951 21879
rect 28166 21876 28172 21888
rect 27939 21848 28172 21876
rect 27939 21845 27951 21848
rect 27893 21839 27951 21845
rect 28166 21836 28172 21848
rect 28224 21836 28230 21888
rect 28920 21885 28948 21916
rect 30576 21888 30604 21916
rect 28905 21879 28963 21885
rect 28905 21845 28917 21879
rect 28951 21845 28963 21879
rect 28905 21839 28963 21845
rect 28994 21836 29000 21888
rect 29052 21876 29058 21888
rect 29089 21879 29147 21885
rect 29089 21876 29101 21879
rect 29052 21848 29101 21876
rect 29052 21836 29058 21848
rect 29089 21845 29101 21848
rect 29135 21845 29147 21879
rect 29089 21839 29147 21845
rect 30558 21836 30564 21888
rect 30616 21836 30622 21888
rect 32398 21836 32404 21888
rect 32456 21836 32462 21888
rect 2760 21786 34316 21808
rect 2760 21734 6550 21786
rect 6602 21734 6614 21786
rect 6666 21734 6678 21786
rect 6730 21734 6742 21786
rect 6794 21734 6806 21786
rect 6858 21734 14439 21786
rect 14491 21734 14503 21786
rect 14555 21734 14567 21786
rect 14619 21734 14631 21786
rect 14683 21734 14695 21786
rect 14747 21734 22328 21786
rect 22380 21734 22392 21786
rect 22444 21734 22456 21786
rect 22508 21734 22520 21786
rect 22572 21734 22584 21786
rect 22636 21734 30217 21786
rect 30269 21734 30281 21786
rect 30333 21734 30345 21786
rect 30397 21734 30409 21786
rect 30461 21734 30473 21786
rect 30525 21734 34316 21786
rect 2760 21712 34316 21734
rect 4522 21632 4528 21684
rect 4580 21672 4586 21684
rect 5445 21675 5503 21681
rect 5445 21672 5457 21675
rect 4580 21644 5457 21672
rect 4580 21632 4586 21644
rect 5445 21641 5457 21644
rect 5491 21641 5503 21675
rect 5810 21672 5816 21684
rect 5445 21635 5503 21641
rect 5552 21644 5816 21672
rect 5261 21607 5319 21613
rect 5261 21573 5273 21607
rect 5307 21604 5319 21607
rect 5552 21604 5580 21644
rect 5810 21632 5816 21644
rect 5868 21632 5874 21684
rect 7837 21675 7895 21681
rect 7837 21641 7849 21675
rect 7883 21672 7895 21675
rect 8018 21672 8024 21684
rect 7883 21644 8024 21672
rect 7883 21641 7895 21644
rect 7837 21635 7895 21641
rect 8018 21632 8024 21644
rect 8076 21632 8082 21684
rect 9674 21632 9680 21684
rect 9732 21672 9738 21684
rect 9861 21675 9919 21681
rect 9861 21672 9873 21675
rect 9732 21644 9873 21672
rect 9732 21632 9738 21644
rect 9861 21641 9873 21644
rect 9907 21672 9919 21675
rect 10502 21672 10508 21684
rect 9907 21644 10508 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 10502 21632 10508 21644
rect 10560 21632 10566 21684
rect 12342 21632 12348 21684
rect 12400 21672 12406 21684
rect 14001 21675 14059 21681
rect 12400 21644 13952 21672
rect 12400 21632 12406 21644
rect 5307 21576 5580 21604
rect 5307 21573 5319 21576
rect 5261 21567 5319 21573
rect 6914 21564 6920 21616
rect 6972 21604 6978 21616
rect 12250 21604 12256 21616
rect 6972 21576 12256 21604
rect 6972 21564 6978 21576
rect 12250 21564 12256 21576
rect 12308 21564 12314 21616
rect 13924 21604 13952 21644
rect 14001 21641 14013 21675
rect 14047 21672 14059 21675
rect 14366 21672 14372 21684
rect 14047 21644 14372 21672
rect 14047 21641 14059 21644
rect 14001 21635 14059 21641
rect 14366 21632 14372 21644
rect 14424 21632 14430 21684
rect 15010 21632 15016 21684
rect 15068 21672 15074 21684
rect 15105 21675 15163 21681
rect 15105 21672 15117 21675
rect 15068 21644 15117 21672
rect 15068 21632 15074 21644
rect 15105 21641 15117 21644
rect 15151 21641 15163 21675
rect 15105 21635 15163 21641
rect 15838 21632 15844 21684
rect 15896 21632 15902 21684
rect 18138 21632 18144 21684
rect 18196 21632 18202 21684
rect 21358 21672 21364 21684
rect 18248 21644 21364 21672
rect 13924 21576 14688 21604
rect 14660 21548 14688 21576
rect 17862 21564 17868 21616
rect 17920 21604 17926 21616
rect 18248 21604 18276 21644
rect 21358 21632 21364 21644
rect 21416 21632 21422 21684
rect 23382 21632 23388 21684
rect 23440 21672 23446 21684
rect 23477 21675 23535 21681
rect 23477 21672 23489 21675
rect 23440 21644 23489 21672
rect 23440 21632 23446 21644
rect 23477 21641 23489 21644
rect 23523 21672 23535 21675
rect 29270 21672 29276 21684
rect 23523 21644 29276 21672
rect 23523 21641 23535 21644
rect 23477 21635 23535 21641
rect 17920 21576 18276 21604
rect 19429 21607 19487 21613
rect 17920 21564 17926 21576
rect 19429 21573 19441 21607
rect 19475 21604 19487 21607
rect 19518 21604 19524 21616
rect 19475 21576 19524 21604
rect 19475 21573 19487 21576
rect 19429 21567 19487 21573
rect 19518 21564 19524 21576
rect 19576 21564 19582 21616
rect 22554 21564 22560 21616
rect 22612 21604 22618 21616
rect 22922 21604 22928 21616
rect 22612 21576 22928 21604
rect 22612 21564 22618 21576
rect 22922 21564 22928 21576
rect 22980 21564 22986 21616
rect 5629 21539 5687 21545
rect 5629 21505 5641 21539
rect 5675 21536 5687 21539
rect 5994 21536 6000 21548
rect 5675 21508 6000 21536
rect 5675 21505 5687 21508
rect 5629 21499 5687 21505
rect 5994 21496 6000 21508
rect 6052 21496 6058 21548
rect 6086 21496 6092 21548
rect 6144 21496 6150 21548
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21536 6791 21539
rect 9858 21536 9864 21548
rect 6779 21508 9864 21536
rect 6779 21505 6791 21508
rect 6733 21499 6791 21505
rect 4798 21428 4804 21480
rect 4856 21428 4862 21480
rect 5721 21471 5779 21477
rect 5721 21468 5733 21471
rect 5644 21440 5733 21468
rect 3234 21360 3240 21412
rect 3292 21400 3298 21412
rect 3292 21372 3358 21400
rect 3292 21360 3298 21372
rect 4522 21360 4528 21412
rect 4580 21360 4586 21412
rect 5644 21344 5672 21440
rect 5721 21437 5733 21440
rect 5767 21468 5779 21471
rect 6181 21471 6239 21477
rect 6181 21468 6193 21471
rect 5767 21440 6193 21468
rect 5767 21437 5779 21440
rect 5721 21431 5779 21437
rect 6181 21437 6193 21440
rect 6227 21437 6239 21471
rect 6181 21431 6239 21437
rect 6365 21471 6423 21477
rect 6365 21437 6377 21471
rect 6411 21468 6423 21471
rect 6748 21468 6776 21499
rect 9858 21496 9864 21508
rect 9916 21496 9922 21548
rect 10594 21536 10600 21548
rect 10060 21508 10600 21536
rect 6411 21440 6776 21468
rect 9585 21471 9643 21477
rect 6411 21437 6423 21440
rect 6365 21431 6423 21437
rect 9585 21437 9597 21471
rect 9631 21468 9643 21471
rect 10060 21468 10088 21508
rect 10594 21496 10600 21508
rect 10652 21496 10658 21548
rect 11333 21539 11391 21545
rect 11333 21505 11345 21539
rect 11379 21536 11391 21539
rect 12066 21536 12072 21548
rect 11379 21508 12072 21536
rect 11379 21505 11391 21508
rect 11333 21499 11391 21505
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 12618 21536 12624 21548
rect 12268 21508 12624 21536
rect 9631 21440 10088 21468
rect 9631 21437 9643 21440
rect 9585 21431 9643 21437
rect 10134 21428 10140 21480
rect 10192 21468 10198 21480
rect 11425 21471 11483 21477
rect 11425 21468 11437 21471
rect 10192 21440 11437 21468
rect 10192 21428 10198 21440
rect 11425 21437 11437 21440
rect 11471 21437 11483 21471
rect 11425 21431 11483 21437
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 5997 21403 6055 21409
rect 5997 21400 6009 21403
rect 5920 21372 6009 21400
rect 3053 21335 3111 21341
rect 3053 21301 3065 21335
rect 3099 21332 3111 21335
rect 4338 21332 4344 21344
rect 3099 21304 4344 21332
rect 3099 21301 3111 21304
rect 3053 21295 3111 21301
rect 4338 21292 4344 21304
rect 4396 21292 4402 21344
rect 5626 21292 5632 21344
rect 5684 21292 5690 21344
rect 5920 21332 5948 21372
rect 5997 21369 6009 21372
rect 6043 21369 6055 21403
rect 5997 21363 6055 21369
rect 6086 21360 6092 21412
rect 6144 21400 6150 21412
rect 6273 21403 6331 21409
rect 6273 21400 6285 21403
rect 6144 21372 6285 21400
rect 6144 21360 6150 21372
rect 6273 21369 6285 21372
rect 6319 21400 6331 21403
rect 7650 21400 7656 21412
rect 6319 21372 7656 21400
rect 6319 21369 6331 21372
rect 6273 21363 6331 21369
rect 7650 21360 7656 21372
rect 7708 21360 7714 21412
rect 9122 21360 9128 21412
rect 9180 21360 9186 21412
rect 9766 21360 9772 21412
rect 9824 21400 9830 21412
rect 11330 21400 11336 21412
rect 9824 21372 11336 21400
rect 9824 21360 9830 21372
rect 11330 21360 11336 21372
rect 11388 21360 11394 21412
rect 11532 21400 11560 21431
rect 11606 21428 11612 21480
rect 11664 21428 11670 21480
rect 11698 21428 11704 21480
rect 11756 21468 11762 21480
rect 12268 21477 12296 21508
rect 12618 21496 12624 21508
rect 12676 21496 12682 21548
rect 13998 21536 14004 21548
rect 13648 21508 14004 21536
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 11756 21440 12265 21468
rect 11756 21428 11762 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 13648 21454 13676 21508
rect 13998 21496 14004 21508
rect 14056 21496 14062 21548
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14461 21539 14519 21545
rect 14461 21536 14473 21539
rect 14240 21508 14473 21536
rect 14240 21496 14246 21508
rect 14461 21505 14473 21508
rect 14507 21505 14519 21539
rect 14461 21499 14519 21505
rect 14642 21496 14648 21548
rect 14700 21496 14706 21548
rect 14918 21496 14924 21548
rect 14976 21536 14982 21548
rect 16393 21539 16451 21545
rect 16393 21536 16405 21539
rect 14976 21508 16405 21536
rect 14976 21496 14982 21508
rect 16393 21505 16405 21508
rect 16439 21505 16451 21539
rect 16393 21499 16451 21505
rect 16666 21496 16672 21548
rect 16724 21496 16730 21548
rect 17126 21496 17132 21548
rect 17184 21536 17190 21548
rect 22741 21539 22799 21545
rect 17184 21508 19380 21536
rect 17184 21496 17190 21508
rect 12253 21431 12311 21437
rect 13906 21428 13912 21480
rect 13964 21468 13970 21480
rect 14200 21468 14228 21496
rect 13964 21440 14228 21468
rect 15933 21471 15991 21477
rect 13964 21428 13970 21440
rect 15933 21437 15945 21471
rect 15979 21437 15991 21471
rect 18782 21468 18788 21480
rect 17802 21440 18788 21468
rect 15933 21431 15991 21437
rect 12529 21403 12587 21409
rect 12529 21400 12541 21403
rect 11532 21372 11652 21400
rect 6178 21332 6184 21344
rect 5920 21304 6184 21332
rect 6178 21292 6184 21304
rect 6236 21332 6242 21344
rect 7006 21332 7012 21344
rect 6236 21304 7012 21332
rect 6236 21292 6242 21304
rect 7006 21292 7012 21304
rect 7064 21332 7070 21344
rect 7101 21335 7159 21341
rect 7101 21332 7113 21335
rect 7064 21304 7113 21332
rect 7064 21292 7070 21304
rect 7101 21301 7113 21304
rect 7147 21332 7159 21335
rect 7834 21332 7840 21344
rect 7147 21304 7840 21332
rect 7147 21301 7159 21304
rect 7101 21295 7159 21301
rect 7834 21292 7840 21304
rect 7892 21292 7898 21344
rect 9140 21332 9168 21360
rect 11624 21344 11652 21372
rect 11808 21372 12541 21400
rect 9493 21335 9551 21341
rect 9493 21332 9505 21335
rect 9140 21304 9505 21332
rect 9493 21301 9505 21304
rect 9539 21332 9551 21335
rect 11054 21332 11060 21344
rect 9539 21304 11060 21332
rect 9539 21301 9551 21304
rect 9493 21295 9551 21301
rect 11054 21292 11060 21304
rect 11112 21292 11118 21344
rect 11606 21292 11612 21344
rect 11664 21292 11670 21344
rect 11808 21341 11836 21372
rect 12529 21369 12541 21372
rect 12575 21369 12587 21403
rect 15948 21400 15976 21431
rect 18782 21428 18788 21440
rect 18840 21428 18846 21480
rect 18966 21428 18972 21480
rect 19024 21468 19030 21480
rect 19352 21478 19380 21508
rect 22741 21505 22753 21539
rect 22787 21536 22799 21539
rect 23474 21536 23480 21548
rect 22787 21508 23480 21536
rect 22787 21505 22799 21508
rect 22741 21499 22799 21505
rect 23474 21496 23480 21508
rect 23532 21496 23538 21548
rect 19352 21477 19472 21478
rect 19153 21471 19211 21477
rect 19153 21468 19165 21471
rect 19024 21440 19165 21468
rect 19024 21428 19030 21440
rect 19153 21437 19165 21440
rect 19199 21437 19211 21471
rect 19352 21471 19487 21477
rect 19352 21450 19441 21471
rect 19153 21431 19211 21437
rect 19429 21437 19441 21450
rect 19475 21468 19487 21471
rect 19475 21440 19932 21468
rect 19475 21437 19487 21440
rect 19429 21431 19487 21437
rect 16758 21400 16764 21412
rect 15948 21372 16764 21400
rect 12529 21363 12587 21369
rect 16758 21360 16764 21372
rect 16816 21360 16822 21412
rect 18708 21372 19564 21400
rect 11793 21335 11851 21341
rect 11793 21301 11805 21335
rect 11839 21301 11851 21335
rect 11793 21295 11851 21301
rect 12250 21292 12256 21344
rect 12308 21332 12314 21344
rect 14737 21335 14795 21341
rect 14737 21332 14749 21335
rect 12308 21304 14749 21332
rect 12308 21292 12314 21304
rect 14737 21301 14749 21304
rect 14783 21332 14795 21335
rect 15010 21332 15016 21344
rect 14783 21304 15016 21332
rect 14783 21301 14795 21304
rect 14737 21295 14795 21301
rect 15010 21292 15016 21304
rect 15068 21332 15074 21344
rect 15381 21335 15439 21341
rect 15381 21332 15393 21335
rect 15068 21304 15393 21332
rect 15068 21292 15074 21304
rect 15381 21301 15393 21304
rect 15427 21332 15439 21335
rect 15654 21332 15660 21344
rect 15427 21304 15660 21332
rect 15427 21301 15439 21304
rect 15381 21295 15439 21301
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 16666 21292 16672 21344
rect 16724 21332 16730 21344
rect 18708 21332 18736 21372
rect 19536 21344 19564 21372
rect 16724 21304 18736 21332
rect 16724 21292 16730 21304
rect 18782 21292 18788 21344
rect 18840 21332 18846 21344
rect 18877 21335 18935 21341
rect 18877 21332 18889 21335
rect 18840 21304 18889 21332
rect 18840 21292 18846 21304
rect 18877 21301 18889 21304
rect 18923 21332 18935 21335
rect 19058 21332 19064 21344
rect 18923 21304 19064 21332
rect 18923 21301 18935 21304
rect 18877 21295 18935 21301
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 19518 21292 19524 21344
rect 19576 21292 19582 21344
rect 19904 21341 19932 21440
rect 20990 21428 20996 21480
rect 21048 21428 21054 21480
rect 23584 21477 23612 21644
rect 29270 21632 29276 21644
rect 29328 21632 29334 21684
rect 29457 21675 29515 21681
rect 29457 21641 29469 21675
rect 29503 21672 29515 21675
rect 30098 21672 30104 21684
rect 29503 21644 30104 21672
rect 29503 21641 29515 21644
rect 29457 21635 29515 21641
rect 30098 21632 30104 21644
rect 30156 21632 30162 21684
rect 31573 21675 31631 21681
rect 31573 21641 31585 21675
rect 31619 21672 31631 21675
rect 31938 21672 31944 21684
rect 31619 21644 31944 21672
rect 31619 21641 31631 21644
rect 31573 21635 31631 21641
rect 31938 21632 31944 21644
rect 31996 21632 32002 21684
rect 32398 21632 32404 21684
rect 32456 21632 32462 21684
rect 24026 21564 24032 21616
rect 24084 21604 24090 21616
rect 24857 21607 24915 21613
rect 24857 21604 24869 21607
rect 24084 21576 24869 21604
rect 24084 21564 24090 21576
rect 24857 21573 24869 21576
rect 24903 21573 24915 21607
rect 24857 21567 24915 21573
rect 26050 21496 26056 21548
rect 26108 21496 26114 21548
rect 29638 21496 29644 21548
rect 29696 21496 29702 21548
rect 29917 21539 29975 21545
rect 29917 21505 29929 21539
rect 29963 21536 29975 21539
rect 30193 21539 30251 21545
rect 30193 21536 30205 21539
rect 29963 21508 30205 21536
rect 29963 21505 29975 21508
rect 29917 21499 29975 21505
rect 30193 21505 30205 21508
rect 30239 21505 30251 21539
rect 32416 21536 32444 21632
rect 30193 21499 30251 21505
rect 30300 21508 32444 21536
rect 23569 21471 23627 21477
rect 23569 21437 23581 21471
rect 23615 21437 23627 21471
rect 23569 21431 23627 21437
rect 23750 21428 23756 21480
rect 23808 21468 23814 21480
rect 25685 21471 25743 21477
rect 23808 21440 25360 21468
rect 23808 21428 23814 21440
rect 21266 21360 21272 21412
rect 21324 21360 21330 21412
rect 22002 21360 22008 21412
rect 22060 21360 22066 21412
rect 19889 21335 19947 21341
rect 19889 21301 19901 21335
rect 19935 21332 19947 21335
rect 20622 21332 20628 21344
rect 19935 21304 20628 21332
rect 19935 21301 19947 21304
rect 19889 21295 19947 21301
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 22646 21292 22652 21344
rect 22704 21332 22710 21344
rect 23017 21335 23075 21341
rect 23017 21332 23029 21335
rect 22704 21304 23029 21332
rect 22704 21292 22710 21304
rect 23017 21301 23029 21304
rect 23063 21301 23075 21335
rect 25332 21332 25360 21440
rect 25685 21437 25697 21471
rect 25731 21468 25743 21471
rect 25774 21468 25780 21480
rect 25731 21440 25780 21468
rect 25731 21437 25743 21440
rect 25685 21431 25743 21437
rect 25774 21428 25780 21440
rect 25832 21428 25838 21480
rect 25869 21471 25927 21477
rect 25869 21437 25881 21471
rect 25915 21468 25927 21471
rect 26142 21468 26148 21480
rect 25915 21440 26148 21468
rect 25915 21437 25927 21440
rect 25869 21431 25927 21437
rect 26142 21428 26148 21440
rect 26200 21428 26206 21480
rect 26605 21471 26663 21477
rect 26605 21468 26617 21471
rect 26344 21440 26617 21468
rect 25685 21335 25743 21341
rect 25685 21332 25697 21335
rect 25332 21304 25697 21332
rect 23017 21295 23075 21301
rect 25685 21301 25697 21304
rect 25731 21332 25743 21335
rect 26344 21332 26372 21440
rect 26605 21437 26617 21440
rect 26651 21437 26663 21471
rect 26605 21431 26663 21437
rect 28166 21428 28172 21480
rect 28224 21468 28230 21480
rect 29733 21471 29791 21477
rect 29733 21468 29745 21471
rect 28224 21440 29745 21468
rect 28224 21428 28230 21440
rect 29733 21437 29745 21440
rect 29779 21437 29791 21471
rect 29733 21431 29791 21437
rect 29822 21428 29828 21480
rect 29880 21468 29886 21480
rect 30300 21477 30328 21508
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29880 21440 30113 21468
rect 29880 21428 29886 21440
rect 30101 21437 30113 21440
rect 30147 21437 30159 21471
rect 30101 21431 30159 21437
rect 30285 21471 30343 21477
rect 30285 21437 30297 21471
rect 30331 21437 30343 21471
rect 30285 21431 30343 21437
rect 26510 21360 26516 21412
rect 26568 21400 26574 21412
rect 28184 21400 28212 21428
rect 26568 21372 28212 21400
rect 30116 21400 30144 21431
rect 30650 21428 30656 21480
rect 30708 21428 30714 21480
rect 31021 21471 31079 21477
rect 31021 21437 31033 21471
rect 31067 21468 31079 21471
rect 31110 21468 31116 21480
rect 31067 21440 31116 21468
rect 31067 21437 31079 21440
rect 31021 21431 31079 21437
rect 31110 21428 31116 21440
rect 31168 21428 31174 21480
rect 31665 21471 31723 21477
rect 31665 21468 31677 21471
rect 31312 21440 31677 21468
rect 30668 21400 30696 21428
rect 31312 21412 31340 21440
rect 31665 21437 31677 21440
rect 31711 21437 31723 21471
rect 31665 21431 31723 21437
rect 31849 21471 31907 21477
rect 31849 21437 31861 21471
rect 31895 21437 31907 21471
rect 31849 21431 31907 21437
rect 30116 21372 30696 21400
rect 31205 21403 31263 21409
rect 26568 21360 26574 21372
rect 31205 21369 31217 21403
rect 31251 21400 31263 21403
rect 31294 21400 31300 21412
rect 31251 21372 31300 21400
rect 31251 21369 31263 21372
rect 31205 21363 31263 21369
rect 31294 21360 31300 21372
rect 31352 21360 31358 21412
rect 31389 21403 31447 21409
rect 31389 21369 31401 21403
rect 31435 21400 31447 21403
rect 31864 21400 31892 21431
rect 31435 21372 31892 21400
rect 31435 21369 31447 21372
rect 31389 21363 31447 21369
rect 25731 21304 26372 21332
rect 25731 21301 25743 21304
rect 25685 21295 25743 21301
rect 29454 21292 29460 21344
rect 29512 21332 29518 21344
rect 30377 21335 30435 21341
rect 30377 21332 30389 21335
rect 29512 21304 30389 21332
rect 29512 21292 29518 21304
rect 30377 21301 30389 21304
rect 30423 21332 30435 21335
rect 31404 21332 31432 21363
rect 30423 21304 31432 21332
rect 31849 21335 31907 21341
rect 30423 21301 30435 21304
rect 30377 21295 30435 21301
rect 31849 21301 31861 21335
rect 31895 21332 31907 21335
rect 31956 21332 31984 21508
rect 32582 21428 32588 21480
rect 32640 21428 32646 21480
rect 33781 21403 33839 21409
rect 33781 21369 33793 21403
rect 33827 21400 33839 21403
rect 34882 21400 34888 21412
rect 33827 21372 34888 21400
rect 33827 21369 33839 21372
rect 33781 21363 33839 21369
rect 34882 21360 34888 21372
rect 34940 21360 34946 21412
rect 31895 21304 31984 21332
rect 31895 21301 31907 21304
rect 31849 21295 31907 21301
rect 2760 21242 34316 21264
rect 2760 21190 7210 21242
rect 7262 21190 7274 21242
rect 7326 21190 7338 21242
rect 7390 21190 7402 21242
rect 7454 21190 7466 21242
rect 7518 21190 15099 21242
rect 15151 21190 15163 21242
rect 15215 21190 15227 21242
rect 15279 21190 15291 21242
rect 15343 21190 15355 21242
rect 15407 21190 22988 21242
rect 23040 21190 23052 21242
rect 23104 21190 23116 21242
rect 23168 21190 23180 21242
rect 23232 21190 23244 21242
rect 23296 21190 30877 21242
rect 30929 21190 30941 21242
rect 30993 21190 31005 21242
rect 31057 21190 31069 21242
rect 31121 21190 31133 21242
rect 31185 21190 34316 21242
rect 2760 21168 34316 21190
rect 4522 21088 4528 21140
rect 4580 21128 4586 21140
rect 4617 21131 4675 21137
rect 4617 21128 4629 21131
rect 4580 21100 4629 21128
rect 4580 21088 4586 21100
rect 4617 21097 4629 21100
rect 4663 21097 4675 21131
rect 6086 21128 6092 21140
rect 4617 21091 4675 21097
rect 5736 21100 6092 21128
rect 1302 21020 1308 21072
rect 1360 21060 1366 21072
rect 3237 21063 3295 21069
rect 3237 21060 3249 21063
rect 1360 21032 3249 21060
rect 1360 21020 1366 21032
rect 3237 21029 3249 21032
rect 3283 21029 3295 21063
rect 3237 21023 3295 21029
rect 5166 21020 5172 21072
rect 5224 21060 5230 21072
rect 5736 21069 5764 21100
rect 6086 21088 6092 21100
rect 6144 21088 6150 21140
rect 6196 21100 8064 21128
rect 5629 21063 5687 21069
rect 5629 21060 5641 21063
rect 5224 21032 5641 21060
rect 5224 21020 5230 21032
rect 5629 21029 5641 21032
rect 5675 21029 5687 21063
rect 5629 21023 5687 21029
rect 5721 21063 5779 21069
rect 5721 21029 5733 21063
rect 5767 21029 5779 21063
rect 6196 21060 6224 21100
rect 8036 21072 8064 21100
rect 8110 21088 8116 21140
rect 8168 21088 8174 21140
rect 9582 21088 9588 21140
rect 9640 21088 9646 21140
rect 10870 21088 10876 21140
rect 10928 21128 10934 21140
rect 10965 21131 11023 21137
rect 10965 21128 10977 21131
rect 10928 21100 10977 21128
rect 10928 21088 10934 21100
rect 10965 21097 10977 21100
rect 11011 21128 11023 21131
rect 13541 21131 13599 21137
rect 11011 21100 11100 21128
rect 11011 21097 11023 21100
rect 10965 21091 11023 21097
rect 5721 21023 5779 21029
rect 6104 21032 6224 21060
rect 4430 20952 4436 21004
rect 4488 20952 4494 21004
rect 5534 20952 5540 21004
rect 5592 20952 5598 21004
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 6104 21001 6132 21032
rect 8018 21020 8024 21072
rect 8076 21020 8082 21072
rect 8128 21060 8156 21088
rect 9493 21063 9551 21069
rect 8128 21032 8984 21060
rect 8956 21001 8984 21032
rect 9493 21029 9505 21063
rect 9539 21060 9551 21063
rect 9600 21060 9628 21088
rect 9539 21032 9628 21060
rect 11072 21060 11100 21100
rect 13541 21097 13553 21131
rect 13587 21128 13599 21131
rect 14182 21128 14188 21140
rect 13587 21100 14188 21128
rect 13587 21097 13599 21100
rect 13541 21091 13599 21097
rect 14182 21088 14188 21100
rect 14240 21128 14246 21140
rect 15470 21128 15476 21140
rect 14240 21100 15476 21128
rect 14240 21088 14246 21100
rect 15470 21088 15476 21100
rect 15528 21088 15534 21140
rect 17773 21131 17831 21137
rect 17773 21097 17785 21131
rect 17819 21128 17831 21131
rect 17954 21128 17960 21140
rect 17819 21100 17960 21128
rect 17819 21097 17831 21100
rect 17773 21091 17831 21097
rect 17954 21088 17960 21100
rect 18012 21088 18018 21140
rect 19610 21128 19616 21140
rect 18340 21100 19616 21128
rect 11514 21060 11520 21072
rect 11072 21032 11520 21060
rect 9539 21029 9551 21032
rect 9493 21023 9551 21029
rect 11514 21020 11520 21032
rect 11572 21020 11578 21072
rect 11606 21020 11612 21072
rect 11664 21060 11670 21072
rect 11664 21032 12296 21060
rect 11664 21020 11670 21032
rect 12268 21004 12296 21032
rect 14366 21020 14372 21072
rect 14424 21060 14430 21072
rect 14424 21032 14504 21060
rect 14424 21020 14430 21032
rect 5905 20995 5963 21001
rect 5905 20992 5917 20995
rect 5868 20964 5917 20992
rect 5868 20952 5874 20964
rect 5905 20961 5917 20964
rect 5951 20961 5963 20995
rect 5905 20955 5963 20961
rect 6089 20995 6147 21001
rect 6089 20961 6101 20995
rect 6135 20961 6147 20995
rect 8941 20995 8999 21001
rect 7498 20964 8340 20992
rect 6089 20955 6147 20961
rect 5261 20927 5319 20933
rect 5261 20893 5273 20927
rect 5307 20924 5319 20927
rect 5307 20896 5396 20924
rect 5307 20893 5319 20896
rect 5261 20887 5319 20893
rect 5368 20865 5396 20896
rect 5353 20859 5411 20865
rect 5353 20825 5365 20859
rect 5399 20825 5411 20859
rect 5353 20819 5411 20825
rect 5920 20788 5948 20955
rect 6365 20927 6423 20933
rect 6365 20893 6377 20927
rect 6411 20924 6423 20927
rect 7837 20927 7895 20933
rect 6411 20896 7788 20924
rect 6411 20893 6423 20896
rect 6365 20887 6423 20893
rect 7760 20856 7788 20896
rect 7837 20893 7849 20927
rect 7883 20924 7895 20927
rect 8205 20927 8263 20933
rect 8205 20924 8217 20927
rect 7883 20896 8217 20924
rect 7883 20893 7895 20896
rect 7837 20887 7895 20893
rect 8205 20893 8217 20896
rect 8251 20893 8263 20927
rect 8312 20924 8340 20964
rect 8941 20961 8953 20995
rect 8987 20961 8999 20995
rect 8941 20955 8999 20961
rect 9858 20952 9864 21004
rect 9916 20992 9922 21004
rect 10505 20995 10563 21001
rect 10505 20992 10517 20995
rect 9916 20964 10517 20992
rect 9916 20952 9922 20964
rect 10505 20961 10517 20964
rect 10551 20961 10563 20995
rect 10505 20955 10563 20961
rect 10873 20995 10931 21001
rect 10873 20961 10885 20995
rect 10919 20961 10931 20995
rect 10873 20955 10931 20961
rect 9033 20927 9091 20933
rect 9033 20924 9045 20927
rect 8312 20896 9045 20924
rect 8205 20887 8263 20893
rect 9033 20893 9045 20896
rect 9079 20893 9091 20927
rect 9033 20887 9091 20893
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20924 9367 20927
rect 9950 20924 9956 20936
rect 9355 20896 9956 20924
rect 9355 20893 9367 20896
rect 9309 20887 9367 20893
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10134 20884 10140 20936
rect 10192 20884 10198 20936
rect 10226 20884 10232 20936
rect 10284 20884 10290 20936
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 10414 20927 10472 20933
rect 10414 20893 10426 20927
rect 10460 20924 10472 20927
rect 10778 20924 10784 20936
rect 10460 20896 10784 20924
rect 10460 20893 10472 20896
rect 10414 20887 10472 20893
rect 10045 20859 10103 20865
rect 10045 20856 10057 20859
rect 7760 20828 10057 20856
rect 10045 20825 10057 20828
rect 10091 20825 10103 20859
rect 10152 20856 10180 20884
rect 10336 20856 10364 20887
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 10152 20828 10364 20856
rect 10888 20856 10916 20955
rect 10962 20952 10968 21004
rect 11020 20992 11026 21004
rect 11057 20995 11115 21001
rect 11057 20992 11069 20995
rect 11020 20964 11069 20992
rect 11020 20952 11026 20964
rect 11057 20961 11069 20964
rect 11103 20961 11115 20995
rect 11057 20955 11115 20961
rect 11330 20952 11336 21004
rect 11388 20992 11394 21004
rect 11425 20995 11483 21001
rect 11425 20992 11437 20995
rect 11388 20964 11437 20992
rect 11388 20952 11394 20964
rect 11425 20961 11437 20964
rect 11471 20992 11483 20995
rect 11974 20992 11980 21004
rect 11471 20964 11980 20992
rect 11471 20961 11483 20964
rect 11425 20955 11483 20961
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 12250 20952 12256 21004
rect 12308 20952 12314 21004
rect 12434 20952 12440 21004
rect 12492 20952 12498 21004
rect 14476 21001 14504 21032
rect 14642 21020 14648 21072
rect 14700 21060 14706 21072
rect 15013 21063 15071 21069
rect 15013 21060 15025 21063
rect 14700 21032 15025 21060
rect 14700 21020 14706 21032
rect 15013 21029 15025 21032
rect 15059 21029 15071 21063
rect 15013 21023 15071 21029
rect 14461 20995 14519 21001
rect 14461 20961 14473 20995
rect 14507 20961 14519 20995
rect 14461 20955 14519 20961
rect 16850 20952 16856 21004
rect 16908 20952 16914 21004
rect 11149 20927 11207 20933
rect 11149 20893 11161 20927
rect 11195 20893 11207 20927
rect 11149 20887 11207 20893
rect 10962 20856 10968 20868
rect 10888 20828 10968 20856
rect 10045 20819 10103 20825
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 6454 20788 6460 20800
rect 5920 20760 6460 20788
rect 6454 20748 6460 20760
rect 6512 20748 6518 20800
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 8849 20791 8907 20797
rect 8849 20788 8861 20791
rect 8536 20760 8861 20788
rect 8536 20748 8542 20760
rect 8849 20757 8861 20760
rect 8895 20757 8907 20791
rect 8849 20751 8907 20757
rect 9674 20748 9680 20800
rect 9732 20788 9738 20800
rect 11164 20788 11192 20887
rect 11514 20884 11520 20936
rect 11572 20924 11578 20936
rect 11793 20927 11851 20933
rect 11793 20924 11805 20927
rect 11572 20896 11805 20924
rect 11572 20884 11578 20896
rect 11793 20893 11805 20896
rect 11839 20924 11851 20927
rect 12452 20924 12480 20952
rect 11839 20896 12480 20924
rect 11839 20893 11851 20896
rect 11793 20887 11851 20893
rect 13630 20884 13636 20936
rect 13688 20884 13694 20936
rect 17972 20924 18000 21088
rect 18340 21001 18368 21100
rect 19610 21088 19616 21100
rect 19668 21088 19674 21140
rect 21266 21088 21272 21140
rect 21324 21128 21330 21140
rect 21361 21131 21419 21137
rect 21361 21128 21373 21131
rect 21324 21100 21373 21128
rect 21324 21088 21330 21100
rect 21361 21097 21373 21100
rect 21407 21097 21419 21131
rect 21361 21091 21419 21097
rect 23753 21131 23811 21137
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 26878 21128 26884 21140
rect 23799 21100 26884 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 20714 21060 20720 21072
rect 19826 21032 20720 21060
rect 20714 21020 20720 21032
rect 20772 21020 20778 21072
rect 20916 21032 21220 21060
rect 18325 20995 18383 21001
rect 18325 20961 18337 20995
rect 18371 20961 18383 20995
rect 18325 20955 18383 20961
rect 20622 20952 20628 21004
rect 20680 20992 20686 21004
rect 20916 20992 20944 21032
rect 21192 21001 21220 21032
rect 22370 21020 22376 21072
rect 22428 21060 22434 21072
rect 23860 21060 23888 21100
rect 26878 21088 26884 21100
rect 26936 21088 26942 21140
rect 27801 21131 27859 21137
rect 27801 21097 27813 21131
rect 27847 21128 27859 21131
rect 27982 21128 27988 21140
rect 27847 21100 27988 21128
rect 27847 21097 27859 21100
rect 27801 21091 27859 21097
rect 27982 21088 27988 21100
rect 28040 21128 28046 21140
rect 28040 21100 28396 21128
rect 28040 21088 28046 21100
rect 28368 21072 28396 21100
rect 28442 21088 28448 21140
rect 28500 21128 28506 21140
rect 29546 21128 29552 21140
rect 28500 21100 29552 21128
rect 28500 21088 28506 21100
rect 29546 21088 29552 21100
rect 29604 21128 29610 21140
rect 30301 21131 30359 21137
rect 30301 21128 30313 21131
rect 29604 21100 30313 21128
rect 29604 21088 29610 21100
rect 30301 21097 30313 21100
rect 30347 21097 30359 21131
rect 30301 21091 30359 21097
rect 30469 21131 30527 21137
rect 30469 21097 30481 21131
rect 30515 21128 30527 21131
rect 30853 21131 30911 21137
rect 30853 21128 30865 21131
rect 30515 21100 30865 21128
rect 30515 21097 30527 21100
rect 30469 21091 30527 21097
rect 30853 21097 30865 21100
rect 30899 21128 30911 21131
rect 31294 21128 31300 21140
rect 30899 21100 31300 21128
rect 30899 21097 30911 21100
rect 30853 21091 30911 21097
rect 31294 21088 31300 21100
rect 31352 21088 31358 21140
rect 32582 21128 32588 21140
rect 31726 21100 32588 21128
rect 22428 21032 23888 21060
rect 22428 21020 22434 21032
rect 20680 20964 20944 20992
rect 20993 20995 21051 21001
rect 20680 20952 20686 20964
rect 20993 20961 21005 20995
rect 21039 20992 21051 20995
rect 21177 20995 21235 21001
rect 21039 20964 21073 20992
rect 21039 20961 21051 20964
rect 20993 20955 21051 20961
rect 21177 20961 21189 20995
rect 21223 20992 21235 20995
rect 21266 20992 21272 21004
rect 21223 20964 21272 20992
rect 21223 20961 21235 20964
rect 21177 20955 21235 20961
rect 17972 20896 18368 20924
rect 18340 20868 18368 20896
rect 18598 20884 18604 20936
rect 18656 20884 18662 20936
rect 20073 20927 20131 20933
rect 20073 20893 20085 20927
rect 20119 20924 20131 20927
rect 20809 20927 20867 20933
rect 20809 20924 20821 20927
rect 20119 20896 20821 20924
rect 20119 20893 20131 20896
rect 20073 20887 20131 20893
rect 20809 20893 20821 20896
rect 20855 20893 20867 20927
rect 20809 20887 20867 20893
rect 12894 20816 12900 20868
rect 12952 20856 12958 20868
rect 16666 20856 16672 20868
rect 12952 20828 16672 20856
rect 12952 20816 12958 20828
rect 16666 20816 16672 20828
rect 16724 20816 16730 20868
rect 16758 20816 16764 20868
rect 16816 20856 16822 20868
rect 17954 20856 17960 20868
rect 16816 20828 17960 20856
rect 16816 20816 16822 20828
rect 17954 20816 17960 20828
rect 18012 20816 18018 20868
rect 18322 20816 18328 20868
rect 18380 20816 18386 20868
rect 20824 20856 20852 20887
rect 20898 20884 20904 20936
rect 20956 20924 20962 20936
rect 21008 20924 21036 20955
rect 21266 20952 21272 20964
rect 21324 20952 21330 21004
rect 21358 20952 21364 21004
rect 21416 20992 21422 21004
rect 21637 20995 21695 21001
rect 21637 20992 21649 20995
rect 21416 20964 21649 20992
rect 21416 20952 21422 20964
rect 21637 20961 21649 20964
rect 21683 20992 21695 20995
rect 22646 20992 22652 21004
rect 21683 20964 22652 20992
rect 21683 20961 21695 20964
rect 21637 20955 21695 20961
rect 22646 20952 22652 20964
rect 22704 20952 22710 21004
rect 23860 21001 23888 21032
rect 23937 21063 23995 21069
rect 23937 21029 23949 21063
rect 23983 21060 23995 21063
rect 24486 21060 24492 21072
rect 23983 21032 24492 21060
rect 23983 21029 23995 21032
rect 23937 21023 23995 21029
rect 24486 21020 24492 21032
rect 24544 21060 24550 21072
rect 24762 21060 24768 21072
rect 24544 21032 24768 21060
rect 24544 21020 24550 21032
rect 24762 21020 24768 21032
rect 24820 21020 24826 21072
rect 26050 21060 26056 21072
rect 25792 21032 26056 21060
rect 23845 20995 23903 21001
rect 23845 20961 23857 20995
rect 23891 20961 23903 20995
rect 23845 20955 23903 20961
rect 24026 20952 24032 21004
rect 24084 20952 24090 21004
rect 25590 20952 25596 21004
rect 25648 20952 25654 21004
rect 25792 21001 25820 21032
rect 26050 21020 26056 21032
rect 26108 21020 26114 21072
rect 26160 21032 28120 21060
rect 25777 20995 25835 21001
rect 25777 20961 25789 20995
rect 25823 20961 25835 20995
rect 25777 20955 25835 20961
rect 21545 20927 21603 20933
rect 21545 20924 21557 20927
rect 20956 20896 21557 20924
rect 20956 20884 20962 20896
rect 21545 20893 21557 20896
rect 21591 20893 21603 20927
rect 21545 20887 21603 20893
rect 21910 20884 21916 20936
rect 21968 20884 21974 20936
rect 22005 20927 22063 20933
rect 22005 20893 22017 20927
rect 22051 20924 22063 20927
rect 23658 20924 23664 20936
rect 22051 20896 23664 20924
rect 22051 20893 22063 20896
rect 22005 20887 22063 20893
rect 23658 20884 23664 20896
rect 23716 20884 23722 20936
rect 25317 20927 25375 20933
rect 23768 20896 24072 20924
rect 23768 20856 23796 20896
rect 20824 20828 23796 20856
rect 24044 20856 24072 20896
rect 25317 20893 25329 20927
rect 25363 20924 25375 20927
rect 25409 20927 25467 20933
rect 25409 20924 25421 20927
rect 25363 20896 25421 20924
rect 25363 20893 25375 20896
rect 25317 20887 25375 20893
rect 25409 20893 25421 20896
rect 25455 20893 25467 20927
rect 25409 20887 25467 20893
rect 26160 20856 26188 21032
rect 26970 20952 26976 21004
rect 27028 20952 27034 21004
rect 27062 20952 27068 21004
rect 27120 20952 27126 21004
rect 27338 20952 27344 21004
rect 27396 20992 27402 21004
rect 27433 20995 27491 21001
rect 27433 20992 27445 20995
rect 27396 20964 27445 20992
rect 27396 20952 27402 20964
rect 27433 20961 27445 20964
rect 27479 20961 27491 20995
rect 27433 20955 27491 20961
rect 27706 20952 27712 21004
rect 27764 20952 27770 21004
rect 27798 20952 27804 21004
rect 27856 20992 27862 21004
rect 27985 20995 28043 21001
rect 27985 20992 27997 20995
rect 27856 20964 27997 20992
rect 27856 20952 27862 20964
rect 27985 20961 27997 20964
rect 28031 20961 28043 20995
rect 28092 20992 28120 21032
rect 28166 21020 28172 21072
rect 28224 21020 28230 21072
rect 28350 21020 28356 21072
rect 28408 21020 28414 21072
rect 29362 21020 29368 21072
rect 29420 21060 29426 21072
rect 29914 21060 29920 21072
rect 29420 21032 29920 21060
rect 29420 21020 29426 21032
rect 29914 21020 29920 21032
rect 29972 21060 29978 21072
rect 30101 21063 30159 21069
rect 30101 21060 30113 21063
rect 29972 21032 30113 21060
rect 29972 21020 29978 21032
rect 30101 21029 30113 21032
rect 30147 21029 30159 21063
rect 30101 21023 30159 21029
rect 30650 21020 30656 21072
rect 30708 21020 30714 21072
rect 31726 20992 31754 21100
rect 32582 21088 32588 21100
rect 32640 21088 32646 21140
rect 33410 20992 33416 21004
rect 28092 20964 31754 20992
rect 33152 20964 33416 20992
rect 27985 20955 28043 20961
rect 26513 20927 26571 20933
rect 26513 20893 26525 20927
rect 26559 20924 26571 20927
rect 26694 20924 26700 20936
rect 26559 20896 26700 20924
rect 26559 20893 26571 20896
rect 26513 20887 26571 20893
rect 26694 20884 26700 20896
rect 26752 20884 26758 20936
rect 27246 20884 27252 20936
rect 27304 20924 27310 20936
rect 27816 20924 27844 20952
rect 33152 20936 33180 20964
rect 33410 20952 33416 20964
rect 33468 20992 33474 21004
rect 33781 20995 33839 21001
rect 33781 20992 33793 20995
rect 33468 20964 33793 20992
rect 33468 20952 33474 20964
rect 33781 20961 33793 20964
rect 33827 20961 33839 20995
rect 33781 20955 33839 20961
rect 27304 20896 27844 20924
rect 27304 20884 27310 20896
rect 30466 20884 30472 20936
rect 30524 20924 30530 20936
rect 30650 20924 30656 20936
rect 30524 20896 30656 20924
rect 30524 20884 30530 20896
rect 30650 20884 30656 20896
rect 30708 20884 30714 20936
rect 31018 20884 31024 20936
rect 31076 20924 31082 20936
rect 31113 20927 31171 20933
rect 31113 20924 31125 20927
rect 31076 20896 31125 20924
rect 31076 20884 31082 20896
rect 31113 20893 31125 20896
rect 31159 20893 31171 20927
rect 31113 20887 31171 20893
rect 31754 20884 31760 20936
rect 31812 20884 31818 20936
rect 32306 20884 32312 20936
rect 32364 20924 32370 20936
rect 32585 20927 32643 20933
rect 32585 20924 32597 20927
rect 32364 20896 32597 20924
rect 32364 20884 32370 20896
rect 32585 20893 32597 20896
rect 32631 20893 32643 20927
rect 32585 20887 32643 20893
rect 33134 20884 33140 20936
rect 33192 20884 33198 20936
rect 33318 20884 33324 20936
rect 33376 20884 33382 20936
rect 24044 20828 26188 20856
rect 9732 20760 11192 20788
rect 11241 20791 11299 20797
rect 9732 20748 9738 20760
rect 11241 20757 11253 20791
rect 11287 20788 11299 20791
rect 11514 20788 11520 20800
rect 11287 20760 11520 20788
rect 11287 20757 11299 20760
rect 11241 20751 11299 20757
rect 11514 20748 11520 20760
rect 11572 20748 11578 20800
rect 12345 20791 12403 20797
rect 12345 20757 12357 20791
rect 12391 20788 12403 20791
rect 13078 20788 13084 20800
rect 12391 20760 13084 20788
rect 12391 20757 12403 20760
rect 12345 20751 12403 20757
rect 13078 20748 13084 20760
rect 13136 20788 13142 20800
rect 13354 20788 13360 20800
rect 13136 20760 13360 20788
rect 13136 20748 13142 20760
rect 13354 20748 13360 20760
rect 13412 20748 13418 20800
rect 14274 20748 14280 20800
rect 14332 20748 14338 20800
rect 15930 20748 15936 20800
rect 15988 20788 15994 20800
rect 16301 20791 16359 20797
rect 16301 20788 16313 20791
rect 15988 20760 16313 20788
rect 15988 20748 15994 20760
rect 16301 20757 16313 20760
rect 16347 20757 16359 20791
rect 16301 20751 16359 20757
rect 18138 20748 18144 20800
rect 18196 20788 18202 20800
rect 18690 20788 18696 20800
rect 18196 20760 18696 20788
rect 18196 20748 18202 20760
rect 18690 20748 18696 20760
rect 18748 20748 18754 20800
rect 20254 20748 20260 20800
rect 20312 20748 20318 20800
rect 21174 20748 21180 20800
rect 21232 20748 21238 20800
rect 21266 20748 21272 20800
rect 21324 20788 21330 20800
rect 22370 20788 22376 20800
rect 21324 20760 22376 20788
rect 21324 20748 21330 20760
rect 22370 20748 22376 20760
rect 22428 20748 22434 20800
rect 22646 20748 22652 20800
rect 22704 20788 22710 20800
rect 24026 20788 24032 20800
rect 22704 20760 24032 20788
rect 22704 20748 22710 20760
rect 24026 20748 24032 20760
rect 24084 20788 24090 20800
rect 24305 20791 24363 20797
rect 24305 20788 24317 20791
rect 24084 20760 24317 20788
rect 24084 20748 24090 20760
rect 24305 20757 24317 20760
rect 24351 20757 24363 20791
rect 24305 20751 24363 20757
rect 24486 20748 24492 20800
rect 24544 20788 24550 20800
rect 24673 20791 24731 20797
rect 24673 20788 24685 20791
rect 24544 20760 24685 20788
rect 24544 20748 24550 20760
rect 24673 20757 24685 20760
rect 24719 20757 24731 20791
rect 24673 20751 24731 20757
rect 25774 20748 25780 20800
rect 25832 20788 25838 20800
rect 25869 20791 25927 20797
rect 25869 20788 25881 20791
rect 25832 20760 25881 20788
rect 25832 20748 25838 20760
rect 25869 20757 25881 20760
rect 25915 20788 25927 20791
rect 26326 20788 26332 20800
rect 25915 20760 26332 20788
rect 25915 20757 25927 20760
rect 25869 20751 25927 20757
rect 26326 20748 26332 20760
rect 26384 20748 26390 20800
rect 26712 20788 26740 20884
rect 30852 20828 31248 20856
rect 27341 20791 27399 20797
rect 27341 20788 27353 20791
rect 26712 20760 27353 20788
rect 27341 20757 27353 20760
rect 27387 20757 27399 20791
rect 27341 20751 27399 20757
rect 27617 20791 27675 20797
rect 27617 20757 27629 20791
rect 27663 20788 27675 20791
rect 27982 20788 27988 20800
rect 27663 20760 27988 20788
rect 27663 20757 27675 20760
rect 27617 20751 27675 20757
rect 27982 20748 27988 20760
rect 28040 20748 28046 20800
rect 28350 20748 28356 20800
rect 28408 20788 28414 20800
rect 30852 20797 30880 20828
rect 31220 20800 31248 20828
rect 30285 20791 30343 20797
rect 30285 20788 30297 20791
rect 28408 20760 30297 20788
rect 28408 20748 28414 20760
rect 30285 20757 30297 20760
rect 30331 20757 30343 20791
rect 30285 20751 30343 20757
rect 30837 20791 30895 20797
rect 30837 20757 30849 20791
rect 30883 20757 30895 20791
rect 30837 20751 30895 20757
rect 30926 20748 30932 20800
rect 30984 20788 30990 20800
rect 31021 20791 31079 20797
rect 31021 20788 31033 20791
rect 30984 20760 31033 20788
rect 30984 20748 30990 20760
rect 31021 20757 31033 20760
rect 31067 20757 31079 20791
rect 31021 20751 31079 20757
rect 31202 20748 31208 20800
rect 31260 20748 31266 20800
rect 32030 20748 32036 20800
rect 32088 20748 32094 20800
rect 32582 20748 32588 20800
rect 32640 20788 32646 20800
rect 32769 20791 32827 20797
rect 32769 20788 32781 20791
rect 32640 20760 32781 20788
rect 32640 20748 32646 20760
rect 32769 20757 32781 20760
rect 32815 20757 32827 20791
rect 32769 20751 32827 20757
rect 33870 20748 33876 20800
rect 33928 20748 33934 20800
rect 2760 20698 34316 20720
rect 2760 20646 6550 20698
rect 6602 20646 6614 20698
rect 6666 20646 6678 20698
rect 6730 20646 6742 20698
rect 6794 20646 6806 20698
rect 6858 20646 14439 20698
rect 14491 20646 14503 20698
rect 14555 20646 14567 20698
rect 14619 20646 14631 20698
rect 14683 20646 14695 20698
rect 14747 20646 22328 20698
rect 22380 20646 22392 20698
rect 22444 20646 22456 20698
rect 22508 20646 22520 20698
rect 22572 20646 22584 20698
rect 22636 20646 30217 20698
rect 30269 20646 30281 20698
rect 30333 20646 30345 20698
rect 30397 20646 30409 20698
rect 30461 20646 30473 20698
rect 30525 20646 34316 20698
rect 2760 20624 34316 20646
rect 5166 20544 5172 20596
rect 5224 20544 5230 20596
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 9033 20587 9091 20593
rect 9033 20584 9045 20587
rect 6880 20556 9045 20584
rect 6880 20544 6886 20556
rect 9033 20553 9045 20556
rect 9079 20553 9091 20587
rect 9033 20547 9091 20553
rect 9858 20544 9864 20596
rect 9916 20544 9922 20596
rect 9953 20587 10011 20593
rect 9953 20553 9965 20587
rect 9999 20584 10011 20587
rect 10226 20584 10232 20596
rect 9999 20556 10232 20584
rect 9999 20553 10011 20556
rect 9953 20547 10011 20553
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 10778 20544 10784 20596
rect 10836 20584 10842 20596
rect 11330 20584 11336 20596
rect 10836 20556 11336 20584
rect 10836 20544 10842 20556
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20448 3663 20451
rect 4246 20448 4252 20460
rect 3651 20420 4252 20448
rect 3651 20417 3663 20420
rect 3605 20411 3663 20417
rect 4246 20408 4252 20420
rect 4304 20408 4310 20460
rect 4338 20408 4344 20460
rect 4396 20448 4402 20460
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 4396 20420 4537 20448
rect 4396 20408 4402 20420
rect 4525 20417 4537 20420
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 5184 20380 5212 20544
rect 9490 20476 9496 20528
rect 9548 20476 9554 20528
rect 9585 20519 9643 20525
rect 9585 20485 9597 20519
rect 9631 20516 9643 20519
rect 9674 20516 9680 20528
rect 9631 20488 9680 20516
rect 9631 20485 9643 20488
rect 9585 20479 9643 20485
rect 9674 20476 9680 20488
rect 9732 20476 9738 20528
rect 10137 20519 10195 20525
rect 10137 20485 10149 20519
rect 10183 20516 10195 20519
rect 10962 20516 10968 20528
rect 10183 20488 10968 20516
rect 10183 20485 10195 20488
rect 10137 20479 10195 20485
rect 10962 20476 10968 20488
rect 11020 20476 11026 20528
rect 5626 20408 5632 20460
rect 5684 20448 5690 20460
rect 5902 20448 5908 20460
rect 5684 20420 5908 20448
rect 5684 20408 5690 20420
rect 5902 20408 5908 20420
rect 5960 20408 5966 20460
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7469 20451 7527 20457
rect 7469 20448 7481 20451
rect 7156 20420 7481 20448
rect 7156 20408 7162 20420
rect 7469 20417 7481 20420
rect 7515 20448 7527 20451
rect 8018 20448 8024 20460
rect 7515 20420 8024 20448
rect 7515 20417 7527 20420
rect 7469 20411 7527 20417
rect 8018 20408 8024 20420
rect 8076 20408 8082 20460
rect 8478 20408 8484 20460
rect 8536 20408 8542 20460
rect 8665 20451 8723 20457
rect 8665 20417 8677 20451
rect 8711 20448 8723 20451
rect 8846 20448 8852 20460
rect 8711 20420 8852 20448
rect 8711 20417 8723 20420
rect 8665 20411 8723 20417
rect 8846 20408 8852 20420
rect 8904 20448 8910 20460
rect 10042 20448 10048 20460
rect 8904 20420 10048 20448
rect 8904 20408 8910 20420
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 10413 20451 10471 20457
rect 10413 20417 10425 20451
rect 10459 20448 10471 20451
rect 10686 20448 10692 20460
rect 10459 20420 10692 20448
rect 10459 20417 10471 20420
rect 10413 20411 10471 20417
rect 10686 20408 10692 20420
rect 10744 20408 10750 20460
rect 10870 20408 10876 20460
rect 10928 20408 10934 20460
rect 11072 20457 11100 20556
rect 11330 20544 11336 20556
rect 11388 20544 11394 20596
rect 13814 20544 13820 20596
rect 13872 20544 13878 20596
rect 18598 20544 18604 20596
rect 18656 20544 18662 20596
rect 19058 20544 19064 20596
rect 19116 20584 19122 20596
rect 19886 20584 19892 20596
rect 19116 20556 19892 20584
rect 19116 20544 19122 20556
rect 19886 20544 19892 20556
rect 19944 20544 19950 20596
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 20993 20587 21051 20593
rect 20993 20584 21005 20587
rect 20772 20556 21005 20584
rect 20772 20544 20778 20556
rect 20993 20553 21005 20556
rect 21039 20553 21051 20587
rect 20993 20547 21051 20553
rect 21361 20587 21419 20593
rect 21361 20553 21373 20587
rect 21407 20584 21419 20587
rect 21542 20584 21548 20596
rect 21407 20556 21548 20584
rect 21407 20553 21419 20556
rect 21361 20547 21419 20553
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 22373 20587 22431 20593
rect 22373 20584 22385 20587
rect 21876 20556 22385 20584
rect 21876 20544 21882 20556
rect 22373 20553 22385 20556
rect 22419 20584 22431 20587
rect 23566 20584 23572 20596
rect 22419 20556 23572 20584
rect 22419 20553 22431 20556
rect 22373 20547 22431 20553
rect 23566 20544 23572 20556
rect 23624 20544 23630 20596
rect 24228 20556 25452 20584
rect 19613 20519 19671 20525
rect 11348 20488 11836 20516
rect 11348 20457 11376 20488
rect 11057 20451 11115 20457
rect 11057 20417 11069 20451
rect 11103 20417 11115 20451
rect 11057 20411 11115 20417
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20417 11391 20451
rect 11333 20411 11391 20417
rect 11698 20408 11704 20460
rect 11756 20408 11762 20460
rect 11808 20448 11836 20488
rect 19613 20485 19625 20519
rect 19659 20516 19671 20519
rect 24228 20516 24256 20556
rect 19659 20488 24256 20516
rect 19659 20485 19671 20488
rect 19613 20479 19671 20485
rect 12342 20448 12348 20460
rect 11808 20420 12348 20448
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 14826 20408 14832 20460
rect 14884 20448 14890 20460
rect 15562 20448 15568 20460
rect 14884 20420 15568 20448
rect 14884 20408 14890 20420
rect 15562 20408 15568 20420
rect 15620 20448 15626 20460
rect 15749 20451 15807 20457
rect 15749 20448 15761 20451
rect 15620 20420 15761 20448
rect 15620 20408 15626 20420
rect 15749 20417 15761 20420
rect 15795 20417 15807 20451
rect 15749 20411 15807 20417
rect 17497 20451 17555 20457
rect 17497 20417 17509 20451
rect 17543 20448 17555 20451
rect 17589 20451 17647 20457
rect 17589 20448 17601 20451
rect 17543 20420 17601 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 17589 20417 17601 20420
rect 17635 20417 17647 20451
rect 17589 20411 17647 20417
rect 18046 20408 18052 20460
rect 18104 20448 18110 20460
rect 19150 20448 19156 20460
rect 18104 20420 19156 20448
rect 18104 20408 18110 20420
rect 19150 20408 19156 20420
rect 19208 20408 19214 20460
rect 20254 20448 20260 20460
rect 19352 20420 20260 20448
rect 4111 20352 5212 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 7834 20340 7840 20392
rect 7892 20380 7898 20392
rect 8110 20380 8116 20392
rect 7892 20352 8116 20380
rect 7892 20340 7898 20352
rect 8110 20340 8116 20352
rect 8168 20340 8174 20392
rect 8496 20380 8524 20408
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 8496 20352 9413 20380
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9677 20383 9735 20389
rect 9677 20349 9689 20383
rect 9723 20380 9735 20383
rect 9950 20380 9956 20392
rect 9723 20352 9956 20380
rect 9723 20349 9735 20352
rect 9677 20343 9735 20349
rect 9950 20340 9956 20352
rect 10008 20340 10014 20392
rect 7193 20315 7251 20321
rect 6762 20284 7052 20312
rect 7024 20256 7052 20284
rect 7193 20281 7205 20315
rect 7239 20312 7251 20315
rect 7650 20312 7656 20324
rect 7239 20284 7656 20312
rect 7239 20281 7251 20284
rect 7193 20275 7251 20281
rect 7650 20272 7656 20284
rect 7708 20272 7714 20324
rect 7926 20272 7932 20324
rect 7984 20312 7990 20324
rect 8389 20315 8447 20321
rect 8389 20312 8401 20315
rect 7984 20284 8401 20312
rect 7984 20272 7990 20284
rect 8389 20281 8401 20284
rect 8435 20281 8447 20315
rect 8389 20275 8447 20281
rect 10042 20272 10048 20324
rect 10100 20312 10106 20324
rect 10410 20312 10416 20324
rect 10100 20284 10416 20312
rect 10100 20272 10106 20284
rect 10410 20272 10416 20284
rect 10468 20272 10474 20324
rect 10704 20312 10732 20408
rect 10888 20380 10916 20408
rect 10965 20383 11023 20389
rect 10965 20380 10977 20383
rect 10888 20352 10977 20380
rect 10965 20349 10977 20352
rect 11011 20349 11023 20383
rect 10965 20343 11023 20349
rect 11422 20340 11428 20392
rect 11480 20340 11486 20392
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18012 20352 18521 20380
rect 18012 20340 18018 20352
rect 18509 20349 18521 20352
rect 18555 20380 18567 20383
rect 18874 20380 18880 20392
rect 18555 20352 18880 20380
rect 18555 20349 18567 20352
rect 18509 20343 18567 20349
rect 18874 20340 18880 20352
rect 18932 20340 18938 20392
rect 19061 20383 19119 20389
rect 19061 20349 19073 20383
rect 19107 20380 19119 20383
rect 19352 20380 19380 20420
rect 20254 20408 20260 20420
rect 20312 20408 20318 20460
rect 21450 20408 21456 20460
rect 21508 20448 21514 20460
rect 21508 20420 22094 20448
rect 21508 20408 21514 20420
rect 19107 20352 19380 20380
rect 19107 20349 19119 20352
rect 19061 20343 19119 20349
rect 19426 20340 19432 20392
rect 19484 20340 19490 20392
rect 19702 20340 19708 20392
rect 19760 20380 19766 20392
rect 20165 20383 20223 20389
rect 20165 20380 20177 20383
rect 19760 20352 20177 20380
rect 19760 20340 19766 20352
rect 20165 20349 20177 20352
rect 20211 20349 20223 20383
rect 20165 20343 20223 20349
rect 21082 20340 21088 20392
rect 21140 20340 21146 20392
rect 21266 20340 21272 20392
rect 21324 20380 21330 20392
rect 21545 20383 21603 20389
rect 21545 20380 21557 20383
rect 21324 20352 21557 20380
rect 21324 20340 21330 20352
rect 21545 20349 21557 20352
rect 21591 20349 21603 20383
rect 21545 20343 21603 20349
rect 21637 20383 21695 20389
rect 21637 20349 21649 20383
rect 21683 20380 21695 20383
rect 21818 20380 21824 20392
rect 21683 20352 21824 20380
rect 21683 20349 21695 20352
rect 21637 20343 21695 20349
rect 11609 20315 11667 20321
rect 10704 20284 11560 20312
rect 3694 20204 3700 20256
rect 3752 20204 3758 20256
rect 4157 20247 4215 20253
rect 4157 20213 4169 20247
rect 4203 20244 4215 20247
rect 5350 20244 5356 20256
rect 4203 20216 5356 20244
rect 4203 20213 4215 20216
rect 4157 20207 4215 20213
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 5718 20204 5724 20256
rect 5776 20204 5782 20256
rect 6362 20204 6368 20256
rect 6420 20244 6426 20256
rect 6822 20244 6828 20256
rect 6420 20216 6828 20244
rect 6420 20204 6426 20216
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7006 20204 7012 20256
rect 7064 20204 7070 20256
rect 8018 20204 8024 20256
rect 8076 20204 8082 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 10594 20244 10600 20256
rect 9456 20216 10600 20244
rect 9456 20204 9462 20216
rect 10594 20204 10600 20216
rect 10652 20204 10658 20256
rect 10870 20204 10876 20256
rect 10928 20244 10934 20256
rect 11149 20247 11207 20253
rect 11149 20244 11161 20247
rect 10928 20216 11161 20244
rect 10928 20204 10934 20216
rect 11149 20213 11161 20216
rect 11195 20213 11207 20247
rect 11532 20244 11560 20284
rect 11609 20281 11621 20315
rect 11655 20312 11667 20315
rect 11977 20315 12035 20321
rect 11977 20312 11989 20315
rect 11655 20284 11989 20312
rect 11655 20281 11667 20284
rect 11609 20275 11667 20281
rect 11977 20281 11989 20284
rect 12023 20281 12035 20315
rect 11977 20275 12035 20281
rect 12986 20272 12992 20324
rect 13044 20272 13050 20324
rect 15194 20312 15200 20324
rect 14858 20284 15200 20312
rect 15194 20272 15200 20284
rect 15252 20272 15258 20324
rect 15289 20315 15347 20321
rect 15289 20281 15301 20315
rect 15335 20281 15347 20315
rect 15289 20275 15347 20281
rect 12066 20244 12072 20256
rect 11532 20216 12072 20244
rect 11149 20207 11207 20213
rect 12066 20204 12072 20216
rect 12124 20204 12130 20256
rect 13446 20204 13452 20256
rect 13504 20204 13510 20256
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 15304 20244 15332 20275
rect 16022 20272 16028 20324
rect 16080 20272 16086 20324
rect 18417 20315 18475 20321
rect 18417 20312 18429 20315
rect 17250 20284 18429 20312
rect 18417 20281 18429 20284
rect 18463 20281 18475 20315
rect 18417 20275 18475 20281
rect 19978 20272 19984 20324
rect 20036 20312 20042 20324
rect 20441 20315 20499 20321
rect 20441 20312 20453 20315
rect 20036 20284 20453 20312
rect 20036 20272 20042 20284
rect 20441 20281 20453 20284
rect 20487 20281 20499 20315
rect 20441 20275 20499 20281
rect 14332 20216 15332 20244
rect 14332 20204 14338 20216
rect 16758 20204 16764 20256
rect 16816 20244 16822 20256
rect 17862 20244 17868 20256
rect 16816 20216 17868 20244
rect 16816 20204 16822 20216
rect 17862 20204 17868 20216
rect 17920 20244 17926 20256
rect 18233 20247 18291 20253
rect 18233 20244 18245 20247
rect 17920 20216 18245 20244
rect 17920 20204 17926 20216
rect 18233 20213 18245 20216
rect 18279 20213 18291 20247
rect 18233 20207 18291 20213
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 18969 20247 19027 20253
rect 18969 20244 18981 20247
rect 18932 20216 18981 20244
rect 18932 20204 18938 20216
rect 18969 20213 18981 20216
rect 19015 20213 19027 20247
rect 18969 20207 19027 20213
rect 19886 20204 19892 20256
rect 19944 20244 19950 20256
rect 20073 20247 20131 20253
rect 20073 20244 20085 20247
rect 19944 20216 20085 20244
rect 19944 20204 19950 20216
rect 20073 20213 20085 20216
rect 20119 20244 20131 20247
rect 21744 20244 21772 20352
rect 21818 20340 21824 20352
rect 21876 20340 21882 20392
rect 21910 20340 21916 20392
rect 21968 20340 21974 20392
rect 22066 20380 22094 20420
rect 22554 20408 22560 20460
rect 22612 20448 22618 20460
rect 23934 20448 23940 20460
rect 22612 20420 23940 20448
rect 22612 20408 22618 20420
rect 23934 20408 23940 20420
rect 23992 20448 23998 20460
rect 24118 20448 24124 20460
rect 23992 20420 24124 20448
rect 23992 20408 23998 20420
rect 24118 20408 24124 20420
rect 24176 20408 24182 20460
rect 24397 20451 24455 20457
rect 24397 20417 24409 20451
rect 24443 20448 24455 20451
rect 24486 20448 24492 20460
rect 24443 20420 24492 20448
rect 24443 20417 24455 20420
rect 24397 20411 24455 20417
rect 24486 20408 24492 20420
rect 24544 20408 24550 20460
rect 25424 20448 25452 20556
rect 25590 20544 25596 20596
rect 25648 20584 25654 20596
rect 26053 20587 26111 20593
rect 26053 20584 26065 20587
rect 25648 20556 26065 20584
rect 25648 20544 25654 20556
rect 26053 20553 26065 20556
rect 26099 20553 26111 20587
rect 26053 20547 26111 20553
rect 26234 20544 26240 20596
rect 26292 20584 26298 20596
rect 26418 20584 26424 20596
rect 26292 20556 26424 20584
rect 26292 20544 26298 20556
rect 26418 20544 26424 20556
rect 26476 20544 26482 20596
rect 26694 20544 26700 20596
rect 26752 20544 26758 20596
rect 26973 20587 27031 20593
rect 26973 20553 26985 20587
rect 27019 20584 27031 20587
rect 27154 20584 27160 20596
rect 27019 20556 27160 20584
rect 27019 20553 27031 20556
rect 26973 20547 27031 20553
rect 27154 20544 27160 20556
rect 27212 20544 27218 20596
rect 27614 20544 27620 20596
rect 27672 20544 27678 20596
rect 27706 20544 27712 20596
rect 27764 20584 27770 20596
rect 27893 20587 27951 20593
rect 27893 20584 27905 20587
rect 27764 20556 27905 20584
rect 27764 20544 27770 20556
rect 27893 20553 27905 20556
rect 27939 20553 27951 20587
rect 27893 20547 27951 20553
rect 29454 20544 29460 20596
rect 29512 20544 29518 20596
rect 29822 20544 29828 20596
rect 29880 20584 29886 20596
rect 29917 20587 29975 20593
rect 29917 20584 29929 20587
rect 29880 20556 29929 20584
rect 29880 20544 29886 20556
rect 29917 20553 29929 20556
rect 29963 20553 29975 20587
rect 29917 20547 29975 20553
rect 31754 20544 31760 20596
rect 31812 20584 31818 20596
rect 31941 20587 31999 20593
rect 31941 20584 31953 20587
rect 31812 20556 31953 20584
rect 31812 20544 31818 20556
rect 31941 20553 31953 20556
rect 31987 20553 31999 20587
rect 31941 20547 31999 20553
rect 25869 20519 25927 20525
rect 25869 20485 25881 20519
rect 25915 20516 25927 20519
rect 26712 20516 26740 20544
rect 27724 20516 27752 20544
rect 25915 20488 26740 20516
rect 27172 20488 27752 20516
rect 28997 20519 29055 20525
rect 25915 20485 25927 20488
rect 25869 20479 25927 20485
rect 25424 20420 25912 20448
rect 23661 20383 23719 20389
rect 23661 20380 23673 20383
rect 22066 20352 23673 20380
rect 23661 20349 23673 20352
rect 23707 20349 23719 20383
rect 23661 20343 23719 20349
rect 22005 20315 22063 20321
rect 22005 20281 22017 20315
rect 22051 20312 22063 20315
rect 25774 20312 25780 20324
rect 22051 20284 24808 20312
rect 25622 20284 25780 20312
rect 22051 20281 22063 20284
rect 22005 20275 22063 20281
rect 20119 20216 21772 20244
rect 23753 20247 23811 20253
rect 20119 20213 20131 20216
rect 20073 20207 20131 20213
rect 23753 20213 23765 20247
rect 23799 20244 23811 20247
rect 23842 20244 23848 20256
rect 23799 20216 23848 20244
rect 23799 20213 23811 20216
rect 23753 20207 23811 20213
rect 23842 20204 23848 20216
rect 23900 20204 23906 20256
rect 24118 20204 24124 20256
rect 24176 20244 24182 20256
rect 24670 20244 24676 20256
rect 24176 20216 24676 20244
rect 24176 20204 24182 20216
rect 24670 20204 24676 20216
rect 24728 20204 24734 20256
rect 24780 20244 24808 20284
rect 25774 20272 25780 20284
rect 25832 20272 25838 20324
rect 25884 20312 25912 20420
rect 26326 20408 26332 20460
rect 26384 20408 26390 20460
rect 26050 20340 26056 20392
rect 26108 20380 26114 20392
rect 26237 20383 26295 20389
rect 26237 20380 26249 20383
rect 26108 20352 26249 20380
rect 26108 20340 26114 20352
rect 26237 20349 26249 20352
rect 26283 20349 26295 20383
rect 26344 20380 26372 20408
rect 26513 20383 26571 20389
rect 26513 20380 26525 20383
rect 26344 20352 26525 20380
rect 26237 20343 26295 20349
rect 26513 20349 26525 20352
rect 26559 20380 26571 20383
rect 26602 20380 26608 20392
rect 26559 20352 26608 20380
rect 26559 20349 26571 20352
rect 26513 20343 26571 20349
rect 26602 20340 26608 20352
rect 26660 20340 26666 20392
rect 27172 20389 27200 20488
rect 28997 20485 29009 20519
rect 29043 20485 29055 20519
rect 28997 20479 29055 20485
rect 30653 20519 30711 20525
rect 30653 20485 30665 20519
rect 30699 20516 30711 20519
rect 31478 20516 31484 20528
rect 30699 20488 31484 20516
rect 30699 20485 30711 20488
rect 30653 20479 30711 20485
rect 27985 20451 28043 20457
rect 27985 20448 27997 20451
rect 27264 20420 27997 20448
rect 27157 20383 27215 20389
rect 27157 20349 27169 20383
rect 27203 20349 27215 20383
rect 27157 20343 27215 20349
rect 26142 20312 26148 20324
rect 25884 20284 26148 20312
rect 26142 20272 26148 20284
rect 26200 20272 26206 20324
rect 26326 20272 26332 20324
rect 26384 20312 26390 20324
rect 27264 20312 27292 20420
rect 27985 20417 27997 20420
rect 28031 20417 28043 20451
rect 27985 20411 28043 20417
rect 27341 20383 27399 20389
rect 27341 20349 27353 20383
rect 27387 20380 27399 20383
rect 27522 20380 27528 20392
rect 27387 20352 27528 20380
rect 27387 20349 27399 20352
rect 27341 20343 27399 20349
rect 27522 20340 27528 20352
rect 27580 20340 27586 20392
rect 27614 20340 27620 20392
rect 27672 20340 27678 20392
rect 27709 20383 27767 20389
rect 27709 20349 27721 20383
rect 27755 20380 27767 20383
rect 29012 20380 29040 20479
rect 31478 20476 31484 20488
rect 31536 20476 31542 20528
rect 29273 20451 29331 20457
rect 29273 20417 29285 20451
rect 29319 20448 29331 20451
rect 29362 20448 29368 20460
rect 29319 20420 29368 20448
rect 29319 20417 29331 20420
rect 29273 20411 29331 20417
rect 29362 20408 29368 20420
rect 29420 20408 29426 20460
rect 30116 20420 30788 20448
rect 27755 20352 29040 20380
rect 29181 20383 29239 20389
rect 27755 20349 27767 20352
rect 27709 20343 27767 20349
rect 29181 20349 29193 20383
rect 29227 20349 29239 20383
rect 29181 20343 29239 20349
rect 26384 20284 27292 20312
rect 26384 20272 26390 20284
rect 27430 20272 27436 20324
rect 27488 20272 27494 20324
rect 29196 20312 29224 20343
rect 29638 20340 29644 20392
rect 29696 20340 29702 20392
rect 30116 20380 30144 20420
rect 29748 20352 30144 20380
rect 30561 20383 30619 20389
rect 29748 20321 29776 20352
rect 30561 20349 30573 20383
rect 30607 20380 30619 20383
rect 30650 20380 30656 20392
rect 30607 20352 30656 20380
rect 30607 20349 30619 20352
rect 30561 20343 30619 20349
rect 30650 20340 30656 20352
rect 30708 20340 30714 20392
rect 30760 20389 30788 20420
rect 30926 20408 30932 20460
rect 30984 20448 30990 20460
rect 31297 20451 31355 20457
rect 31297 20448 31309 20451
rect 30984 20420 31309 20448
rect 30984 20408 30990 20420
rect 31297 20417 31309 20420
rect 31343 20417 31355 20451
rect 32217 20451 32275 20457
rect 32217 20448 32229 20451
rect 31297 20411 31355 20417
rect 31680 20420 32229 20448
rect 30745 20383 30803 20389
rect 30745 20349 30757 20383
rect 30791 20380 30803 20383
rect 30834 20380 30840 20392
rect 30791 20352 30840 20380
rect 30791 20349 30803 20352
rect 30745 20343 30803 20349
rect 30834 20340 30840 20352
rect 30892 20340 30898 20392
rect 31018 20340 31024 20392
rect 31076 20340 31082 20392
rect 31386 20340 31392 20392
rect 31444 20380 31450 20392
rect 31680 20380 31708 20420
rect 32217 20417 32229 20420
rect 32263 20417 32275 20451
rect 32217 20411 32275 20417
rect 32493 20451 32551 20457
rect 32493 20417 32505 20451
rect 32539 20448 32551 20451
rect 32582 20448 32588 20460
rect 32539 20420 32588 20448
rect 32539 20417 32551 20420
rect 32493 20411 32551 20417
rect 32582 20408 32588 20420
rect 32640 20408 32646 20460
rect 31444 20352 31708 20380
rect 31444 20340 31450 20352
rect 32030 20340 32036 20392
rect 32088 20340 32094 20392
rect 33870 20380 33876 20392
rect 33626 20352 33876 20380
rect 33870 20340 33876 20352
rect 33928 20340 33934 20392
rect 29733 20315 29791 20321
rect 29733 20312 29745 20315
rect 29196 20284 29745 20312
rect 29733 20281 29745 20284
rect 29779 20281 29791 20315
rect 29733 20275 29791 20281
rect 29914 20272 29920 20324
rect 29972 20321 29978 20324
rect 29972 20315 30007 20321
rect 29995 20281 30007 20315
rect 31404 20312 31432 20340
rect 29972 20275 30007 20281
rect 30576 20284 31432 20312
rect 29972 20272 29978 20275
rect 30576 20256 30604 20284
rect 31570 20272 31576 20324
rect 31628 20272 31634 20324
rect 28629 20247 28687 20253
rect 28629 20244 28641 20247
rect 24780 20216 28641 20244
rect 28629 20213 28641 20216
rect 28675 20244 28687 20247
rect 29822 20244 29828 20256
rect 28675 20216 29828 20244
rect 28675 20213 28687 20216
rect 28629 20207 28687 20213
rect 29822 20204 29828 20216
rect 29880 20204 29886 20256
rect 30098 20204 30104 20256
rect 30156 20204 30162 20256
rect 30558 20204 30564 20256
rect 30616 20204 30622 20256
rect 30742 20204 30748 20256
rect 30800 20244 30806 20256
rect 30929 20247 30987 20253
rect 30929 20244 30941 20247
rect 30800 20216 30941 20244
rect 30800 20204 30806 20216
rect 30929 20213 30941 20216
rect 30975 20213 30987 20247
rect 30929 20207 30987 20213
rect 31018 20204 31024 20256
rect 31076 20244 31082 20256
rect 31481 20247 31539 20253
rect 31481 20244 31493 20247
rect 31076 20216 31493 20244
rect 31076 20204 31082 20216
rect 31481 20213 31493 20216
rect 31527 20244 31539 20247
rect 32048 20244 32076 20340
rect 31527 20216 32076 20244
rect 33965 20247 34023 20253
rect 31527 20213 31539 20216
rect 31481 20207 31539 20213
rect 33965 20213 33977 20247
rect 34011 20244 34023 20247
rect 34011 20216 34376 20244
rect 34011 20213 34023 20216
rect 33965 20207 34023 20213
rect 2760 20154 34316 20176
rect 2760 20102 7210 20154
rect 7262 20102 7274 20154
rect 7326 20102 7338 20154
rect 7390 20102 7402 20154
rect 7454 20102 7466 20154
rect 7518 20102 15099 20154
rect 15151 20102 15163 20154
rect 15215 20102 15227 20154
rect 15279 20102 15291 20154
rect 15343 20102 15355 20154
rect 15407 20102 22988 20154
rect 23040 20102 23052 20154
rect 23104 20102 23116 20154
rect 23168 20102 23180 20154
rect 23232 20102 23244 20154
rect 23296 20102 30877 20154
rect 30929 20102 30941 20154
rect 30993 20102 31005 20154
rect 31057 20102 31069 20154
rect 31121 20102 31133 20154
rect 31185 20102 34316 20154
rect 2760 20080 34316 20102
rect 5261 20043 5319 20049
rect 5261 20040 5273 20043
rect 4172 20012 5273 20040
rect 4172 19972 4200 20012
rect 5261 20009 5273 20012
rect 5307 20009 5319 20043
rect 5261 20003 5319 20009
rect 5350 20000 5356 20052
rect 5408 20040 5414 20052
rect 6181 20043 6239 20049
rect 6181 20040 6193 20043
rect 5408 20012 6193 20040
rect 5408 20000 5414 20012
rect 6181 20009 6193 20012
rect 6227 20009 6239 20043
rect 6181 20003 6239 20009
rect 7650 20000 7656 20052
rect 7708 20000 7714 20052
rect 7745 20043 7803 20049
rect 7745 20009 7757 20043
rect 7791 20040 7803 20043
rect 7926 20040 7932 20052
rect 7791 20012 7932 20040
rect 7791 20009 7803 20012
rect 7745 20003 7803 20009
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 8018 20000 8024 20052
rect 8076 20000 8082 20052
rect 9030 20000 9036 20052
rect 9088 20040 9094 20052
rect 9125 20043 9183 20049
rect 9125 20040 9137 20043
rect 9088 20012 9137 20040
rect 9088 20000 9094 20012
rect 9125 20009 9137 20012
rect 9171 20009 9183 20043
rect 9125 20003 9183 20009
rect 10410 20000 10416 20052
rect 10468 20000 10474 20052
rect 10597 20043 10655 20049
rect 10597 20009 10609 20043
rect 10643 20040 10655 20043
rect 11422 20040 11428 20052
rect 10643 20012 11428 20040
rect 10643 20009 10655 20012
rect 10597 20003 10655 20009
rect 11422 20000 11428 20012
rect 11480 20000 11486 20052
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 11609 20043 11667 20049
rect 11609 20040 11621 20043
rect 11572 20012 11621 20040
rect 11572 20000 11578 20012
rect 11609 20009 11621 20012
rect 11655 20040 11667 20043
rect 12897 20043 12955 20049
rect 11655 20012 12296 20040
rect 11655 20009 11667 20012
rect 11609 20003 11667 20009
rect 4094 19944 4200 19972
rect 4614 19932 4620 19984
rect 4672 19972 4678 19984
rect 4672 19944 6776 19972
rect 4672 19932 4678 19944
rect 4522 19796 4528 19848
rect 4580 19796 4586 19848
rect 4798 19796 4804 19848
rect 4856 19796 4862 19848
rect 3053 19703 3111 19709
rect 3053 19669 3065 19703
rect 3099 19700 3111 19703
rect 4908 19700 4936 19944
rect 5258 19864 5264 19916
rect 5316 19904 5322 19916
rect 5353 19907 5411 19913
rect 5353 19904 5365 19907
rect 5316 19876 5365 19904
rect 5316 19864 5322 19876
rect 5353 19873 5365 19876
rect 5399 19873 5411 19907
rect 5353 19867 5411 19873
rect 5721 19907 5779 19913
rect 5721 19873 5733 19907
rect 5767 19904 5779 19907
rect 5810 19904 5816 19916
rect 5767 19876 5816 19904
rect 5767 19873 5779 19876
rect 5721 19867 5779 19873
rect 5810 19864 5816 19876
rect 5868 19864 5874 19916
rect 5997 19907 6055 19913
rect 5997 19873 6009 19907
rect 6043 19904 6055 19907
rect 6178 19904 6184 19916
rect 6043 19876 6184 19904
rect 6043 19873 6055 19876
rect 5997 19867 6055 19873
rect 6178 19864 6184 19876
rect 6236 19864 6242 19916
rect 6748 19913 6776 19944
rect 6733 19907 6791 19913
rect 6733 19873 6745 19907
rect 6779 19873 6791 19907
rect 6733 19867 6791 19873
rect 5534 19796 5540 19848
rect 5592 19836 5598 19848
rect 5629 19839 5687 19845
rect 5629 19836 5641 19839
rect 5592 19808 5641 19836
rect 5592 19796 5598 19808
rect 5629 19805 5641 19808
rect 5675 19805 5687 19839
rect 5629 19799 5687 19805
rect 6086 19796 6092 19848
rect 6144 19796 6150 19848
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19805 7159 19839
rect 7668 19836 7696 20000
rect 8036 19904 8064 20000
rect 8680 19944 9168 19972
rect 8573 19907 8631 19913
rect 8573 19904 8585 19907
rect 8036 19876 8585 19904
rect 8573 19873 8585 19876
rect 8619 19873 8631 19907
rect 8573 19867 8631 19873
rect 8021 19839 8079 19845
rect 8021 19836 8033 19839
rect 7668 19808 8033 19836
rect 7101 19799 7159 19805
rect 8021 19805 8033 19808
rect 8067 19805 8079 19839
rect 8680 19836 8708 19944
rect 9140 19904 9168 19944
rect 9490 19932 9496 19984
rect 9548 19972 9554 19984
rect 9585 19975 9643 19981
rect 9585 19972 9597 19975
rect 9548 19944 9597 19972
rect 9548 19932 9554 19944
rect 9585 19941 9597 19944
rect 9631 19941 9643 19975
rect 10428 19972 10456 20000
rect 11793 19975 11851 19981
rect 11793 19972 11805 19975
rect 10428 19944 11805 19972
rect 9585 19935 9643 19941
rect 11793 19941 11805 19944
rect 11839 19941 11851 19975
rect 11793 19935 11851 19941
rect 12066 19932 12072 19984
rect 12124 19932 12130 19984
rect 9692 19904 9812 19905
rect 9140 19877 10272 19904
rect 9140 19876 9720 19877
rect 9784 19876 10272 19877
rect 8021 19799 8079 19805
rect 8128 19808 8708 19836
rect 5718 19728 5724 19780
rect 5776 19768 5782 19780
rect 7116 19768 7144 19799
rect 5776 19740 7144 19768
rect 5776 19728 5782 19740
rect 7650 19728 7656 19780
rect 7708 19768 7714 19780
rect 8128 19768 8156 19808
rect 9030 19796 9036 19848
rect 9088 19796 9094 19848
rect 10244 19836 10272 19876
rect 10318 19864 10324 19916
rect 10376 19904 10382 19916
rect 10413 19907 10471 19913
rect 10413 19904 10425 19907
rect 10376 19876 10425 19904
rect 10376 19864 10382 19876
rect 10413 19873 10425 19876
rect 10459 19873 10471 19907
rect 10413 19867 10471 19873
rect 10502 19864 10508 19916
rect 10560 19864 10566 19916
rect 10870 19864 10876 19916
rect 10928 19864 10934 19916
rect 10962 19864 10968 19916
rect 11020 19864 11026 19916
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 11379 19902 11560 19904
rect 11379 19876 11589 19902
rect 11379 19873 11391 19876
rect 11532 19874 11589 19876
rect 11333 19867 11391 19873
rect 10520 19836 10548 19864
rect 10244 19808 10548 19836
rect 10778 19796 10784 19848
rect 10836 19836 10842 19848
rect 11561 19836 11589 19874
rect 11698 19864 11704 19916
rect 11756 19864 11762 19916
rect 12268 19913 12296 20012
rect 12897 20009 12909 20043
rect 12943 20040 12955 20043
rect 12986 20040 12992 20052
rect 12943 20012 12992 20040
rect 12943 20009 12955 20012
rect 12897 20003 12955 20009
rect 12986 20000 12992 20012
rect 13044 20000 13050 20052
rect 13357 20043 13415 20049
rect 13357 20009 13369 20043
rect 13403 20040 13415 20043
rect 13630 20040 13636 20052
rect 13403 20012 13636 20040
rect 13403 20009 13415 20012
rect 13357 20003 13415 20009
rect 13630 20000 13636 20012
rect 13688 20000 13694 20052
rect 13725 20043 13783 20049
rect 13725 20009 13737 20043
rect 13771 20040 13783 20043
rect 15473 20043 15531 20049
rect 13771 20012 14044 20040
rect 13771 20009 13783 20012
rect 13725 20003 13783 20009
rect 14016 19984 14044 20012
rect 15473 20009 15485 20043
rect 15519 20040 15531 20043
rect 15562 20040 15568 20052
rect 15519 20012 15568 20040
rect 15519 20009 15531 20012
rect 15473 20003 15531 20009
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 16022 20000 16028 20052
rect 16080 20040 16086 20052
rect 16301 20043 16359 20049
rect 16301 20040 16313 20043
rect 16080 20012 16313 20040
rect 16080 20000 16086 20012
rect 16301 20009 16313 20012
rect 16347 20009 16359 20043
rect 16301 20003 16359 20009
rect 16758 20000 16764 20052
rect 16816 20000 16822 20052
rect 17034 20000 17040 20052
rect 17092 20000 17098 20052
rect 18877 20043 18935 20049
rect 18877 20009 18889 20043
rect 18923 20040 18935 20043
rect 18966 20040 18972 20052
rect 18923 20012 18972 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 18966 20000 18972 20012
rect 19024 20040 19030 20052
rect 19150 20040 19156 20052
rect 19024 20012 19156 20040
rect 19024 20000 19030 20012
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 19337 20043 19395 20049
rect 19337 20009 19349 20043
rect 19383 20040 19395 20043
rect 20898 20040 20904 20052
rect 19383 20012 20904 20040
rect 19383 20009 19395 20012
rect 19337 20003 19395 20009
rect 20898 20000 20904 20012
rect 20956 20040 20962 20052
rect 21266 20040 21272 20052
rect 20956 20012 21272 20040
rect 20956 20000 20962 20012
rect 21266 20000 21272 20012
rect 21324 20000 21330 20052
rect 22186 20040 22192 20052
rect 21744 20012 22192 20040
rect 13814 19932 13820 19984
rect 13872 19932 13878 19984
rect 13998 19932 14004 19984
rect 14056 19932 14062 19984
rect 14182 19932 14188 19984
rect 14240 19932 14246 19984
rect 16390 19932 16396 19984
rect 16448 19972 16454 19984
rect 16669 19975 16727 19981
rect 16669 19972 16681 19975
rect 16448 19944 16681 19972
rect 16448 19932 16454 19944
rect 16669 19941 16681 19944
rect 16715 19972 16727 19975
rect 17052 19972 17080 20000
rect 19426 19972 19432 19984
rect 16715 19944 17080 19972
rect 18064 19944 19432 19972
rect 16715 19941 16727 19944
rect 16669 19935 16727 19941
rect 12253 19907 12311 19913
rect 12253 19873 12265 19907
rect 12299 19873 12311 19907
rect 12253 19867 12311 19873
rect 12342 19864 12348 19916
rect 12400 19864 12406 19916
rect 12989 19907 13047 19913
rect 12989 19873 13001 19907
rect 13035 19904 13047 19907
rect 13538 19904 13544 19916
rect 13035 19876 13544 19904
rect 13035 19873 13047 19876
rect 12989 19867 13047 19873
rect 13538 19864 13544 19876
rect 13596 19864 13602 19916
rect 17405 19907 17463 19913
rect 17405 19904 17417 19907
rect 13832 19876 14044 19904
rect 10836 19808 11468 19836
rect 11561 19808 11652 19836
rect 10836 19796 10842 19808
rect 9585 19771 9643 19777
rect 7708 19740 8156 19768
rect 8312 19740 8984 19768
rect 7708 19728 7714 19740
rect 3099 19672 4936 19700
rect 3099 19669 3111 19672
rect 3053 19663 3111 19669
rect 4982 19660 4988 19712
rect 5040 19700 5046 19712
rect 5445 19703 5503 19709
rect 5445 19700 5457 19703
rect 5040 19672 5457 19700
rect 5040 19660 5046 19672
rect 5445 19669 5457 19672
rect 5491 19669 5503 19703
rect 5445 19663 5503 19669
rect 5810 19660 5816 19712
rect 5868 19700 5874 19712
rect 7668 19700 7696 19728
rect 8312 19712 8340 19740
rect 5868 19672 7696 19700
rect 5868 19660 5874 19672
rect 8294 19660 8300 19712
rect 8352 19660 8358 19712
rect 8386 19660 8392 19712
rect 8444 19700 8450 19712
rect 8849 19703 8907 19709
rect 8849 19700 8861 19703
rect 8444 19672 8861 19700
rect 8444 19660 8450 19672
rect 8849 19669 8861 19672
rect 8895 19669 8907 19703
rect 8956 19700 8984 19740
rect 9585 19737 9597 19771
rect 9631 19768 9643 19771
rect 10042 19768 10048 19780
rect 9631 19740 10048 19768
rect 9631 19737 9643 19740
rect 9585 19731 9643 19737
rect 10042 19728 10048 19740
rect 10100 19728 10106 19780
rect 10870 19728 10876 19780
rect 10928 19768 10934 19780
rect 11057 19771 11115 19777
rect 11057 19768 11069 19771
rect 10928 19740 11069 19768
rect 10928 19728 10934 19740
rect 11057 19737 11069 19740
rect 11103 19737 11115 19771
rect 11440 19768 11468 19808
rect 11624 19768 11652 19808
rect 12158 19796 12164 19848
rect 12216 19836 12222 19848
rect 13832 19836 13860 19876
rect 12216 19808 13860 19836
rect 12216 19796 12222 19808
rect 13906 19796 13912 19848
rect 13964 19796 13970 19848
rect 11977 19771 12035 19777
rect 11977 19768 11989 19771
rect 11440 19740 11589 19768
rect 11624 19740 11989 19768
rect 11057 19731 11115 19737
rect 9769 19703 9827 19709
rect 9769 19700 9781 19703
rect 8956 19672 9781 19700
rect 8849 19663 8907 19669
rect 9769 19669 9781 19672
rect 9815 19669 9827 19703
rect 9769 19663 9827 19669
rect 10686 19660 10692 19712
rect 10744 19700 10750 19712
rect 11149 19703 11207 19709
rect 11149 19700 11161 19703
rect 10744 19672 11161 19700
rect 10744 19660 10750 19672
rect 11149 19669 11161 19672
rect 11195 19669 11207 19703
rect 11149 19663 11207 19669
rect 11422 19660 11428 19712
rect 11480 19660 11486 19712
rect 11561 19700 11589 19740
rect 11977 19737 11989 19740
rect 12023 19768 12035 19771
rect 13262 19768 13268 19780
rect 12023 19740 13268 19768
rect 12023 19737 12035 19740
rect 11977 19731 12035 19737
rect 13262 19728 13268 19740
rect 13320 19728 13326 19780
rect 14016 19768 14044 19876
rect 16776 19876 17417 19904
rect 16482 19796 16488 19848
rect 16540 19836 16546 19848
rect 16776 19836 16804 19876
rect 17405 19873 17417 19876
rect 17451 19904 17463 19907
rect 17954 19904 17960 19916
rect 17451 19876 17960 19904
rect 17451 19873 17463 19876
rect 17405 19867 17463 19873
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 16540 19808 16804 19836
rect 16945 19839 17003 19845
rect 16540 19796 16546 19808
rect 16945 19805 16957 19839
rect 16991 19836 17003 19839
rect 17218 19836 17224 19848
rect 16991 19808 17224 19836
rect 16991 19805 17003 19808
rect 16945 19799 17003 19805
rect 17218 19796 17224 19808
rect 17276 19796 17282 19848
rect 18064 19768 18092 19944
rect 19426 19932 19432 19944
rect 19484 19932 19490 19984
rect 19886 19932 19892 19984
rect 19944 19932 19950 19984
rect 19981 19975 20039 19981
rect 19981 19941 19993 19975
rect 20027 19972 20039 19975
rect 20441 19975 20499 19981
rect 20441 19972 20453 19975
rect 20027 19944 20453 19972
rect 20027 19941 20039 19944
rect 19981 19935 20039 19941
rect 20441 19941 20453 19944
rect 20487 19972 20499 19975
rect 20530 19972 20536 19984
rect 20487 19944 20536 19972
rect 20487 19941 20499 19944
rect 20441 19935 20499 19941
rect 20530 19932 20536 19944
rect 20588 19932 20594 19984
rect 21744 19972 21772 20012
rect 22186 20000 22192 20012
rect 22244 20000 22250 20052
rect 22833 20043 22891 20049
rect 22833 20009 22845 20043
rect 22879 20040 22891 20043
rect 26326 20040 26332 20052
rect 22879 20012 26332 20040
rect 22879 20009 22891 20012
rect 22833 20003 22891 20009
rect 26326 20000 26332 20012
rect 26384 20000 26390 20052
rect 27065 20043 27123 20049
rect 27065 20009 27077 20043
rect 27111 20040 27123 20043
rect 27430 20040 27436 20052
rect 27111 20012 27436 20040
rect 27111 20009 27123 20012
rect 27065 20003 27123 20009
rect 27430 20000 27436 20012
rect 27488 20000 27494 20052
rect 28905 20043 28963 20049
rect 28905 20009 28917 20043
rect 28951 20009 28963 20043
rect 28905 20003 28963 20009
rect 20916 19944 21772 19972
rect 18325 19907 18383 19913
rect 18325 19873 18337 19907
rect 18371 19873 18383 19907
rect 18325 19867 18383 19873
rect 18345 19836 18373 19867
rect 18690 19864 18696 19916
rect 18748 19904 18754 19916
rect 18969 19907 19027 19913
rect 18969 19904 18981 19907
rect 18748 19876 18981 19904
rect 18748 19864 18754 19876
rect 18969 19873 18981 19876
rect 19015 19873 19027 19907
rect 18969 19867 19027 19873
rect 19150 19864 19156 19916
rect 19208 19904 19214 19916
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 19208 19876 19625 19904
rect 19208 19864 19214 19876
rect 19613 19873 19625 19876
rect 19659 19873 19671 19907
rect 19613 19867 19671 19873
rect 19705 19907 19763 19913
rect 19705 19873 19717 19907
rect 19751 19904 19763 19907
rect 19904 19904 19932 19932
rect 20916 19913 20944 19944
rect 22094 19932 22100 19984
rect 22152 19932 22158 19984
rect 24670 19932 24676 19984
rect 24728 19972 24734 19984
rect 24728 19944 25268 19972
rect 24728 19932 24734 19944
rect 20165 19907 20223 19913
rect 20165 19904 20177 19907
rect 19751 19876 19932 19904
rect 19996 19876 20177 19904
rect 19751 19873 19763 19876
rect 19705 19867 19763 19873
rect 19996 19848 20024 19876
rect 20165 19873 20177 19876
rect 20211 19904 20223 19907
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20211 19876 20913 19904
rect 20211 19873 20223 19876
rect 20165 19867 20223 19873
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 23109 19907 23167 19913
rect 23109 19873 23121 19907
rect 23155 19873 23167 19907
rect 23109 19867 23167 19873
rect 23293 19907 23351 19913
rect 23293 19873 23305 19907
rect 23339 19904 23351 19907
rect 23658 19904 23664 19916
rect 23339 19876 23664 19904
rect 23339 19873 23351 19876
rect 23293 19867 23351 19873
rect 18414 19836 18420 19848
rect 18345 19808 18420 19836
rect 18414 19796 18420 19808
rect 18472 19796 18478 19848
rect 18601 19839 18659 19845
rect 18601 19805 18613 19839
rect 18647 19805 18659 19839
rect 18601 19799 18659 19805
rect 14016 19740 18092 19768
rect 18230 19728 18236 19780
rect 18288 19768 18294 19780
rect 18616 19768 18644 19799
rect 19058 19796 19064 19848
rect 19116 19796 19122 19848
rect 19978 19796 19984 19848
rect 20036 19796 20042 19848
rect 20070 19796 20076 19848
rect 20128 19796 20134 19848
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21085 19839 21143 19845
rect 21085 19836 21097 19839
rect 21048 19808 21097 19836
rect 21048 19796 21054 19808
rect 21085 19805 21097 19808
rect 21131 19836 21143 19839
rect 21131 19808 21220 19836
rect 21131 19805 21143 19808
rect 21085 19799 21143 19805
rect 18288 19740 19196 19768
rect 18288 19728 18294 19740
rect 12069 19703 12127 19709
rect 12069 19700 12081 19703
rect 11561 19672 12081 19700
rect 12069 19669 12081 19672
rect 12115 19669 12127 19703
rect 12069 19663 12127 19669
rect 12526 19660 12532 19712
rect 12584 19660 12590 19712
rect 17034 19660 17040 19712
rect 17092 19700 17098 19712
rect 17310 19700 17316 19712
rect 17092 19672 17316 19700
rect 17092 19660 17098 19672
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 17497 19703 17555 19709
rect 17497 19700 17509 19703
rect 17460 19672 17509 19700
rect 17460 19660 17466 19672
rect 17497 19669 17509 19672
rect 17543 19669 17555 19703
rect 17497 19663 17555 19669
rect 17954 19660 17960 19712
rect 18012 19700 18018 19712
rect 18049 19703 18107 19709
rect 18049 19700 18061 19703
rect 18012 19672 18061 19700
rect 18012 19660 18018 19672
rect 18049 19669 18061 19672
rect 18095 19669 18107 19703
rect 18049 19663 18107 19669
rect 18322 19660 18328 19712
rect 18380 19700 18386 19712
rect 19168 19709 19196 19740
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 19429 19771 19487 19777
rect 19429 19768 19441 19771
rect 19300 19740 19441 19768
rect 19300 19728 19306 19740
rect 19429 19737 19441 19740
rect 19475 19737 19487 19771
rect 19429 19731 19487 19737
rect 18417 19703 18475 19709
rect 18417 19700 18429 19703
rect 18380 19672 18429 19700
rect 18380 19660 18386 19672
rect 18417 19669 18429 19672
rect 18463 19669 18475 19703
rect 18417 19663 18475 19669
rect 19153 19703 19211 19709
rect 19153 19669 19165 19703
rect 19199 19700 19211 19703
rect 19886 19700 19892 19712
rect 19199 19672 19892 19700
rect 19199 19669 19211 19672
rect 19153 19663 19211 19669
rect 19886 19660 19892 19672
rect 19944 19660 19950 19712
rect 21192 19700 21220 19808
rect 21358 19796 21364 19848
rect 21416 19796 21422 19848
rect 22554 19728 22560 19780
rect 22612 19728 22618 19780
rect 23124 19768 23152 19867
rect 23658 19864 23664 19876
rect 23716 19864 23722 19916
rect 23842 19864 23848 19916
rect 23900 19864 23906 19916
rect 25240 19913 25268 19944
rect 25314 19932 25320 19984
rect 25372 19972 25378 19984
rect 27985 19975 28043 19981
rect 25372 19944 27292 19972
rect 25372 19932 25378 19944
rect 25225 19907 25283 19913
rect 25225 19873 25237 19907
rect 25271 19873 25283 19907
rect 25225 19867 25283 19873
rect 25682 19864 25688 19916
rect 25740 19904 25746 19916
rect 26053 19907 26111 19913
rect 26053 19904 26065 19907
rect 25740 19876 26065 19904
rect 25740 19864 25746 19876
rect 26053 19873 26065 19876
rect 26099 19873 26111 19907
rect 26053 19867 26111 19873
rect 26234 19864 26240 19916
rect 26292 19904 26298 19916
rect 26786 19904 26792 19916
rect 26292 19876 26792 19904
rect 26292 19864 26298 19876
rect 26786 19864 26792 19876
rect 26844 19864 26850 19916
rect 27264 19913 27292 19944
rect 27985 19941 27997 19975
rect 28031 19972 28043 19975
rect 28920 19972 28948 20003
rect 30742 20000 30748 20052
rect 30800 20000 30806 20052
rect 32306 20000 32312 20052
rect 32364 20000 32370 20052
rect 32398 20000 32404 20052
rect 32456 20040 32462 20052
rect 33045 20043 33103 20049
rect 33045 20040 33057 20043
rect 32456 20012 33057 20040
rect 32456 20000 32462 20012
rect 33045 20009 33057 20012
rect 33091 20009 33103 20043
rect 33045 20003 33103 20009
rect 33137 20043 33195 20049
rect 33137 20009 33149 20043
rect 33183 20040 33195 20043
rect 34348 20040 34376 20216
rect 33183 20012 34376 20040
rect 33183 20009 33195 20012
rect 33137 20003 33195 20009
rect 29362 19972 29368 19984
rect 28031 19944 28948 19972
rect 29012 19944 29368 19972
rect 28031 19941 28043 19944
rect 27985 19935 28043 19941
rect 27249 19907 27307 19913
rect 27249 19873 27261 19907
rect 27295 19873 27307 19907
rect 27249 19867 27307 19873
rect 27338 19864 27344 19916
rect 27396 19864 27402 19916
rect 27709 19907 27767 19913
rect 27709 19873 27721 19907
rect 27755 19904 27767 19907
rect 27890 19904 27896 19916
rect 27755 19876 27896 19904
rect 27755 19873 27767 19876
rect 27709 19867 27767 19873
rect 27890 19864 27896 19876
rect 27948 19864 27954 19916
rect 28261 19907 28319 19913
rect 28261 19873 28273 19907
rect 28307 19904 28319 19907
rect 29012 19904 29040 19944
rect 29362 19932 29368 19944
rect 29420 19932 29426 19984
rect 29549 19975 29607 19981
rect 29549 19941 29561 19975
rect 29595 19972 29607 19975
rect 29638 19972 29644 19984
rect 29595 19944 29644 19972
rect 29595 19941 29607 19944
rect 29549 19935 29607 19941
rect 29638 19932 29644 19944
rect 29696 19932 29702 19984
rect 30760 19972 30788 20000
rect 30837 19975 30895 19981
rect 30837 19972 30849 19975
rect 30760 19944 30849 19972
rect 30837 19941 30849 19944
rect 30883 19941 30895 19975
rect 32493 19975 32551 19981
rect 32493 19972 32505 19975
rect 32062 19944 32505 19972
rect 30837 19935 30895 19941
rect 32493 19941 32505 19944
rect 32539 19941 32551 19975
rect 32493 19935 32551 19941
rect 32766 19932 32772 19984
rect 32824 19972 32830 19984
rect 33152 19972 33180 20003
rect 32824 19944 33180 19972
rect 32824 19932 32830 19944
rect 28307 19876 29040 19904
rect 29089 19907 29147 19913
rect 28307 19873 28319 19876
rect 28261 19867 28319 19873
rect 29089 19873 29101 19907
rect 29135 19904 29147 19907
rect 29730 19904 29736 19916
rect 29135 19876 29736 19904
rect 29135 19873 29147 19876
rect 29089 19867 29147 19873
rect 29730 19864 29736 19876
rect 29788 19864 29794 19916
rect 30558 19864 30564 19916
rect 30616 19864 30622 19916
rect 32585 19907 32643 19913
rect 32585 19873 32597 19907
rect 32631 19904 32643 19907
rect 33134 19904 33140 19916
rect 32631 19876 33140 19904
rect 32631 19873 32643 19876
rect 32585 19867 32643 19873
rect 33134 19864 33140 19876
rect 33192 19864 33198 19916
rect 23201 19839 23259 19845
rect 23201 19805 23213 19839
rect 23247 19836 23259 19839
rect 23474 19836 23480 19848
rect 23247 19808 23480 19836
rect 23247 19805 23259 19808
rect 23201 19799 23259 19805
rect 23474 19796 23480 19808
rect 23532 19796 23538 19848
rect 25961 19839 26019 19845
rect 25961 19836 25973 19839
rect 23952 19808 25973 19836
rect 23566 19768 23572 19780
rect 23124 19740 23572 19768
rect 23566 19728 23572 19740
rect 23624 19728 23630 19780
rect 22572 19700 22600 19728
rect 21192 19672 22600 19700
rect 23477 19703 23535 19709
rect 23477 19669 23489 19703
rect 23523 19700 23535 19703
rect 23952 19700 23980 19808
rect 25961 19805 25973 19808
rect 26007 19836 26019 19839
rect 27356 19836 27384 19864
rect 26007 19808 27384 19836
rect 27433 19839 27491 19845
rect 26007 19805 26019 19808
rect 25961 19799 26019 19805
rect 27433 19805 27445 19839
rect 27479 19836 27491 19839
rect 28074 19836 28080 19848
rect 27479 19808 28080 19836
rect 27479 19805 27491 19808
rect 27433 19799 27491 19805
rect 28074 19796 28080 19808
rect 28132 19796 28138 19848
rect 28169 19839 28227 19845
rect 28169 19805 28181 19839
rect 28215 19836 28227 19839
rect 28994 19836 29000 19848
rect 28215 19808 29000 19836
rect 28215 19805 28227 19808
rect 28169 19799 28227 19805
rect 28994 19796 29000 19808
rect 29052 19796 29058 19848
rect 29273 19839 29331 19845
rect 29273 19805 29285 19839
rect 29319 19836 29331 19839
rect 32306 19836 32312 19848
rect 29319 19808 32312 19836
rect 29319 19805 29331 19808
rect 29273 19799 29331 19805
rect 32306 19796 32312 19808
rect 32364 19796 32370 19848
rect 33042 19796 33048 19848
rect 33100 19836 33106 19848
rect 33229 19839 33287 19845
rect 33229 19836 33241 19839
rect 33100 19808 33241 19836
rect 33100 19796 33106 19808
rect 33229 19805 33241 19808
rect 33275 19805 33287 19839
rect 33229 19799 33287 19805
rect 33318 19796 33324 19848
rect 33376 19796 33382 19848
rect 26050 19728 26056 19780
rect 26108 19768 26114 19780
rect 27062 19768 27068 19780
rect 26108 19740 27068 19768
rect 26108 19728 26114 19740
rect 27062 19728 27068 19740
rect 27120 19728 27126 19780
rect 29638 19768 29644 19780
rect 27540 19740 29644 19768
rect 27540 19712 27568 19740
rect 29638 19728 29644 19740
rect 29696 19728 29702 19780
rect 32677 19771 32735 19777
rect 32677 19737 32689 19771
rect 32723 19768 32735 19771
rect 33336 19768 33364 19796
rect 32723 19740 33364 19768
rect 32723 19737 32735 19740
rect 32677 19731 32735 19737
rect 23523 19672 23980 19700
rect 23523 19669 23535 19672
rect 23477 19663 23535 19669
rect 24946 19660 24952 19712
rect 25004 19709 25010 19712
rect 25004 19703 25019 19709
rect 25007 19669 25019 19703
rect 25004 19663 25019 19669
rect 25004 19660 25010 19663
rect 25774 19660 25780 19712
rect 25832 19700 25838 19712
rect 26145 19703 26203 19709
rect 26145 19700 26157 19703
rect 25832 19672 26157 19700
rect 25832 19660 25838 19672
rect 26145 19669 26157 19672
rect 26191 19669 26203 19703
rect 26145 19663 26203 19669
rect 26602 19660 26608 19712
rect 26660 19700 26666 19712
rect 27249 19703 27307 19709
rect 27249 19700 27261 19703
rect 26660 19672 27261 19700
rect 26660 19660 26666 19672
rect 27249 19669 27261 19672
rect 27295 19669 27307 19703
rect 27249 19663 27307 19669
rect 27522 19660 27528 19712
rect 27580 19660 27586 19712
rect 27982 19660 27988 19712
rect 28040 19660 28046 19712
rect 28445 19703 28503 19709
rect 28445 19669 28457 19703
rect 28491 19700 28503 19703
rect 28994 19700 29000 19712
rect 28491 19672 29000 19700
rect 28491 19669 28503 19672
rect 28445 19663 28503 19669
rect 28994 19660 29000 19672
rect 29052 19660 29058 19712
rect 29457 19703 29515 19709
rect 29457 19669 29469 19703
rect 29503 19700 29515 19703
rect 30650 19700 30656 19712
rect 29503 19672 30656 19700
rect 29503 19669 29515 19672
rect 29457 19663 29515 19669
rect 30650 19660 30656 19672
rect 30708 19660 30714 19712
rect 2760 19610 34316 19632
rect 2760 19558 6550 19610
rect 6602 19558 6614 19610
rect 6666 19558 6678 19610
rect 6730 19558 6742 19610
rect 6794 19558 6806 19610
rect 6858 19558 14439 19610
rect 14491 19558 14503 19610
rect 14555 19558 14567 19610
rect 14619 19558 14631 19610
rect 14683 19558 14695 19610
rect 14747 19558 22328 19610
rect 22380 19558 22392 19610
rect 22444 19558 22456 19610
rect 22508 19558 22520 19610
rect 22572 19558 22584 19610
rect 22636 19558 30217 19610
rect 30269 19558 30281 19610
rect 30333 19558 30345 19610
rect 30397 19558 30409 19610
rect 30461 19558 30473 19610
rect 30525 19558 34316 19610
rect 2760 19536 34316 19558
rect 5077 19499 5135 19505
rect 5077 19465 5089 19499
rect 5123 19496 5135 19499
rect 5166 19496 5172 19508
rect 5123 19468 5172 19496
rect 5123 19465 5135 19468
rect 5077 19459 5135 19465
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 5261 19499 5319 19505
rect 5261 19465 5273 19499
rect 5307 19496 5319 19499
rect 5534 19496 5540 19508
rect 5307 19468 5540 19496
rect 5307 19465 5319 19468
rect 5261 19459 5319 19465
rect 5534 19456 5540 19468
rect 5592 19456 5598 19508
rect 6996 19499 7054 19505
rect 6996 19465 7008 19499
rect 7042 19496 7054 19499
rect 8573 19499 8631 19505
rect 8573 19496 8585 19499
rect 7042 19468 8585 19496
rect 7042 19465 7054 19468
rect 6996 19459 7054 19465
rect 8573 19465 8585 19468
rect 8619 19465 8631 19499
rect 8573 19459 8631 19465
rect 10229 19499 10287 19505
rect 10229 19465 10241 19499
rect 10275 19496 10287 19499
rect 10962 19496 10968 19508
rect 10275 19468 10968 19496
rect 10275 19465 10287 19468
rect 10229 19459 10287 19465
rect 10962 19456 10968 19468
rect 11020 19456 11026 19508
rect 11330 19456 11336 19508
rect 11388 19456 11394 19508
rect 13262 19456 13268 19508
rect 13320 19456 13326 19508
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 14277 19499 14335 19505
rect 14277 19496 14289 19499
rect 13872 19468 14289 19496
rect 13872 19456 13878 19468
rect 14277 19465 14289 19468
rect 14323 19465 14335 19499
rect 14277 19459 14335 19465
rect 15470 19456 15476 19508
rect 15528 19496 15534 19508
rect 15841 19499 15899 19505
rect 15841 19496 15853 19499
rect 15528 19468 15853 19496
rect 15528 19456 15534 19468
rect 15841 19465 15853 19468
rect 15887 19465 15899 19499
rect 15841 19459 15899 19465
rect 16301 19499 16359 19505
rect 16301 19465 16313 19499
rect 16347 19496 16359 19499
rect 16390 19496 16396 19508
rect 16347 19468 16396 19496
rect 16347 19465 16359 19468
rect 16301 19459 16359 19465
rect 16390 19456 16396 19468
rect 16448 19456 16454 19508
rect 16669 19499 16727 19505
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 17037 19499 17095 19505
rect 17037 19496 17049 19499
rect 16715 19468 17049 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 17037 19465 17049 19468
rect 17083 19496 17095 19499
rect 17218 19496 17224 19508
rect 17083 19468 17224 19496
rect 17083 19465 17095 19468
rect 17037 19459 17095 19465
rect 5626 19428 5632 19440
rect 5092 19400 5632 19428
rect 3234 19252 3240 19304
rect 3292 19252 3298 19304
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 4614 19292 4620 19304
rect 4479 19264 4620 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4614 19252 4620 19264
rect 4672 19252 4678 19304
rect 5092 19301 5120 19400
rect 5626 19388 5632 19400
rect 5684 19428 5690 19440
rect 6730 19428 6736 19440
rect 5684 19400 6736 19428
rect 5684 19388 5690 19400
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 8110 19388 8116 19440
rect 8168 19428 8174 19440
rect 16684 19428 16712 19459
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 21174 19456 21180 19508
rect 21232 19496 21238 19508
rect 21450 19496 21456 19508
rect 21232 19468 21456 19496
rect 21232 19456 21238 19468
rect 21450 19456 21456 19468
rect 21508 19456 21514 19508
rect 22094 19456 22100 19508
rect 22152 19456 22158 19508
rect 24946 19456 24952 19508
rect 25004 19496 25010 19508
rect 25041 19499 25099 19505
rect 25041 19496 25053 19499
rect 25004 19468 25053 19496
rect 25004 19456 25010 19468
rect 25041 19465 25053 19468
rect 25087 19465 25099 19499
rect 25041 19459 25099 19465
rect 26418 19456 26424 19508
rect 26476 19496 26482 19508
rect 26786 19496 26792 19508
rect 26476 19468 26792 19496
rect 26476 19456 26482 19468
rect 26786 19456 26792 19468
rect 26844 19496 26850 19508
rect 27525 19499 27583 19505
rect 27525 19496 27537 19499
rect 26844 19468 27537 19496
rect 26844 19456 26850 19468
rect 27525 19465 27537 19468
rect 27571 19465 27583 19499
rect 27525 19459 27583 19465
rect 29178 19456 29184 19508
rect 29236 19496 29242 19508
rect 30098 19496 30104 19508
rect 29236 19468 30104 19496
rect 29236 19456 29242 19468
rect 30098 19456 30104 19468
rect 30156 19456 30162 19508
rect 8168 19400 16712 19428
rect 8168 19388 8174 19400
rect 26326 19388 26332 19440
rect 26384 19428 26390 19440
rect 26694 19428 26700 19440
rect 26384 19400 26700 19428
rect 26384 19388 26390 19400
rect 26694 19388 26700 19400
rect 26752 19388 26758 19440
rect 28074 19388 28080 19440
rect 28132 19428 28138 19440
rect 28810 19428 28816 19440
rect 28132 19400 28816 19428
rect 28132 19388 28138 19400
rect 28810 19388 28816 19400
rect 28868 19428 28874 19440
rect 28905 19431 28963 19437
rect 28905 19428 28917 19431
rect 28868 19400 28917 19428
rect 28868 19388 28874 19400
rect 28905 19397 28917 19400
rect 28951 19397 28963 19431
rect 28905 19391 28963 19397
rect 29454 19388 29460 19440
rect 29512 19428 29518 19440
rect 29641 19431 29699 19437
rect 29641 19428 29653 19431
rect 29512 19400 29653 19428
rect 29512 19388 29518 19400
rect 29641 19397 29653 19400
rect 29687 19428 29699 19431
rect 29914 19428 29920 19440
rect 29687 19400 29920 19428
rect 29687 19397 29699 19400
rect 29641 19391 29699 19397
rect 29914 19388 29920 19400
rect 29972 19388 29978 19440
rect 5258 19320 5264 19372
rect 5316 19320 5322 19372
rect 5718 19320 5724 19372
rect 5776 19360 5782 19372
rect 5997 19363 6055 19369
rect 5997 19360 6009 19363
rect 5776 19332 6009 19360
rect 5776 19320 5782 19332
rect 5997 19329 6009 19332
rect 6043 19329 6055 19363
rect 7098 19360 7104 19372
rect 5997 19323 6055 19329
rect 6748 19332 7104 19360
rect 4709 19295 4767 19301
rect 4709 19261 4721 19295
rect 4755 19292 4767 19295
rect 5077 19295 5135 19301
rect 4755 19264 5028 19292
rect 4755 19261 4767 19264
rect 4709 19255 4767 19261
rect 5000 19224 5028 19264
rect 5077 19261 5089 19295
rect 5123 19261 5135 19295
rect 5276 19292 5304 19320
rect 6748 19301 6776 19332
rect 7098 19320 7104 19332
rect 7156 19320 7162 19372
rect 9766 19320 9772 19372
rect 9824 19360 9830 19372
rect 9861 19363 9919 19369
rect 9861 19360 9873 19363
rect 9824 19332 9873 19360
rect 9824 19320 9830 19332
rect 9861 19329 9873 19332
rect 9907 19329 9919 19363
rect 9861 19323 9919 19329
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5276 19264 5641 19292
rect 5077 19255 5135 19261
rect 5629 19261 5641 19264
rect 5675 19261 5687 19295
rect 5629 19255 5687 19261
rect 6733 19295 6791 19301
rect 6733 19261 6745 19295
rect 6779 19261 6791 19295
rect 6733 19255 6791 19261
rect 9122 19252 9128 19304
rect 9180 19252 9186 19304
rect 5000 19196 7420 19224
rect 5534 19116 5540 19168
rect 5592 19116 5598 19168
rect 6641 19159 6699 19165
rect 6641 19125 6653 19159
rect 6687 19156 6699 19159
rect 6914 19156 6920 19168
rect 6687 19128 6920 19156
rect 6687 19125 6699 19128
rect 6641 19119 6699 19125
rect 6914 19116 6920 19128
rect 6972 19116 6978 19168
rect 7392 19156 7420 19196
rect 7742 19184 7748 19236
rect 7800 19184 7806 19236
rect 8570 19224 8576 19236
rect 8404 19196 8576 19224
rect 8404 19156 8432 19196
rect 8570 19184 8576 19196
rect 8628 19224 8634 19236
rect 9490 19224 9496 19236
rect 8628 19196 9496 19224
rect 8628 19184 8634 19196
rect 9490 19184 9496 19196
rect 9548 19184 9554 19236
rect 9876 19224 9904 19323
rect 10778 19320 10784 19372
rect 10836 19360 10842 19372
rect 11333 19363 11391 19369
rect 11333 19360 11345 19363
rect 10836 19332 11345 19360
rect 10836 19320 10842 19332
rect 11333 19329 11345 19332
rect 11379 19360 11391 19363
rect 11701 19363 11759 19369
rect 11701 19360 11713 19363
rect 11379 19332 11713 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 11701 19329 11713 19332
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11974 19320 11980 19372
rect 12032 19320 12038 19372
rect 12526 19320 12532 19372
rect 12584 19360 12590 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12584 19332 13001 19360
rect 12584 19320 12590 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13446 19320 13452 19372
rect 13504 19360 13510 19372
rect 13633 19363 13691 19369
rect 13633 19360 13645 19363
rect 13504 19332 13645 19360
rect 13504 19320 13510 19332
rect 13633 19329 13645 19332
rect 13679 19329 13691 19363
rect 13998 19360 14004 19372
rect 13633 19323 13691 19329
rect 13740 19332 14004 19360
rect 9950 19252 9956 19304
rect 10008 19292 10014 19304
rect 10597 19295 10655 19301
rect 10597 19292 10609 19295
rect 10008 19264 10609 19292
rect 10008 19252 10014 19264
rect 10597 19261 10609 19264
rect 10643 19261 10655 19295
rect 10597 19255 10655 19261
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 11146 19292 11152 19304
rect 10735 19264 11152 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 11146 19252 11152 19264
rect 11204 19292 11210 19304
rect 11241 19295 11299 19301
rect 11241 19292 11253 19295
rect 11204 19264 11253 19292
rect 11204 19252 11210 19264
rect 11241 19261 11253 19264
rect 11287 19261 11299 19295
rect 11606 19292 11612 19304
rect 11241 19255 11299 19261
rect 11348 19264 11612 19292
rect 11348 19236 11376 19264
rect 11606 19252 11612 19264
rect 11664 19292 11670 19304
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11664 19264 11805 19292
rect 11664 19252 11670 19264
rect 11793 19261 11805 19264
rect 11839 19261 11851 19295
rect 11793 19255 11851 19261
rect 9876 19196 11192 19224
rect 7392 19128 8432 19156
rect 8478 19116 8484 19168
rect 8536 19116 8542 19168
rect 10778 19116 10784 19168
rect 10836 19156 10842 19168
rect 11057 19159 11115 19165
rect 11057 19156 11069 19159
rect 10836 19128 11069 19156
rect 10836 19116 10842 19128
rect 11057 19125 11069 19128
rect 11103 19125 11115 19159
rect 11164 19156 11192 19196
rect 11330 19184 11336 19236
rect 11388 19184 11394 19236
rect 11514 19184 11520 19236
rect 11572 19224 11578 19236
rect 11992 19224 12020 19320
rect 12342 19292 12348 19304
rect 11572 19196 12020 19224
rect 12084 19264 12348 19292
rect 11572 19184 11578 19196
rect 12084 19156 12112 19264
rect 12342 19252 12348 19264
rect 12400 19292 12406 19304
rect 13173 19295 13231 19301
rect 12400 19264 12848 19292
rect 12400 19252 12406 19264
rect 12820 19224 12848 19264
rect 13173 19261 13185 19295
rect 13219 19261 13231 19295
rect 13173 19255 13231 19261
rect 13188 19224 13216 19255
rect 12268 19196 12664 19224
rect 12820 19196 13216 19224
rect 11164 19128 12112 19156
rect 11057 19119 11115 19125
rect 12158 19116 12164 19168
rect 12216 19156 12222 19168
rect 12268 19165 12296 19196
rect 12253 19159 12311 19165
rect 12253 19156 12265 19159
rect 12216 19128 12265 19156
rect 12216 19116 12222 19128
rect 12253 19125 12265 19128
rect 12299 19125 12311 19159
rect 12253 19119 12311 19125
rect 12434 19116 12440 19168
rect 12492 19116 12498 19168
rect 12636 19156 12664 19196
rect 13740 19156 13768 19332
rect 13998 19320 14004 19332
rect 14056 19360 14062 19372
rect 15746 19360 15752 19372
rect 14056 19332 15752 19360
rect 14056 19320 14062 19332
rect 15746 19320 15752 19332
rect 15804 19360 15810 19372
rect 16390 19360 16396 19372
rect 15804 19332 16396 19360
rect 15804 19320 15810 19332
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 18874 19320 18880 19372
rect 18932 19320 18938 19372
rect 19242 19320 19248 19372
rect 19300 19320 19306 19372
rect 23474 19320 23480 19372
rect 23532 19320 23538 19372
rect 23750 19320 23756 19372
rect 23808 19320 23814 19372
rect 23952 19332 24532 19360
rect 14918 19252 14924 19304
rect 14976 19292 14982 19304
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14976 19264 15117 19292
rect 14976 19252 14982 19264
rect 15105 19261 15117 19264
rect 15151 19261 15163 19295
rect 15105 19255 15163 19261
rect 15289 19295 15347 19301
rect 15289 19261 15301 19295
rect 15335 19292 15347 19295
rect 15933 19295 15991 19301
rect 15933 19292 15945 19295
rect 15335 19264 15945 19292
rect 15335 19261 15347 19264
rect 15289 19255 15347 19261
rect 15933 19261 15945 19264
rect 15979 19292 15991 19295
rect 16482 19292 16488 19304
rect 15979 19264 16488 19292
rect 15979 19261 15991 19264
rect 15933 19255 15991 19261
rect 16482 19252 16488 19264
rect 16540 19252 16546 19304
rect 17126 19252 17132 19304
rect 17184 19252 17190 19304
rect 18969 19295 19027 19301
rect 18969 19261 18981 19295
rect 19015 19261 19027 19295
rect 20378 19264 21036 19292
rect 18969 19255 19027 19261
rect 18984 19224 19012 19255
rect 21008 19233 21036 19264
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 21140 19264 22017 19292
rect 21140 19252 21146 19264
rect 22005 19261 22017 19264
rect 22051 19261 22063 19295
rect 23492 19292 23520 19320
rect 23845 19295 23903 19301
rect 23845 19292 23857 19295
rect 23492 19264 23857 19292
rect 22005 19255 22063 19261
rect 23845 19261 23857 19264
rect 23891 19261 23903 19295
rect 23845 19255 23903 19261
rect 20993 19227 21051 19233
rect 18984 19196 19656 19224
rect 12636 19128 13768 19156
rect 14550 19116 14556 19168
rect 14608 19116 14614 19168
rect 15381 19159 15439 19165
rect 15381 19125 15393 19159
rect 15427 19156 15439 19159
rect 15562 19156 15568 19168
rect 15427 19128 15568 19156
rect 15427 19125 15439 19128
rect 15381 19119 15439 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 19628 19156 19656 19196
rect 20993 19193 21005 19227
rect 21039 19193 21051 19227
rect 20993 19187 21051 19193
rect 23658 19184 23664 19236
rect 23716 19224 23722 19236
rect 23952 19233 23980 19332
rect 24397 19295 24455 19301
rect 24397 19292 24409 19295
rect 24320 19264 24409 19292
rect 23937 19227 23995 19233
rect 23937 19224 23949 19227
rect 23716 19196 23949 19224
rect 23716 19184 23722 19196
rect 23937 19193 23949 19196
rect 23983 19193 23995 19227
rect 23937 19187 23995 19193
rect 20254 19156 20260 19168
rect 19628 19128 20260 19156
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 20714 19116 20720 19168
rect 20772 19116 20778 19168
rect 24320 19165 24348 19264
rect 24397 19261 24409 19264
rect 24443 19261 24455 19295
rect 24504 19292 24532 19332
rect 27080 19332 27292 19360
rect 25225 19295 25283 19301
rect 25225 19292 25237 19295
rect 24504 19264 25237 19292
rect 24397 19255 24455 19261
rect 25225 19261 25237 19264
rect 25271 19261 25283 19295
rect 25225 19255 25283 19261
rect 25314 19252 25320 19304
rect 25372 19252 25378 19304
rect 26697 19295 26755 19301
rect 26697 19261 26709 19295
rect 26743 19292 26755 19295
rect 26789 19295 26847 19301
rect 26789 19292 26801 19295
rect 26743 19264 26801 19292
rect 26743 19261 26755 19264
rect 26697 19255 26755 19261
rect 26789 19261 26801 19264
rect 26835 19261 26847 19295
rect 26789 19255 26847 19261
rect 26973 19295 27031 19301
rect 26973 19261 26985 19295
rect 27019 19292 27031 19295
rect 27080 19292 27108 19332
rect 27019 19264 27108 19292
rect 27019 19261 27031 19264
rect 26973 19255 27031 19261
rect 27154 19252 27160 19304
rect 27212 19252 27218 19304
rect 27264 19292 27292 19332
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 27433 19363 27491 19369
rect 27433 19360 27445 19363
rect 27396 19332 27445 19360
rect 27396 19320 27402 19332
rect 27433 19329 27445 19332
rect 27479 19360 27491 19363
rect 27890 19360 27896 19372
rect 27479 19332 27896 19360
rect 27479 19329 27491 19332
rect 27433 19323 27491 19329
rect 27890 19320 27896 19332
rect 27948 19320 27954 19372
rect 28184 19332 30144 19360
rect 28184 19292 28212 19332
rect 27264 19264 28212 19292
rect 28258 19252 28264 19304
rect 28316 19252 28322 19304
rect 30116 19301 30144 19332
rect 33778 19320 33784 19372
rect 33836 19320 33842 19372
rect 30101 19295 30159 19301
rect 30101 19261 30113 19295
rect 30147 19261 30159 19295
rect 30101 19255 30159 19261
rect 30650 19252 30656 19304
rect 30708 19292 30714 19304
rect 31294 19292 31300 19304
rect 30708 19264 31300 19292
rect 30708 19252 30714 19264
rect 31294 19252 31300 19264
rect 31352 19292 31358 19304
rect 31757 19295 31815 19301
rect 31757 19292 31769 19295
rect 31352 19264 31769 19292
rect 31352 19252 31358 19264
rect 31757 19261 31769 19264
rect 31803 19261 31815 19295
rect 31757 19255 31815 19261
rect 32766 19252 32772 19304
rect 32824 19252 32830 19304
rect 27065 19227 27123 19233
rect 27065 19193 27077 19227
rect 27111 19193 27123 19227
rect 27065 19187 27123 19193
rect 24305 19159 24363 19165
rect 24305 19125 24317 19159
rect 24351 19125 24363 19159
rect 24305 19119 24363 19125
rect 26050 19116 26056 19168
rect 26108 19116 26114 19168
rect 27080 19156 27108 19187
rect 27246 19184 27252 19236
rect 27304 19233 27310 19236
rect 27304 19227 27333 19233
rect 27321 19193 27333 19227
rect 29733 19227 29791 19233
rect 27304 19187 27333 19193
rect 27724 19196 28120 19224
rect 27304 19184 27310 19187
rect 27724 19168 27752 19196
rect 27430 19156 27436 19168
rect 27080 19128 27436 19156
rect 27430 19116 27436 19128
rect 27488 19116 27494 19168
rect 27706 19116 27712 19168
rect 27764 19116 27770 19168
rect 27798 19116 27804 19168
rect 27856 19116 27862 19168
rect 27890 19116 27896 19168
rect 27948 19116 27954 19168
rect 28092 19156 28120 19196
rect 29733 19193 29745 19227
rect 29779 19224 29791 19227
rect 29822 19224 29828 19236
rect 29779 19196 29828 19224
rect 29779 19193 29791 19196
rect 29733 19187 29791 19193
rect 29822 19184 29828 19196
rect 29880 19184 29886 19236
rect 29917 19227 29975 19233
rect 29917 19193 29929 19227
rect 29963 19193 29975 19227
rect 29917 19187 29975 19193
rect 29086 19156 29092 19168
rect 28092 19128 29092 19156
rect 29086 19116 29092 19128
rect 29144 19116 29150 19168
rect 29270 19116 29276 19168
rect 29328 19116 29334 19168
rect 29362 19116 29368 19168
rect 29420 19116 29426 19168
rect 29457 19159 29515 19165
rect 29457 19125 29469 19159
rect 29503 19156 29515 19159
rect 29546 19156 29552 19168
rect 29503 19128 29552 19156
rect 29503 19125 29515 19128
rect 29457 19119 29515 19125
rect 29546 19116 29552 19128
rect 29604 19116 29610 19168
rect 29932 19156 29960 19187
rect 30006 19156 30012 19168
rect 29932 19128 30012 19156
rect 30006 19116 30012 19128
rect 30064 19116 30070 19168
rect 30282 19116 30288 19168
rect 30340 19156 30346 19168
rect 31205 19159 31263 19165
rect 31205 19156 31217 19159
rect 30340 19128 31217 19156
rect 30340 19116 30346 19128
rect 31205 19125 31217 19128
rect 31251 19125 31263 19159
rect 31205 19119 31263 19125
rect 32490 19116 32496 19168
rect 32548 19156 32554 19168
rect 33042 19156 33048 19168
rect 32548 19128 33048 19156
rect 32548 19116 32554 19128
rect 33042 19116 33048 19128
rect 33100 19156 33106 19168
rect 33686 19156 33692 19168
rect 33100 19128 33692 19156
rect 33100 19116 33106 19128
rect 33686 19116 33692 19128
rect 33744 19116 33750 19168
rect 2760 19066 34316 19088
rect 2760 19014 7210 19066
rect 7262 19014 7274 19066
rect 7326 19014 7338 19066
rect 7390 19014 7402 19066
rect 7454 19014 7466 19066
rect 7518 19014 15099 19066
rect 15151 19014 15163 19066
rect 15215 19014 15227 19066
rect 15279 19014 15291 19066
rect 15343 19014 15355 19066
rect 15407 19014 22988 19066
rect 23040 19014 23052 19066
rect 23104 19014 23116 19066
rect 23168 19014 23180 19066
rect 23232 19014 23244 19066
rect 23296 19014 30877 19066
rect 30929 19014 30941 19066
rect 30993 19014 31005 19066
rect 31057 19014 31069 19066
rect 31121 19014 31133 19066
rect 31185 19014 34316 19066
rect 2760 18992 34316 19014
rect 4157 18955 4215 18961
rect 4157 18921 4169 18955
rect 4203 18952 4215 18955
rect 4522 18952 4528 18964
rect 4203 18924 4528 18952
rect 4203 18921 4215 18924
rect 4157 18915 4215 18921
rect 4522 18912 4528 18924
rect 4580 18912 4586 18964
rect 5258 18912 5264 18964
rect 5316 18952 5322 18964
rect 6917 18955 6975 18961
rect 5316 18924 6592 18952
rect 5316 18912 5322 18924
rect 4798 18884 4804 18896
rect 4264 18856 4804 18884
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 3053 18819 3111 18825
rect 3053 18816 3065 18819
rect 1360 18788 3065 18816
rect 1360 18776 1366 18788
rect 3053 18785 3065 18788
rect 3099 18785 3111 18819
rect 3053 18779 3111 18785
rect 3605 18819 3663 18825
rect 3605 18785 3617 18819
rect 3651 18816 3663 18819
rect 3694 18816 3700 18828
rect 3651 18788 3700 18816
rect 3651 18785 3663 18788
rect 3605 18779 3663 18785
rect 3694 18776 3700 18788
rect 3752 18776 3758 18828
rect 4264 18825 4292 18856
rect 4798 18844 4804 18856
rect 4856 18844 4862 18896
rect 5534 18844 5540 18896
rect 5592 18844 5598 18896
rect 5810 18844 5816 18896
rect 5868 18884 5874 18896
rect 6362 18884 6368 18896
rect 5868 18856 6368 18884
rect 5868 18844 5874 18856
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 4249 18819 4307 18825
rect 4249 18785 4261 18819
rect 4295 18785 4307 18819
rect 6564 18816 6592 18924
rect 6917 18921 6929 18955
rect 6963 18952 6975 18955
rect 7006 18952 7012 18964
rect 6963 18924 7012 18952
rect 6963 18921 6975 18924
rect 6917 18915 6975 18921
rect 7006 18912 7012 18924
rect 7064 18912 7070 18964
rect 7377 18955 7435 18961
rect 7377 18921 7389 18955
rect 7423 18952 7435 18955
rect 7650 18952 7656 18964
rect 7423 18924 7656 18952
rect 7423 18921 7435 18924
rect 7377 18915 7435 18921
rect 7650 18912 7656 18924
rect 7708 18912 7714 18964
rect 7742 18912 7748 18964
rect 7800 18912 7806 18964
rect 8478 18912 8484 18964
rect 8536 18912 8542 18964
rect 8941 18955 8999 18961
rect 8941 18921 8953 18955
rect 8987 18952 8999 18955
rect 9122 18952 9128 18964
rect 8987 18924 9128 18952
rect 8987 18921 8999 18924
rect 8941 18915 8999 18921
rect 9122 18912 9128 18924
rect 9180 18912 9186 18964
rect 9490 18912 9496 18964
rect 9548 18952 9554 18964
rect 11882 18952 11888 18964
rect 9548 18924 11888 18952
rect 9548 18912 9554 18924
rect 11882 18912 11888 18924
rect 11940 18952 11946 18964
rect 12158 18952 12164 18964
rect 11940 18924 12164 18952
rect 11940 18912 11946 18924
rect 12158 18912 12164 18924
rect 12216 18912 12222 18964
rect 12250 18912 12256 18964
rect 12308 18912 12314 18964
rect 14826 18952 14832 18964
rect 14384 18924 14832 18952
rect 8496 18884 8524 18912
rect 8496 18856 9628 18884
rect 7009 18819 7067 18825
rect 7009 18816 7021 18819
rect 6564 18788 7021 18816
rect 4249 18779 4307 18785
rect 7009 18785 7021 18788
rect 7055 18785 7067 18819
rect 7009 18779 7067 18785
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18785 7711 18819
rect 7653 18779 7711 18785
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 4982 18748 4988 18760
rect 4571 18720 4988 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 5997 18751 6055 18757
rect 5997 18717 6009 18751
rect 6043 18748 6055 18751
rect 6089 18751 6147 18757
rect 6089 18748 6101 18751
rect 6043 18720 6101 18748
rect 6043 18717 6055 18720
rect 5997 18711 6055 18717
rect 6089 18717 6101 18720
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 3234 18572 3240 18624
rect 3292 18572 3298 18624
rect 6178 18572 6184 18624
rect 6236 18612 6242 18624
rect 6733 18615 6791 18621
rect 6733 18612 6745 18615
rect 6236 18584 6745 18612
rect 6236 18572 6242 18584
rect 6733 18581 6745 18584
rect 6779 18581 6791 18615
rect 7668 18612 7696 18779
rect 8570 18776 8576 18828
rect 8628 18816 8634 18828
rect 9600 18825 9628 18856
rect 9950 18844 9956 18896
rect 10008 18844 10014 18896
rect 10870 18844 10876 18896
rect 10928 18884 10934 18896
rect 11057 18887 11115 18893
rect 11057 18884 11069 18887
rect 10928 18856 11069 18884
rect 10928 18844 10934 18856
rect 11057 18853 11069 18856
rect 11103 18884 11115 18887
rect 11514 18884 11520 18896
rect 11103 18856 11520 18884
rect 11103 18853 11115 18856
rect 11057 18847 11115 18853
rect 11514 18844 11520 18856
rect 11572 18844 11578 18896
rect 14384 18884 14412 18924
rect 14826 18912 14832 18924
rect 14884 18952 14890 18964
rect 14884 18924 16436 18952
rect 14884 18912 14890 18924
rect 12406 18856 14228 18884
rect 9033 18819 9091 18825
rect 9033 18816 9045 18819
rect 8628 18788 9045 18816
rect 8628 18776 8634 18788
rect 9033 18785 9045 18788
rect 9079 18785 9091 18819
rect 9033 18779 9091 18785
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18785 9643 18819
rect 12406 18816 12434 18856
rect 9585 18779 9643 18785
rect 9692 18788 12434 18816
rect 8386 18708 8392 18760
rect 8444 18708 8450 18760
rect 8478 18708 8484 18760
rect 8536 18748 8542 18760
rect 9398 18748 9404 18760
rect 8536 18720 9404 18748
rect 8536 18708 8542 18720
rect 9398 18708 9404 18720
rect 9456 18708 9462 18760
rect 8662 18640 8668 18692
rect 8720 18680 8726 18692
rect 9692 18680 9720 18788
rect 12894 18776 12900 18828
rect 12952 18816 12958 18828
rect 13173 18819 13231 18825
rect 13173 18816 13185 18819
rect 12952 18788 13185 18816
rect 12952 18776 12958 18788
rect 13173 18785 13185 18788
rect 13219 18785 13231 18819
rect 13906 18816 13912 18828
rect 13173 18779 13231 18785
rect 13464 18788 13912 18816
rect 11241 18751 11299 18757
rect 11241 18717 11253 18751
rect 11287 18717 11299 18751
rect 11241 18711 11299 18717
rect 12345 18751 12403 18757
rect 12345 18717 12357 18751
rect 12391 18717 12403 18751
rect 12345 18711 12403 18717
rect 8720 18652 9720 18680
rect 10781 18683 10839 18689
rect 8720 18640 8726 18652
rect 10781 18649 10793 18683
rect 10827 18649 10839 18683
rect 11256 18680 11284 18711
rect 11885 18683 11943 18689
rect 11885 18680 11897 18683
rect 11256 18652 11897 18680
rect 10781 18643 10839 18649
rect 11885 18649 11897 18652
rect 11931 18649 11943 18683
rect 12360 18680 12388 18711
rect 12434 18708 12440 18760
rect 12492 18708 12498 18760
rect 13464 18757 13492 18788
rect 13906 18776 13912 18788
rect 13964 18776 13970 18828
rect 13449 18751 13507 18757
rect 13449 18717 13461 18751
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 13998 18680 14004 18692
rect 12360 18652 14004 18680
rect 11885 18643 11943 18649
rect 9674 18612 9680 18624
rect 7668 18584 9680 18612
rect 6733 18575 6791 18581
rect 9674 18572 9680 18584
rect 9732 18572 9738 18624
rect 10594 18572 10600 18624
rect 10652 18572 10658 18624
rect 10796 18612 10824 18643
rect 13998 18640 14004 18652
rect 14056 18640 14062 18692
rect 11422 18612 11428 18624
rect 10796 18584 11428 18612
rect 11422 18572 11428 18584
rect 11480 18572 11486 18624
rect 11790 18572 11796 18624
rect 11848 18572 11854 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 12894 18612 12900 18624
rect 12216 18584 12900 18612
rect 12216 18572 12222 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 13814 18572 13820 18624
rect 13872 18572 13878 18624
rect 14200 18612 14228 18856
rect 14292 18856 14412 18884
rect 14292 18825 14320 18856
rect 15562 18844 15568 18896
rect 15620 18844 15626 18896
rect 14277 18819 14335 18825
rect 14277 18785 14289 18819
rect 14323 18785 14335 18819
rect 14277 18779 14335 18785
rect 16114 18776 16120 18828
rect 16172 18776 16178 18828
rect 14550 18708 14556 18760
rect 14608 18708 14614 18760
rect 16132 18680 16160 18776
rect 16408 18760 16436 18924
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17552 18924 19380 18952
rect 17552 18912 17558 18924
rect 17402 18844 17408 18896
rect 17460 18844 17466 18896
rect 19352 18884 19380 18924
rect 19426 18912 19432 18964
rect 19484 18912 19490 18964
rect 19518 18912 19524 18964
rect 19576 18912 19582 18964
rect 19613 18955 19671 18961
rect 19613 18921 19625 18955
rect 19659 18952 19671 18955
rect 19794 18952 19800 18964
rect 19659 18924 19800 18952
rect 19659 18921 19671 18924
rect 19613 18915 19671 18921
rect 19794 18912 19800 18924
rect 19852 18952 19858 18964
rect 19852 18924 20208 18952
rect 19852 18912 19858 18924
rect 19536 18884 19564 18912
rect 19352 18856 19564 18884
rect 18506 18776 18512 18828
rect 18564 18816 18570 18828
rect 19061 18819 19119 18825
rect 19061 18816 19073 18819
rect 18564 18788 19073 18816
rect 18564 18776 18570 18788
rect 19061 18785 19073 18788
rect 19107 18816 19119 18819
rect 19150 18816 19156 18828
rect 19107 18788 19156 18816
rect 19107 18785 19119 18788
rect 19061 18779 19119 18785
rect 19150 18776 19156 18788
rect 19208 18816 19214 18828
rect 19208 18788 19656 18816
rect 19208 18776 19214 18788
rect 16390 18708 16396 18760
rect 16448 18708 16454 18760
rect 16666 18708 16672 18760
rect 16724 18708 16730 18760
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18748 18199 18751
rect 18877 18751 18935 18757
rect 18877 18748 18889 18751
rect 18187 18720 18889 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 18877 18717 18889 18720
rect 18923 18717 18935 18751
rect 18877 18711 18935 18717
rect 15580 18652 16160 18680
rect 19628 18680 19656 18788
rect 19794 18776 19800 18828
rect 19852 18776 19858 18828
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18785 19947 18819
rect 19889 18779 19947 18785
rect 19904 18748 19932 18779
rect 20180 18748 20208 18924
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 26050 18952 26056 18964
rect 20772 18924 23244 18952
rect 20772 18912 20778 18924
rect 23216 18884 23244 18924
rect 24596 18924 26056 18952
rect 24596 18893 24624 18924
rect 26050 18912 26056 18924
rect 26108 18912 26114 18964
rect 27982 18912 27988 18964
rect 28040 18952 28046 18964
rect 28077 18955 28135 18961
rect 28077 18952 28089 18955
rect 28040 18924 28089 18952
rect 28040 18912 28046 18924
rect 28077 18921 28089 18924
rect 28123 18952 28135 18955
rect 28902 18952 28908 18964
rect 28123 18924 28908 18952
rect 28123 18921 28135 18924
rect 28077 18915 28135 18921
rect 28902 18912 28908 18924
rect 28960 18912 28966 18964
rect 29365 18955 29423 18961
rect 29365 18921 29377 18955
rect 29411 18952 29423 18955
rect 29454 18952 29460 18964
rect 29411 18924 29460 18952
rect 29411 18921 29423 18924
rect 29365 18915 29423 18921
rect 29454 18912 29460 18924
rect 29512 18912 29518 18964
rect 29546 18912 29552 18964
rect 29604 18952 29610 18964
rect 30193 18955 30251 18961
rect 30193 18952 30205 18955
rect 29604 18924 30205 18952
rect 29604 18912 29610 18924
rect 30193 18921 30205 18924
rect 30239 18921 30251 18955
rect 30193 18915 30251 18921
rect 30285 18955 30343 18961
rect 30285 18921 30297 18955
rect 30331 18921 30343 18955
rect 30285 18915 30343 18921
rect 31849 18955 31907 18961
rect 31849 18921 31861 18955
rect 31895 18952 31907 18955
rect 32490 18952 32496 18964
rect 31895 18924 32496 18952
rect 31895 18921 31907 18924
rect 31849 18915 31907 18921
rect 24581 18887 24639 18893
rect 23216 18856 23612 18884
rect 20346 18776 20352 18828
rect 20404 18816 20410 18828
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 20404 18788 21189 18816
rect 20404 18776 20410 18788
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 19904 18720 20208 18748
rect 20990 18708 20996 18760
rect 21048 18708 21054 18760
rect 23474 18708 23480 18760
rect 23532 18708 23538 18760
rect 23584 18748 23612 18856
rect 24581 18853 24593 18887
rect 24627 18853 24639 18887
rect 27706 18884 27712 18896
rect 24581 18847 24639 18853
rect 26252 18856 27712 18884
rect 24118 18776 24124 18828
rect 24176 18816 24182 18828
rect 24305 18819 24363 18825
rect 24305 18816 24317 18819
rect 24176 18788 24317 18816
rect 24176 18776 24182 18788
rect 24305 18785 24317 18788
rect 24351 18785 24363 18819
rect 24305 18779 24363 18785
rect 25682 18776 25688 18828
rect 25740 18776 25746 18828
rect 26252 18825 26280 18856
rect 27706 18844 27712 18856
rect 27764 18844 27770 18896
rect 28442 18844 28448 18896
rect 28500 18884 28506 18896
rect 28810 18884 28816 18896
rect 28500 18856 28816 18884
rect 28500 18844 28506 18856
rect 28810 18844 28816 18856
rect 28868 18884 28874 18896
rect 28868 18856 29592 18884
rect 28868 18844 28874 18856
rect 26237 18819 26295 18825
rect 26237 18785 26249 18819
rect 26283 18785 26295 18819
rect 26237 18779 26295 18785
rect 26421 18819 26479 18825
rect 26421 18785 26433 18819
rect 26467 18816 26479 18819
rect 26789 18819 26847 18825
rect 26789 18816 26801 18819
rect 26467 18788 26801 18816
rect 26467 18785 26479 18788
rect 26421 18779 26479 18785
rect 26789 18785 26801 18788
rect 26835 18816 26847 18819
rect 27338 18816 27344 18828
rect 26835 18788 27344 18816
rect 26835 18785 26847 18788
rect 26789 18779 26847 18785
rect 27338 18776 27344 18788
rect 27396 18776 27402 18828
rect 27433 18819 27491 18825
rect 27433 18785 27445 18819
rect 27479 18785 27491 18819
rect 27433 18779 27491 18785
rect 26053 18751 26111 18757
rect 23584 18720 25636 18748
rect 20349 18683 20407 18689
rect 20349 18680 20361 18683
rect 19628 18652 20361 18680
rect 15580 18612 15608 18652
rect 20349 18649 20361 18652
rect 20395 18649 20407 18683
rect 23934 18680 23940 18692
rect 20349 18643 20407 18649
rect 21284 18652 23940 18680
rect 14200 18584 15608 18612
rect 16025 18615 16083 18621
rect 16025 18581 16037 18615
rect 16071 18612 16083 18615
rect 16758 18612 16764 18624
rect 16071 18584 16764 18612
rect 16071 18581 16083 18584
rect 16025 18575 16083 18581
rect 16758 18572 16764 18584
rect 16816 18572 16822 18624
rect 17770 18572 17776 18624
rect 17828 18612 17834 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 17828 18584 18337 18612
rect 17828 18572 17834 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 18325 18575 18383 18581
rect 19429 18615 19487 18621
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 19518 18612 19524 18624
rect 19475 18584 19524 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 20073 18615 20131 18621
rect 20073 18581 20085 18615
rect 20119 18612 20131 18615
rect 21284 18612 21312 18652
rect 23934 18640 23940 18652
rect 23992 18640 23998 18692
rect 25608 18680 25636 18720
rect 26053 18717 26065 18751
rect 26099 18748 26111 18751
rect 26513 18751 26571 18757
rect 26513 18748 26525 18751
rect 26099 18720 26525 18748
rect 26099 18717 26111 18720
rect 26053 18711 26111 18717
rect 26513 18717 26525 18720
rect 26559 18717 26571 18751
rect 26513 18711 26571 18717
rect 27448 18680 27476 18779
rect 28994 18776 29000 18828
rect 29052 18816 29058 18828
rect 29564 18825 29592 18856
rect 29638 18844 29644 18896
rect 29696 18884 29702 18896
rect 30300 18884 30328 18915
rect 32490 18912 32496 18924
rect 32548 18912 32554 18964
rect 30650 18884 30656 18896
rect 29696 18856 30656 18884
rect 29696 18844 29702 18856
rect 30650 18844 30656 18856
rect 30708 18844 30714 18896
rect 29181 18819 29239 18825
rect 29181 18816 29193 18819
rect 29052 18788 29193 18816
rect 29052 18776 29058 18788
rect 29181 18785 29193 18788
rect 29227 18785 29239 18819
rect 29181 18779 29239 18785
rect 29549 18819 29607 18825
rect 29549 18785 29561 18819
rect 29595 18785 29607 18819
rect 29549 18779 29607 18785
rect 30006 18776 30012 18828
rect 30064 18776 30070 18828
rect 30098 18776 30104 18828
rect 30156 18776 30162 18828
rect 30282 18776 30288 18828
rect 30340 18816 30346 18828
rect 30561 18819 30619 18825
rect 30561 18816 30573 18819
rect 30340 18788 30573 18816
rect 30340 18776 30346 18788
rect 30561 18785 30573 18788
rect 30607 18785 30619 18819
rect 30561 18779 30619 18785
rect 31941 18819 31999 18825
rect 31941 18785 31953 18819
rect 31987 18816 31999 18819
rect 32950 18816 32956 18828
rect 31987 18788 32956 18816
rect 31987 18785 31999 18788
rect 31941 18779 31999 18785
rect 32950 18776 32956 18788
rect 33008 18776 33014 18828
rect 33502 18776 33508 18828
rect 33560 18776 33566 18828
rect 29638 18708 29644 18760
rect 29696 18708 29702 18760
rect 30024 18748 30052 18776
rect 29748 18720 30052 18748
rect 25608 18652 27476 18680
rect 27890 18640 27896 18692
rect 27948 18680 27954 18692
rect 29748 18680 29776 18720
rect 27948 18652 29776 18680
rect 27948 18640 27954 18652
rect 29822 18640 29828 18692
rect 29880 18680 29886 18692
rect 30300 18680 30328 18776
rect 30469 18751 30527 18757
rect 30469 18717 30481 18751
rect 30515 18717 30527 18751
rect 30469 18711 30527 18717
rect 30745 18751 30803 18757
rect 30745 18717 30757 18751
rect 30791 18748 30803 18751
rect 31389 18751 31447 18757
rect 31389 18748 31401 18751
rect 30791 18720 31401 18748
rect 30791 18717 30803 18720
rect 30745 18711 30803 18717
rect 31389 18717 31401 18720
rect 31435 18717 31447 18751
rect 31389 18711 31447 18717
rect 33045 18751 33103 18757
rect 33045 18717 33057 18751
rect 33091 18748 33103 18751
rect 34514 18748 34520 18760
rect 33091 18720 34520 18748
rect 33091 18717 33103 18720
rect 33045 18711 33103 18717
rect 29880 18652 30328 18680
rect 29880 18640 29886 18652
rect 20119 18584 21312 18612
rect 20119 18581 20131 18584
rect 20073 18575 20131 18581
rect 21358 18572 21364 18624
rect 21416 18572 21422 18624
rect 21634 18572 21640 18624
rect 21692 18612 21698 18624
rect 23201 18615 23259 18621
rect 23201 18612 23213 18615
rect 21692 18584 23213 18612
rect 21692 18572 21698 18584
rect 23201 18581 23213 18584
rect 23247 18612 23259 18615
rect 23382 18612 23388 18624
rect 23247 18584 23388 18612
rect 23247 18581 23259 18584
rect 23201 18575 23259 18581
rect 23382 18572 23388 18584
rect 23440 18572 23446 18624
rect 24121 18615 24179 18621
rect 24121 18581 24133 18615
rect 24167 18612 24179 18615
rect 24394 18612 24400 18624
rect 24167 18584 24400 18612
rect 24167 18581 24179 18584
rect 24121 18575 24179 18581
rect 24394 18572 24400 18584
rect 24452 18572 24458 18624
rect 26329 18615 26387 18621
rect 26329 18581 26341 18615
rect 26375 18612 26387 18615
rect 27430 18612 27436 18624
rect 26375 18584 27436 18612
rect 26375 18581 26387 18584
rect 26329 18575 26387 18581
rect 27430 18572 27436 18584
rect 27488 18572 27494 18624
rect 28166 18572 28172 18624
rect 28224 18612 28230 18624
rect 28629 18615 28687 18621
rect 28629 18612 28641 18615
rect 28224 18584 28641 18612
rect 28224 18572 28230 18584
rect 28629 18581 28641 18584
rect 28675 18581 28687 18615
rect 28629 18575 28687 18581
rect 28810 18572 28816 18624
rect 28868 18612 28874 18624
rect 29549 18615 29607 18621
rect 29549 18612 29561 18615
rect 28868 18584 29561 18612
rect 28868 18572 28874 18584
rect 29549 18581 29561 18584
rect 29595 18581 29607 18615
rect 29549 18575 29607 18581
rect 29914 18572 29920 18624
rect 29972 18612 29978 18624
rect 30484 18612 30512 18711
rect 34514 18708 34520 18720
rect 34572 18708 34578 18760
rect 29972 18584 30512 18612
rect 29972 18572 29978 18584
rect 30834 18572 30840 18624
rect 30892 18572 30898 18624
rect 32030 18572 32036 18624
rect 32088 18572 32094 18624
rect 2760 18522 34316 18544
rect 2760 18470 6550 18522
rect 6602 18470 6614 18522
rect 6666 18470 6678 18522
rect 6730 18470 6742 18522
rect 6794 18470 6806 18522
rect 6858 18470 14439 18522
rect 14491 18470 14503 18522
rect 14555 18470 14567 18522
rect 14619 18470 14631 18522
rect 14683 18470 14695 18522
rect 14747 18470 22328 18522
rect 22380 18470 22392 18522
rect 22444 18470 22456 18522
rect 22508 18470 22520 18522
rect 22572 18470 22584 18522
rect 22636 18470 30217 18522
rect 30269 18470 30281 18522
rect 30333 18470 30345 18522
rect 30397 18470 30409 18522
rect 30461 18470 30473 18522
rect 30525 18470 34316 18522
rect 2760 18448 34316 18470
rect 3234 18368 3240 18420
rect 3292 18368 3298 18420
rect 3602 18368 3608 18420
rect 3660 18408 3666 18420
rect 6546 18408 6552 18420
rect 3660 18380 6552 18408
rect 3660 18368 3666 18380
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 8570 18368 8576 18420
rect 8628 18368 8634 18420
rect 11790 18368 11796 18420
rect 11848 18408 11854 18420
rect 12050 18411 12108 18417
rect 12050 18408 12062 18411
rect 11848 18380 12062 18408
rect 11848 18368 11854 18380
rect 12050 18377 12062 18380
rect 12096 18377 12108 18411
rect 12050 18371 12108 18377
rect 13814 18368 13820 18420
rect 13872 18368 13878 18420
rect 13998 18368 14004 18420
rect 14056 18408 14062 18420
rect 14461 18411 14519 18417
rect 14461 18408 14473 18411
rect 14056 18380 14473 18408
rect 14056 18368 14062 18380
rect 14461 18377 14473 18380
rect 14507 18377 14519 18411
rect 14461 18371 14519 18377
rect 14553 18411 14611 18417
rect 14553 18377 14565 18411
rect 14599 18408 14611 18411
rect 14918 18408 14924 18420
rect 14599 18380 14924 18408
rect 14599 18377 14611 18380
rect 14553 18371 14611 18377
rect 3252 18340 3280 18368
rect 3252 18312 6316 18340
rect 5261 18275 5319 18281
rect 5261 18241 5273 18275
rect 5307 18272 5319 18275
rect 5718 18272 5724 18284
rect 5307 18244 5724 18272
rect 5307 18241 5319 18244
rect 5261 18235 5319 18241
rect 5718 18232 5724 18244
rect 5776 18232 5782 18284
rect 5810 18232 5816 18284
rect 5868 18272 5874 18284
rect 6181 18275 6239 18281
rect 6181 18272 6193 18275
rect 5868 18244 6193 18272
rect 5868 18232 5874 18244
rect 6181 18241 6193 18244
rect 6227 18241 6239 18275
rect 6288 18272 6316 18312
rect 6457 18275 6515 18281
rect 6457 18272 6469 18275
rect 6288 18244 6469 18272
rect 6181 18235 6239 18241
rect 6457 18241 6469 18244
rect 6503 18241 6515 18275
rect 6457 18235 6515 18241
rect 6546 18232 6552 18284
rect 6604 18281 6610 18284
rect 8588 18281 8616 18368
rect 9033 18343 9091 18349
rect 9033 18309 9045 18343
rect 9079 18340 9091 18343
rect 9953 18343 10011 18349
rect 9079 18312 9720 18340
rect 9079 18309 9091 18312
rect 9033 18303 9091 18309
rect 6604 18275 6632 18281
rect 6620 18241 6632 18275
rect 6604 18235 6632 18241
rect 6733 18275 6791 18281
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 8481 18275 8539 18281
rect 6779 18244 7696 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 6604 18232 6610 18235
rect 7668 18216 7696 18244
rect 8481 18241 8493 18275
rect 8527 18241 8539 18275
rect 8481 18235 8539 18241
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18241 8631 18275
rect 8573 18235 8631 18241
rect 3329 18207 3387 18213
rect 3329 18173 3341 18207
rect 3375 18204 3387 18207
rect 3789 18207 3847 18213
rect 3789 18204 3801 18207
rect 3375 18176 3801 18204
rect 3375 18173 3387 18176
rect 3329 18167 3387 18173
rect 3789 18173 3801 18176
rect 3835 18173 3847 18207
rect 3789 18167 3847 18173
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 4706 18204 4712 18216
rect 4663 18176 4712 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 3804 18136 3832 18167
rect 4706 18164 4712 18176
rect 4764 18204 4770 18216
rect 5074 18204 5080 18216
rect 4764 18176 5080 18204
rect 4764 18164 4770 18176
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5537 18207 5595 18213
rect 5537 18173 5549 18207
rect 5583 18173 5595 18207
rect 5537 18167 5595 18173
rect 5258 18136 5264 18148
rect 3804 18108 5264 18136
rect 5258 18096 5264 18108
rect 5316 18096 5322 18148
rect 3418 18028 3424 18080
rect 3476 18028 3482 18080
rect 5552 18068 5580 18167
rect 7650 18164 7656 18216
rect 7708 18164 7714 18216
rect 8496 18204 8524 18235
rect 8846 18232 8852 18284
rect 8904 18232 8910 18284
rect 9692 18281 9720 18312
rect 9953 18309 9965 18343
rect 9999 18340 10011 18343
rect 13832 18340 13860 18368
rect 9999 18312 11468 18340
rect 9999 18309 10011 18312
rect 9953 18303 10011 18309
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 10594 18272 10600 18284
rect 9677 18235 9735 18241
rect 10152 18244 10600 18272
rect 8864 18204 8892 18232
rect 10152 18213 10180 18244
rect 10594 18232 10600 18244
rect 10652 18232 10658 18284
rect 10778 18232 10784 18284
rect 10836 18232 10842 18284
rect 11440 18281 11468 18312
rect 13188 18312 13860 18340
rect 11425 18275 11483 18281
rect 11425 18241 11437 18275
rect 11471 18241 11483 18275
rect 11425 18235 11483 18241
rect 11793 18275 11851 18281
rect 11793 18241 11805 18275
rect 11839 18272 11851 18275
rect 13078 18272 13084 18284
rect 11839 18244 13084 18272
rect 11839 18241 11851 18244
rect 11793 18235 11851 18241
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 8496 18176 8892 18204
rect 10137 18207 10195 18213
rect 10137 18173 10149 18207
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10413 18207 10471 18213
rect 10413 18173 10425 18207
rect 10459 18204 10471 18207
rect 10796 18204 10824 18232
rect 10459 18176 10824 18204
rect 13188 18190 13216 18312
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18272 13599 18275
rect 13817 18275 13875 18281
rect 13817 18272 13829 18275
rect 13587 18244 13829 18272
rect 13587 18241 13599 18244
rect 13541 18235 13599 18241
rect 13817 18241 13829 18244
rect 13863 18241 13875 18275
rect 14476 18272 14504 18371
rect 14918 18368 14924 18380
rect 14976 18368 14982 18420
rect 16666 18368 16672 18420
rect 16724 18408 16730 18420
rect 16761 18411 16819 18417
rect 16761 18408 16773 18411
rect 16724 18380 16773 18408
rect 16724 18368 16730 18380
rect 16761 18377 16773 18380
rect 16807 18377 16819 18411
rect 16761 18371 16819 18377
rect 16960 18380 18368 18408
rect 16960 18340 16988 18380
rect 17589 18343 17647 18349
rect 17589 18340 17601 18343
rect 16224 18312 16988 18340
rect 17052 18312 17601 18340
rect 15013 18275 15071 18281
rect 15013 18272 15025 18275
rect 14476 18244 15025 18272
rect 13817 18235 13875 18241
rect 15013 18241 15025 18244
rect 15059 18241 15071 18275
rect 15013 18235 15071 18241
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18241 15163 18275
rect 15105 18235 15163 18241
rect 15120 18204 15148 18235
rect 13832 18176 15148 18204
rect 10459 18173 10471 18176
rect 10413 18167 10471 18173
rect 13832 18148 13860 18176
rect 7837 18139 7895 18145
rect 7837 18136 7849 18139
rect 7300 18108 7849 18136
rect 5994 18068 6000 18080
rect 5552 18040 6000 18068
rect 5994 18028 6000 18040
rect 6052 18028 6058 18080
rect 6362 18028 6368 18080
rect 6420 18068 6426 18080
rect 7300 18068 7328 18108
rect 7837 18105 7849 18108
rect 7883 18136 7895 18139
rect 8018 18136 8024 18148
rect 7883 18108 8024 18136
rect 7883 18105 7895 18108
rect 7837 18099 7895 18105
rect 8018 18096 8024 18108
rect 8076 18096 8082 18148
rect 8665 18139 8723 18145
rect 8665 18105 8677 18139
rect 8711 18136 8723 18139
rect 8711 18108 9812 18136
rect 8711 18105 8723 18108
rect 8665 18099 8723 18105
rect 9784 18080 9812 18108
rect 10336 18108 11376 18136
rect 6420 18040 7328 18068
rect 7377 18071 7435 18077
rect 6420 18028 6426 18040
rect 7377 18037 7389 18071
rect 7423 18068 7435 18071
rect 7742 18068 7748 18080
rect 7423 18040 7748 18068
rect 7423 18037 7435 18040
rect 7377 18031 7435 18037
rect 7742 18028 7748 18040
rect 7800 18028 7806 18080
rect 9122 18028 9128 18080
rect 9180 18028 9186 18080
rect 9766 18028 9772 18080
rect 9824 18028 9830 18080
rect 10336 18077 10364 18108
rect 10321 18071 10379 18077
rect 10321 18037 10333 18071
rect 10367 18037 10379 18071
rect 10321 18031 10379 18037
rect 10870 18028 10876 18080
rect 10928 18028 10934 18080
rect 11348 18068 11376 18108
rect 13814 18096 13820 18148
rect 13872 18096 13878 18148
rect 14921 18139 14979 18145
rect 14921 18105 14933 18139
rect 14967 18136 14979 18139
rect 15749 18139 15807 18145
rect 15749 18136 15761 18139
rect 14967 18108 15761 18136
rect 14967 18105 14979 18108
rect 14921 18099 14979 18105
rect 15749 18105 15761 18108
rect 15795 18105 15807 18139
rect 15749 18099 15807 18105
rect 12894 18068 12900 18080
rect 11348 18040 12900 18068
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 12986 18028 12992 18080
rect 13044 18068 13050 18080
rect 16224 18068 16252 18312
rect 16298 18232 16304 18284
rect 16356 18272 16362 18284
rect 17052 18272 17080 18312
rect 17589 18309 17601 18312
rect 17635 18309 17647 18343
rect 17589 18303 17647 18309
rect 16356 18244 17080 18272
rect 16356 18232 16362 18244
rect 17310 18232 17316 18284
rect 17368 18232 17374 18284
rect 17770 18281 17776 18284
rect 17748 18275 17776 18281
rect 17748 18241 17760 18275
rect 17748 18235 17776 18241
rect 17763 18232 17776 18235
rect 17828 18232 17834 18284
rect 17862 18232 17868 18284
rect 17920 18232 17926 18284
rect 16393 18207 16451 18213
rect 16393 18173 16405 18207
rect 16439 18204 16451 18207
rect 16758 18204 16764 18216
rect 16439 18176 16764 18204
rect 16439 18173 16451 18176
rect 16393 18167 16451 18173
rect 16758 18164 16764 18176
rect 16816 18204 16822 18216
rect 16942 18204 16948 18216
rect 16816 18176 16948 18204
rect 16816 18164 16822 18176
rect 16942 18164 16948 18176
rect 17000 18164 17006 18216
rect 17221 18207 17279 18213
rect 17221 18173 17233 18207
rect 17267 18204 17279 18207
rect 17763 18204 17791 18232
rect 17267 18176 17791 18204
rect 18233 18207 18291 18213
rect 17267 18173 17279 18176
rect 17221 18167 17279 18173
rect 18233 18173 18245 18207
rect 18279 18173 18291 18207
rect 18233 18167 18291 18173
rect 18248 18136 18276 18167
rect 17236 18108 18276 18136
rect 18340 18136 18368 18380
rect 19058 18368 19064 18420
rect 19116 18368 19122 18420
rect 23017 18411 23075 18417
rect 23017 18377 23029 18411
rect 23063 18408 23075 18411
rect 23474 18408 23480 18420
rect 23063 18380 23480 18408
rect 23063 18377 23075 18380
rect 23017 18371 23075 18377
rect 23474 18368 23480 18380
rect 23532 18368 23538 18420
rect 24044 18380 25636 18408
rect 18782 18300 18788 18352
rect 18840 18340 18846 18352
rect 19521 18343 19579 18349
rect 19521 18340 19533 18343
rect 18840 18312 19533 18340
rect 18840 18300 18846 18312
rect 19521 18309 19533 18312
rect 19567 18340 19579 18343
rect 19794 18340 19800 18352
rect 19567 18312 19800 18340
rect 19567 18309 19579 18312
rect 19521 18303 19579 18309
rect 19794 18300 19800 18312
rect 19852 18300 19858 18352
rect 18690 18232 18696 18284
rect 18748 18272 18754 18284
rect 19058 18272 19064 18284
rect 18748 18244 19064 18272
rect 18748 18232 18754 18244
rect 19058 18232 19064 18244
rect 19116 18232 19122 18284
rect 20254 18232 20260 18284
rect 20312 18272 20318 18284
rect 20806 18272 20812 18284
rect 20312 18244 20812 18272
rect 20312 18232 20318 18244
rect 20806 18232 20812 18244
rect 20864 18272 20870 18284
rect 21269 18275 21327 18281
rect 21269 18272 21281 18275
rect 20864 18244 21281 18272
rect 20864 18232 20870 18244
rect 21269 18241 21281 18244
rect 21315 18241 21327 18275
rect 21269 18235 21327 18241
rect 23566 18232 23572 18284
rect 23624 18232 23630 18284
rect 18506 18164 18512 18216
rect 18564 18164 18570 18216
rect 18598 18164 18604 18216
rect 18656 18164 18662 18216
rect 18782 18164 18788 18216
rect 18840 18164 18846 18216
rect 18966 18164 18972 18216
rect 19024 18164 19030 18216
rect 23293 18207 23351 18213
rect 23293 18173 23305 18207
rect 23339 18204 23351 18207
rect 24044 18204 24072 18380
rect 24121 18343 24179 18349
rect 24121 18309 24133 18343
rect 24167 18309 24179 18343
rect 24121 18303 24179 18309
rect 23339 18176 24072 18204
rect 24136 18204 24164 18303
rect 24394 18232 24400 18284
rect 24452 18272 24458 18284
rect 24765 18275 24823 18281
rect 24765 18272 24777 18275
rect 24452 18244 24777 18272
rect 24452 18232 24458 18244
rect 24765 18241 24777 18244
rect 24811 18241 24823 18275
rect 24765 18235 24823 18241
rect 25501 18207 25559 18213
rect 25501 18204 25513 18207
rect 24136 18176 25513 18204
rect 23339 18173 23351 18176
rect 23293 18167 23351 18173
rect 18984 18136 19012 18164
rect 23492 18148 23520 18176
rect 25501 18173 25513 18176
rect 25547 18173 25559 18207
rect 25608 18204 25636 18380
rect 25682 18368 25688 18420
rect 25740 18408 25746 18420
rect 25777 18411 25835 18417
rect 25777 18408 25789 18411
rect 25740 18380 25789 18408
rect 25740 18368 25746 18380
rect 25777 18377 25789 18380
rect 25823 18377 25835 18411
rect 25777 18371 25835 18377
rect 27798 18368 27804 18420
rect 27856 18408 27862 18420
rect 28350 18408 28356 18420
rect 27856 18380 28356 18408
rect 27856 18368 27862 18380
rect 28350 18368 28356 18380
rect 28408 18368 28414 18420
rect 28460 18380 28856 18408
rect 27522 18300 27528 18352
rect 27580 18340 27586 18352
rect 27985 18343 28043 18349
rect 27985 18340 27997 18343
rect 27580 18312 27997 18340
rect 27580 18300 27586 18312
rect 27985 18309 27997 18312
rect 28031 18309 28043 18343
rect 27985 18303 28043 18309
rect 28074 18300 28080 18352
rect 28132 18340 28138 18352
rect 28460 18340 28488 18380
rect 28132 18312 28488 18340
rect 28537 18343 28595 18349
rect 28132 18300 28138 18312
rect 28537 18309 28549 18343
rect 28583 18309 28595 18343
rect 28537 18303 28595 18309
rect 28552 18272 28580 18303
rect 26988 18244 28580 18272
rect 25685 18207 25743 18213
rect 25685 18204 25697 18207
rect 25608 18176 25697 18204
rect 25501 18167 25559 18173
rect 25685 18173 25697 18176
rect 25731 18173 25743 18207
rect 25685 18167 25743 18173
rect 26602 18164 26608 18216
rect 26660 18164 26666 18216
rect 26786 18164 26792 18216
rect 26844 18164 26850 18216
rect 26988 18213 27016 18244
rect 26973 18207 27031 18213
rect 26973 18173 26985 18207
rect 27019 18173 27031 18207
rect 26973 18167 27031 18173
rect 27157 18207 27215 18213
rect 27157 18173 27169 18207
rect 27203 18173 27215 18207
rect 27157 18167 27215 18173
rect 18340 18108 19012 18136
rect 17236 18080 17264 18108
rect 21542 18096 21548 18148
rect 21600 18096 21606 18148
rect 23201 18139 23259 18145
rect 23201 18136 23213 18139
rect 22770 18108 23213 18136
rect 23201 18105 23213 18108
rect 23247 18105 23259 18139
rect 23201 18099 23259 18105
rect 23474 18096 23480 18148
rect 23532 18096 23538 18148
rect 23753 18139 23811 18145
rect 23753 18105 23765 18139
rect 23799 18136 23811 18139
rect 26053 18139 26111 18145
rect 26053 18136 26065 18139
rect 23799 18108 26065 18136
rect 23799 18105 23811 18108
rect 23753 18099 23811 18105
rect 26053 18105 26065 18108
rect 26099 18105 26111 18139
rect 27172 18136 27200 18167
rect 27430 18164 27436 18216
rect 27488 18204 27494 18216
rect 28442 18213 28448 18216
rect 27893 18207 27951 18213
rect 27893 18204 27905 18207
rect 27488 18176 27905 18204
rect 27488 18164 27494 18176
rect 27893 18173 27905 18176
rect 27939 18173 27951 18207
rect 27893 18167 27951 18173
rect 28412 18207 28448 18213
rect 28412 18173 28424 18207
rect 28412 18167 28448 18173
rect 28442 18164 28448 18167
rect 28500 18164 28506 18216
rect 28828 18213 28856 18380
rect 29270 18368 29276 18420
rect 29328 18408 29334 18420
rect 29457 18411 29515 18417
rect 29457 18408 29469 18411
rect 29328 18380 29469 18408
rect 29328 18368 29334 18380
rect 29457 18377 29469 18380
rect 29503 18377 29515 18411
rect 29457 18371 29515 18377
rect 30653 18411 30711 18417
rect 30653 18377 30665 18411
rect 30699 18408 30711 18411
rect 30742 18408 30748 18420
rect 30699 18380 30748 18408
rect 30699 18377 30711 18380
rect 30653 18371 30711 18377
rect 30742 18368 30748 18380
rect 30800 18368 30806 18420
rect 29362 18300 29368 18352
rect 29420 18340 29426 18352
rect 29549 18343 29607 18349
rect 29549 18340 29561 18343
rect 29420 18312 29561 18340
rect 29420 18300 29426 18312
rect 29549 18309 29561 18312
rect 29595 18340 29607 18343
rect 29822 18340 29828 18352
rect 29595 18312 29828 18340
rect 29595 18309 29607 18312
rect 29549 18303 29607 18309
rect 29822 18300 29828 18312
rect 29880 18300 29886 18352
rect 30837 18343 30895 18349
rect 30837 18309 30849 18343
rect 30883 18340 30895 18343
rect 31202 18340 31208 18352
rect 30883 18312 31208 18340
rect 30883 18309 30895 18312
rect 30837 18303 30895 18309
rect 31202 18300 31208 18312
rect 31260 18300 31266 18352
rect 28902 18232 28908 18284
rect 28960 18272 28966 18284
rect 28960 18244 33456 18272
rect 28960 18232 28966 18244
rect 28813 18207 28871 18213
rect 28813 18173 28825 18207
rect 28859 18173 28871 18207
rect 28813 18167 28871 18173
rect 29089 18207 29147 18213
rect 29089 18173 29101 18207
rect 29135 18204 29147 18207
rect 29638 18204 29644 18216
rect 29135 18176 29644 18204
rect 29135 18173 29147 18176
rect 29089 18167 29147 18173
rect 29638 18164 29644 18176
rect 29696 18164 29702 18216
rect 29917 18207 29975 18213
rect 29917 18173 29929 18207
rect 29963 18204 29975 18207
rect 30098 18204 30104 18216
rect 29963 18176 30104 18204
rect 29963 18173 29975 18176
rect 29917 18167 29975 18173
rect 30098 18164 30104 18176
rect 30156 18164 30162 18216
rect 30834 18164 30840 18216
rect 30892 18164 30898 18216
rect 31294 18164 31300 18216
rect 31352 18164 31358 18216
rect 32950 18164 32956 18216
rect 33008 18164 33014 18216
rect 33428 18213 33456 18244
rect 33502 18232 33508 18284
rect 33560 18232 33566 18284
rect 33686 18232 33692 18284
rect 33744 18232 33750 18284
rect 33413 18207 33471 18213
rect 33413 18173 33425 18207
rect 33459 18173 33471 18207
rect 33413 18167 33471 18173
rect 26053 18099 26111 18105
rect 26988 18108 27200 18136
rect 27709 18139 27767 18145
rect 26988 18080 27016 18108
rect 27709 18105 27721 18139
rect 27755 18136 27767 18139
rect 27982 18136 27988 18148
rect 27755 18108 27988 18136
rect 27755 18105 27767 18108
rect 27709 18099 27767 18105
rect 27982 18096 27988 18108
rect 28040 18096 28046 18148
rect 28288 18139 28346 18145
rect 28288 18136 28300 18139
rect 28092 18108 28300 18136
rect 13044 18040 16252 18068
rect 13044 18028 13050 18040
rect 17126 18028 17132 18080
rect 17184 18028 17190 18080
rect 17218 18028 17224 18080
rect 17276 18028 17282 18080
rect 17678 18028 17684 18080
rect 17736 18068 17742 18080
rect 17957 18071 18015 18077
rect 17957 18068 17969 18071
rect 17736 18040 17969 18068
rect 17736 18028 17742 18040
rect 17957 18037 17969 18040
rect 18003 18037 18015 18071
rect 17957 18031 18015 18037
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 18325 18071 18383 18077
rect 18325 18068 18337 18071
rect 18104 18040 18337 18068
rect 18104 18028 18110 18040
rect 18325 18037 18337 18040
rect 18371 18037 18383 18071
rect 18325 18031 18383 18037
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 19981 18071 20039 18077
rect 19981 18068 19993 18071
rect 18656 18040 19993 18068
rect 18656 18028 18662 18040
rect 19981 18037 19993 18040
rect 20027 18037 20039 18071
rect 19981 18031 20039 18037
rect 20530 18028 20536 18080
rect 20588 18028 20594 18080
rect 22186 18028 22192 18080
rect 22244 18068 22250 18080
rect 23661 18071 23719 18077
rect 23661 18068 23673 18071
rect 22244 18040 23673 18068
rect 22244 18028 22250 18040
rect 23661 18037 23673 18040
rect 23707 18068 23719 18071
rect 24213 18071 24271 18077
rect 24213 18068 24225 18071
rect 23707 18040 24225 18068
rect 23707 18037 23719 18040
rect 23661 18031 23719 18037
rect 24213 18037 24225 18040
rect 24259 18037 24271 18071
rect 24213 18031 24271 18037
rect 24946 18028 24952 18080
rect 25004 18028 25010 18080
rect 26878 18028 26884 18080
rect 26936 18028 26942 18080
rect 26970 18028 26976 18080
rect 27028 18028 27034 18080
rect 27062 18028 27068 18080
rect 27120 18068 27126 18080
rect 28092 18068 28120 18108
rect 28288 18105 28300 18108
rect 28334 18136 28346 18139
rect 28905 18139 28963 18145
rect 28905 18136 28917 18139
rect 28334 18108 28488 18136
rect 28334 18105 28346 18108
rect 28288 18099 28346 18105
rect 28460 18080 28488 18108
rect 28828 18108 28917 18136
rect 28828 18080 28856 18108
rect 28905 18105 28917 18108
rect 28951 18105 28963 18139
rect 28905 18099 28963 18105
rect 29273 18139 29331 18145
rect 29273 18105 29285 18139
rect 29319 18136 29331 18139
rect 29362 18136 29368 18148
rect 29319 18108 29368 18136
rect 29319 18105 29331 18108
rect 29273 18099 29331 18105
rect 29362 18096 29368 18108
rect 29420 18096 29426 18148
rect 29546 18096 29552 18148
rect 29604 18136 29610 18148
rect 29825 18139 29883 18145
rect 29825 18136 29837 18139
rect 29604 18108 29837 18136
rect 29604 18096 29610 18108
rect 29825 18105 29837 18108
rect 29871 18105 29883 18139
rect 29825 18099 29883 18105
rect 30469 18139 30527 18145
rect 30469 18105 30481 18139
rect 30515 18136 30527 18139
rect 30558 18136 30564 18148
rect 30515 18108 30564 18136
rect 30515 18105 30527 18108
rect 30469 18099 30527 18105
rect 30558 18096 30564 18108
rect 30616 18096 30622 18148
rect 30685 18139 30743 18145
rect 30685 18105 30697 18139
rect 30731 18136 30743 18139
rect 30852 18136 30880 18164
rect 30731 18108 30880 18136
rect 30731 18105 30743 18108
rect 30685 18099 30743 18105
rect 27120 18040 28120 18068
rect 27120 18028 27126 18040
rect 28442 18028 28448 18080
rect 28500 18028 28506 18080
rect 28718 18028 28724 18080
rect 28776 18028 28782 18080
rect 28810 18028 28816 18080
rect 28868 18028 28874 18080
rect 29181 18071 29239 18077
rect 29181 18037 29193 18071
rect 29227 18068 29239 18071
rect 29454 18068 29460 18080
rect 29227 18040 29460 18068
rect 29227 18037 29239 18040
rect 29181 18031 29239 18037
rect 29454 18028 29460 18040
rect 29512 18028 29518 18080
rect 29733 18071 29791 18077
rect 29733 18037 29745 18071
rect 29779 18068 29791 18071
rect 29914 18068 29920 18080
rect 29779 18040 29920 18068
rect 29779 18037 29791 18040
rect 29733 18031 29791 18037
rect 29914 18028 29920 18040
rect 29972 18028 29978 18080
rect 30098 18028 30104 18080
rect 30156 18028 30162 18080
rect 31205 18071 31263 18077
rect 31205 18037 31217 18071
rect 31251 18068 31263 18071
rect 31312 18068 31340 18164
rect 32030 18096 32036 18148
rect 32088 18096 32094 18148
rect 32398 18096 32404 18148
rect 32456 18136 32462 18148
rect 32677 18139 32735 18145
rect 32677 18136 32689 18139
rect 32456 18108 32689 18136
rect 32456 18096 32462 18108
rect 32677 18105 32689 18108
rect 32723 18105 32735 18139
rect 32677 18099 32735 18105
rect 31251 18040 31340 18068
rect 33045 18071 33103 18077
rect 31251 18037 31263 18040
rect 31205 18031 31263 18037
rect 33045 18037 33057 18071
rect 33091 18068 33103 18071
rect 33594 18068 33600 18080
rect 33091 18040 33600 18068
rect 33091 18037 33103 18040
rect 33045 18031 33103 18037
rect 33594 18028 33600 18040
rect 33652 18028 33658 18080
rect 2760 17978 34316 18000
rect 2760 17926 7210 17978
rect 7262 17926 7274 17978
rect 7326 17926 7338 17978
rect 7390 17926 7402 17978
rect 7454 17926 7466 17978
rect 7518 17926 15099 17978
rect 15151 17926 15163 17978
rect 15215 17926 15227 17978
rect 15279 17926 15291 17978
rect 15343 17926 15355 17978
rect 15407 17926 22988 17978
rect 23040 17926 23052 17978
rect 23104 17926 23116 17978
rect 23168 17926 23180 17978
rect 23232 17926 23244 17978
rect 23296 17926 30877 17978
rect 30929 17926 30941 17978
rect 30993 17926 31005 17978
rect 31057 17926 31069 17978
rect 31121 17926 31133 17978
rect 31185 17926 34316 17978
rect 2760 17904 34316 17926
rect 4985 17867 5043 17873
rect 4985 17833 4997 17867
rect 5031 17864 5043 17867
rect 5442 17864 5448 17876
rect 5031 17836 5448 17864
rect 5031 17833 5043 17836
rect 4985 17827 5043 17833
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 9122 17864 9128 17876
rect 8312 17836 9128 17864
rect 6914 17756 6920 17808
rect 6972 17756 6978 17808
rect 8312 17805 8340 17836
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 18874 17864 18880 17876
rect 12406 17836 18880 17864
rect 8297 17799 8355 17805
rect 8297 17765 8309 17799
rect 8343 17765 8355 17799
rect 9582 17796 9588 17808
rect 9522 17768 9588 17796
rect 8297 17759 8355 17765
rect 9582 17756 9588 17768
rect 9640 17756 9646 17808
rect 12161 17799 12219 17805
rect 12161 17765 12173 17799
rect 12207 17796 12219 17799
rect 12406 17796 12434 17836
rect 18874 17824 18880 17836
rect 18932 17864 18938 17876
rect 20898 17864 20904 17876
rect 18932 17836 20904 17864
rect 18932 17824 18938 17836
rect 20898 17824 20904 17836
rect 20956 17824 20962 17876
rect 22649 17867 22707 17873
rect 22649 17833 22661 17867
rect 22695 17833 22707 17867
rect 22649 17827 22707 17833
rect 12207 17768 12434 17796
rect 12207 17765 12219 17768
rect 12161 17759 12219 17765
rect 12894 17756 12900 17808
rect 12952 17756 12958 17808
rect 13446 17756 13452 17808
rect 13504 17756 13510 17808
rect 15841 17799 15899 17805
rect 15841 17796 15853 17799
rect 14674 17768 15853 17796
rect 15841 17765 15853 17768
rect 15887 17765 15899 17799
rect 15841 17759 15899 17765
rect 16022 17756 16028 17808
rect 16080 17756 16086 17808
rect 16114 17756 16120 17808
rect 16172 17796 16178 17808
rect 16853 17799 16911 17805
rect 16853 17796 16865 17799
rect 16172 17768 16865 17796
rect 16172 17756 16178 17768
rect 16853 17765 16865 17768
rect 16899 17796 16911 17799
rect 17402 17796 17408 17808
rect 16899 17768 17408 17796
rect 16899 17765 16911 17768
rect 16853 17759 16911 17765
rect 17402 17756 17408 17768
rect 17460 17756 17466 17808
rect 17770 17756 17776 17808
rect 17828 17756 17834 17808
rect 17862 17756 17868 17808
rect 17920 17756 17926 17808
rect 18969 17799 19027 17805
rect 18969 17796 18981 17799
rect 18156 17768 18981 17796
rect 3418 17688 3424 17740
rect 3476 17688 3482 17740
rect 5350 17688 5356 17740
rect 5408 17688 5414 17740
rect 12986 17728 12992 17740
rect 9508 17700 12388 17728
rect 4522 17620 4528 17672
rect 4580 17620 4586 17672
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17629 4859 17663
rect 4801 17623 4859 17629
rect 3050 17484 3056 17536
rect 3108 17484 3114 17536
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 4816 17524 4844 17623
rect 6362 17620 6368 17672
rect 6420 17660 6426 17672
rect 6457 17663 6515 17669
rect 6457 17660 6469 17663
rect 6420 17632 6469 17660
rect 6420 17620 6426 17632
rect 6457 17629 6469 17632
rect 6503 17629 6515 17663
rect 6457 17623 6515 17629
rect 6733 17663 6791 17669
rect 6733 17629 6745 17663
rect 6779 17660 6791 17663
rect 8021 17663 8079 17669
rect 8021 17660 8033 17663
rect 6779 17632 8033 17660
rect 6779 17629 6791 17632
rect 6733 17623 6791 17629
rect 8021 17629 8033 17632
rect 8067 17629 8079 17663
rect 9508 17660 9536 17700
rect 12360 17672 12388 17700
rect 12452 17700 12992 17728
rect 8021 17623 8079 17629
rect 8128 17632 9536 17660
rect 6454 17524 6460 17536
rect 4212 17496 6460 17524
rect 4212 17484 4218 17496
rect 6454 17484 6460 17496
rect 6512 17524 6518 17536
rect 6748 17524 6776 17623
rect 7098 17552 7104 17604
rect 7156 17592 7162 17604
rect 8128 17592 8156 17632
rect 12250 17620 12256 17672
rect 12308 17620 12314 17672
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12452 17660 12480 17700
rect 12986 17688 12992 17700
rect 13044 17688 13050 17740
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 13173 17731 13231 17737
rect 13173 17728 13185 17731
rect 13136 17700 13185 17728
rect 13136 17688 13142 17700
rect 13173 17697 13185 17700
rect 13219 17697 13231 17731
rect 15749 17731 15807 17737
rect 15749 17728 15761 17731
rect 13173 17691 13231 17697
rect 14844 17700 15761 17728
rect 14844 17672 14872 17700
rect 15749 17697 15761 17700
rect 15795 17697 15807 17731
rect 15749 17691 15807 17697
rect 17313 17731 17371 17737
rect 17313 17697 17325 17731
rect 17359 17728 17371 17731
rect 17880 17728 17908 17756
rect 17359 17700 17908 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 12400 17632 12480 17660
rect 13280 17632 14780 17660
rect 12400 17620 12406 17632
rect 13280 17592 13308 17632
rect 7156 17564 8156 17592
rect 9324 17564 13308 17592
rect 14752 17592 14780 17632
rect 14826 17620 14832 17672
rect 14884 17620 14890 17672
rect 14921 17663 14979 17669
rect 14921 17629 14933 17663
rect 14967 17660 14979 17663
rect 15013 17663 15071 17669
rect 15013 17660 15025 17663
rect 14967 17632 15025 17660
rect 14967 17629 14979 17632
rect 14921 17623 14979 17629
rect 15013 17629 15025 17632
rect 15059 17629 15071 17663
rect 16574 17660 16580 17672
rect 15013 17623 15071 17629
rect 15580 17632 16580 17660
rect 15580 17592 15608 17632
rect 16574 17620 16580 17632
rect 16632 17660 16638 17672
rect 16850 17660 16856 17672
rect 16632 17632 16856 17660
rect 16632 17620 16638 17632
rect 16850 17620 16856 17632
rect 16908 17620 16914 17672
rect 17218 17620 17224 17672
rect 17276 17620 17282 17672
rect 17586 17620 17592 17672
rect 17644 17660 17650 17672
rect 18156 17660 18184 17768
rect 18969 17765 18981 17768
rect 19015 17765 19027 17799
rect 18969 17759 19027 17765
rect 20806 17756 20812 17808
rect 20864 17796 20870 17808
rect 21910 17796 21916 17808
rect 20864 17768 21916 17796
rect 20864 17756 20870 17768
rect 21910 17756 21916 17768
rect 21968 17796 21974 17808
rect 22664 17796 22692 17827
rect 22738 17824 22744 17876
rect 22796 17864 22802 17876
rect 23290 17864 23296 17876
rect 22796 17836 23296 17864
rect 22796 17824 22802 17836
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 26878 17864 26884 17876
rect 26252 17836 26884 17864
rect 21968 17768 22692 17796
rect 21968 17756 21974 17768
rect 18230 17688 18236 17740
rect 18288 17728 18294 17740
rect 18509 17731 18567 17737
rect 18509 17728 18521 17731
rect 18288 17700 18521 17728
rect 18288 17688 18294 17700
rect 18509 17697 18521 17700
rect 18555 17697 18567 17731
rect 19058 17728 19064 17740
rect 18509 17691 18567 17697
rect 18616 17700 19064 17728
rect 17644 17632 18184 17660
rect 17644 17620 17650 17632
rect 18322 17620 18328 17672
rect 18380 17660 18386 17672
rect 18616 17660 18644 17700
rect 19058 17688 19064 17700
rect 19116 17688 19122 17740
rect 19518 17688 19524 17740
rect 19576 17688 19582 17740
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17728 19763 17731
rect 20165 17731 20223 17737
rect 20165 17728 20177 17731
rect 19751 17700 20177 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 20165 17697 20177 17700
rect 20211 17697 20223 17731
rect 20165 17691 20223 17697
rect 20530 17688 20536 17740
rect 20588 17728 20594 17740
rect 20625 17731 20683 17737
rect 20625 17728 20637 17731
rect 20588 17700 20637 17728
rect 20588 17688 20594 17700
rect 20625 17697 20637 17700
rect 20671 17697 20683 17731
rect 20625 17691 20683 17697
rect 20901 17731 20959 17737
rect 20901 17697 20913 17731
rect 20947 17728 20959 17731
rect 21266 17728 21272 17740
rect 20947 17700 21272 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 21361 17731 21419 17737
rect 21361 17697 21373 17731
rect 21407 17728 21419 17731
rect 21634 17728 21640 17740
rect 21407 17700 21640 17728
rect 21407 17697 21419 17700
rect 21361 17691 21419 17697
rect 21634 17688 21640 17700
rect 21692 17688 21698 17740
rect 22664 17728 22692 17768
rect 24210 17756 24216 17808
rect 24268 17756 24274 17808
rect 26252 17805 26280 17836
rect 26878 17824 26884 17836
rect 26936 17824 26942 17876
rect 27709 17867 27767 17873
rect 27709 17833 27721 17867
rect 27755 17864 27767 17867
rect 28258 17864 28264 17876
rect 27755 17836 28264 17864
rect 27755 17833 27767 17836
rect 27709 17827 27767 17833
rect 28258 17824 28264 17836
rect 28316 17824 28322 17876
rect 29362 17864 29368 17876
rect 28368 17836 29368 17864
rect 26237 17799 26295 17805
rect 26237 17765 26249 17799
rect 26283 17765 26295 17799
rect 28074 17796 28080 17808
rect 27462 17768 28080 17796
rect 26237 17759 26295 17765
rect 28074 17756 28080 17768
rect 28132 17756 28138 17808
rect 23477 17731 23535 17737
rect 23477 17728 23489 17731
rect 22664 17700 23489 17728
rect 23477 17697 23489 17700
rect 23523 17697 23535 17731
rect 23477 17691 23535 17697
rect 27614 17688 27620 17740
rect 27672 17688 27678 17740
rect 28169 17731 28227 17737
rect 28169 17697 28181 17731
rect 28215 17728 28227 17731
rect 28258 17728 28264 17740
rect 28215 17700 28264 17728
rect 28215 17697 28227 17700
rect 28169 17691 28227 17697
rect 28258 17688 28264 17700
rect 28316 17688 28322 17740
rect 28368 17728 28396 17836
rect 29362 17824 29368 17836
rect 29420 17824 29426 17876
rect 30098 17824 30104 17876
rect 30156 17824 30162 17876
rect 31757 17867 31815 17873
rect 31757 17833 31769 17867
rect 31803 17864 31815 17867
rect 32398 17864 32404 17876
rect 31803 17836 32404 17864
rect 31803 17833 31815 17836
rect 31757 17827 31815 17833
rect 32398 17824 32404 17836
rect 32456 17824 32462 17876
rect 33502 17824 33508 17876
rect 33560 17864 33566 17876
rect 33597 17867 33655 17873
rect 33597 17864 33609 17867
rect 33560 17836 33609 17864
rect 33560 17824 33566 17836
rect 33597 17833 33609 17836
rect 33643 17833 33655 17867
rect 33597 17827 33655 17833
rect 28445 17731 28503 17737
rect 28445 17728 28457 17731
rect 28368 17700 28457 17728
rect 28445 17697 28457 17700
rect 28491 17697 28503 17731
rect 28445 17691 28503 17697
rect 28534 17688 28540 17740
rect 28592 17728 28598 17740
rect 28592 17700 29316 17728
rect 28592 17688 28598 17700
rect 18380 17632 18644 17660
rect 18693 17663 18751 17669
rect 18380 17620 18386 17632
rect 18693 17629 18705 17663
rect 18739 17660 18751 17663
rect 19242 17660 19248 17672
rect 18739 17632 19248 17660
rect 18739 17629 18751 17632
rect 18693 17623 18751 17629
rect 17236 17592 17264 17620
rect 14752 17564 15608 17592
rect 15672 17564 17264 17592
rect 7156 17552 7162 17564
rect 6512 17496 6776 17524
rect 6512 17484 6518 17496
rect 7650 17484 7656 17536
rect 7708 17524 7714 17536
rect 7745 17527 7803 17533
rect 7745 17524 7757 17527
rect 7708 17496 7757 17524
rect 7708 17484 7714 17496
rect 7745 17493 7757 17496
rect 7791 17524 7803 17527
rect 9324 17524 9352 17564
rect 7791 17496 9352 17524
rect 7791 17493 7803 17496
rect 7745 17487 7803 17493
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 10502 17524 10508 17536
rect 9824 17496 10508 17524
rect 9824 17484 9830 17496
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 10873 17527 10931 17533
rect 10873 17493 10885 17527
rect 10919 17524 10931 17527
rect 11054 17524 11060 17536
rect 10919 17496 11060 17524
rect 10919 17493 10931 17496
rect 10873 17487 10931 17493
rect 11054 17484 11060 17496
rect 11112 17484 11118 17536
rect 15470 17484 15476 17536
rect 15528 17524 15534 17536
rect 15672 17533 15700 17564
rect 17678 17552 17684 17604
rect 17736 17592 17742 17604
rect 17773 17595 17831 17601
rect 17773 17592 17785 17595
rect 17736 17564 17785 17592
rect 17736 17552 17742 17564
rect 17773 17561 17785 17564
rect 17819 17561 17831 17595
rect 18708 17592 18736 17623
rect 19242 17620 19248 17632
rect 19300 17620 19306 17672
rect 19337 17663 19395 17669
rect 19337 17629 19349 17663
rect 19383 17660 19395 17663
rect 20070 17660 20076 17672
rect 19383 17632 20076 17660
rect 19383 17629 19395 17632
rect 19337 17623 19395 17629
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20254 17620 20260 17672
rect 20312 17620 20318 17672
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17629 20499 17663
rect 23014 17660 23020 17672
rect 20441 17623 20499 17629
rect 20916 17632 23020 17660
rect 17773 17555 17831 17561
rect 17880 17564 18736 17592
rect 17880 17536 17908 17564
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15528 17496 15669 17524
rect 15528 17484 15534 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 16666 17484 16672 17536
rect 16724 17524 16730 17536
rect 17037 17527 17095 17533
rect 17037 17524 17049 17527
rect 16724 17496 17049 17524
rect 16724 17484 16730 17496
rect 17037 17493 17049 17496
rect 17083 17493 17095 17527
rect 17037 17487 17095 17493
rect 17126 17484 17132 17536
rect 17184 17524 17190 17536
rect 17862 17524 17868 17536
rect 17184 17496 17868 17524
rect 17184 17484 17190 17496
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 18322 17484 18328 17536
rect 18380 17484 18386 17536
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 18509 17527 18567 17533
rect 18509 17524 18521 17527
rect 18472 17496 18521 17524
rect 18472 17484 18478 17496
rect 18509 17493 18521 17496
rect 18555 17493 18567 17527
rect 18509 17487 18567 17493
rect 19794 17484 19800 17536
rect 19852 17484 19858 17536
rect 20088 17524 20116 17620
rect 20456 17592 20484 17623
rect 20916 17592 20944 17632
rect 23014 17620 23020 17632
rect 23072 17620 23078 17672
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17660 23811 17663
rect 24946 17660 24952 17672
rect 23799 17632 24952 17660
rect 23799 17629 23811 17632
rect 23753 17623 23811 17629
rect 24946 17620 24952 17632
rect 25004 17620 25010 17672
rect 25961 17663 26019 17669
rect 25961 17629 25973 17663
rect 26007 17629 26019 17663
rect 25961 17623 26019 17629
rect 20456 17564 20944 17592
rect 20990 17524 20996 17536
rect 20088 17496 20996 17524
rect 20990 17484 20996 17496
rect 21048 17484 21054 17536
rect 21266 17484 21272 17536
rect 21324 17524 21330 17536
rect 23474 17524 23480 17536
rect 21324 17496 23480 17524
rect 21324 17484 21330 17496
rect 23474 17484 23480 17496
rect 23532 17484 23538 17536
rect 25222 17484 25228 17536
rect 25280 17484 25286 17536
rect 25976 17524 26004 17623
rect 27632 17592 27660 17688
rect 28353 17663 28411 17669
rect 28353 17629 28365 17663
rect 28399 17660 28411 17663
rect 28399 17632 28764 17660
rect 28399 17629 28411 17632
rect 28353 17623 28411 17629
rect 27985 17595 28043 17601
rect 27985 17592 27997 17595
rect 27632 17564 27997 17592
rect 27985 17561 27997 17564
rect 28031 17561 28043 17595
rect 27985 17555 28043 17561
rect 27614 17524 27620 17536
rect 25976 17496 27620 17524
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 28445 17527 28503 17533
rect 28445 17493 28457 17527
rect 28491 17524 28503 17527
rect 28534 17524 28540 17536
rect 28491 17496 28540 17524
rect 28491 17493 28503 17496
rect 28445 17487 28503 17493
rect 28534 17484 28540 17496
rect 28592 17484 28598 17536
rect 28626 17484 28632 17536
rect 28684 17484 28690 17536
rect 28736 17524 28764 17632
rect 29178 17620 29184 17672
rect 29236 17620 29242 17672
rect 29288 17660 29316 17700
rect 29362 17688 29368 17740
rect 29420 17688 29426 17740
rect 29549 17731 29607 17737
rect 29549 17697 29561 17731
rect 29595 17728 29607 17731
rect 29914 17728 29920 17740
rect 29595 17700 29920 17728
rect 29595 17697 29607 17700
rect 29549 17691 29607 17697
rect 29914 17688 29920 17700
rect 29972 17688 29978 17740
rect 30122 17737 30150 17824
rect 30650 17796 30656 17808
rect 30300 17768 30656 17796
rect 30300 17737 30328 17768
rect 30650 17756 30656 17768
rect 30708 17756 30714 17808
rect 33873 17799 33931 17805
rect 33873 17796 33885 17799
rect 33350 17768 33885 17796
rect 33873 17765 33885 17768
rect 33919 17765 33931 17799
rect 33873 17759 33931 17765
rect 30101 17731 30159 17737
rect 30101 17697 30113 17731
rect 30147 17697 30159 17731
rect 30101 17691 30159 17697
rect 30285 17731 30343 17737
rect 30285 17697 30297 17731
rect 30331 17697 30343 17731
rect 30285 17691 30343 17697
rect 29638 17660 29644 17672
rect 29288 17632 29644 17660
rect 29638 17620 29644 17632
rect 29696 17620 29702 17672
rect 29822 17620 29828 17672
rect 29880 17660 29886 17672
rect 30300 17660 30328 17691
rect 31202 17688 31208 17740
rect 31260 17688 31266 17740
rect 33134 17688 33140 17740
rect 33192 17688 33198 17740
rect 33781 17731 33839 17737
rect 33781 17697 33793 17731
rect 33827 17697 33839 17731
rect 33781 17691 33839 17697
rect 29880 17632 30328 17660
rect 30469 17663 30527 17669
rect 29880 17620 29886 17632
rect 30469 17629 30481 17663
rect 30515 17660 30527 17663
rect 30650 17660 30656 17672
rect 30515 17632 30656 17660
rect 30515 17629 30527 17632
rect 30469 17623 30527 17629
rect 30650 17620 30656 17632
rect 30708 17620 30714 17672
rect 31849 17663 31907 17669
rect 31849 17660 31861 17663
rect 31726 17632 31861 17660
rect 28902 17552 28908 17604
rect 28960 17592 28966 17604
rect 31726 17592 31754 17632
rect 31849 17629 31861 17632
rect 31895 17629 31907 17663
rect 31849 17623 31907 17629
rect 32122 17620 32128 17672
rect 32180 17620 32186 17672
rect 33152 17660 33180 17688
rect 33796 17660 33824 17691
rect 33152 17632 33824 17660
rect 28960 17564 31754 17592
rect 28960 17552 28966 17564
rect 29454 17524 29460 17536
rect 28736 17496 29460 17524
rect 29454 17484 29460 17496
rect 29512 17484 29518 17536
rect 29546 17484 29552 17536
rect 29604 17484 29610 17536
rect 30193 17527 30251 17533
rect 30193 17493 30205 17527
rect 30239 17524 30251 17527
rect 30742 17524 30748 17536
rect 30239 17496 30748 17524
rect 30239 17493 30251 17496
rect 30193 17487 30251 17493
rect 30742 17484 30748 17496
rect 30800 17484 30806 17536
rect 31018 17484 31024 17536
rect 31076 17484 31082 17536
rect 2760 17434 34316 17456
rect 2760 17382 6550 17434
rect 6602 17382 6614 17434
rect 6666 17382 6678 17434
rect 6730 17382 6742 17434
rect 6794 17382 6806 17434
rect 6858 17382 14439 17434
rect 14491 17382 14503 17434
rect 14555 17382 14567 17434
rect 14619 17382 14631 17434
rect 14683 17382 14695 17434
rect 14747 17382 22328 17434
rect 22380 17382 22392 17434
rect 22444 17382 22456 17434
rect 22508 17382 22520 17434
rect 22572 17382 22584 17434
rect 22636 17382 30217 17434
rect 30269 17382 30281 17434
rect 30333 17382 30345 17434
rect 30397 17382 30409 17434
rect 30461 17382 30473 17434
rect 30525 17382 34316 17434
rect 2760 17360 34316 17382
rect 3050 17280 3056 17332
rect 3108 17280 3114 17332
rect 5537 17323 5595 17329
rect 5537 17289 5549 17323
rect 5583 17320 5595 17323
rect 6086 17320 6092 17332
rect 5583 17292 6092 17320
rect 5583 17289 5595 17292
rect 5537 17283 5595 17289
rect 3068 17116 3096 17280
rect 4338 17144 4344 17196
rect 4396 17184 4402 17196
rect 5074 17184 5080 17196
rect 4396 17156 5080 17184
rect 4396 17144 4402 17156
rect 5074 17144 5080 17156
rect 5132 17144 5138 17196
rect 4249 17119 4307 17125
rect 4249 17116 4261 17119
rect 3068 17088 4261 17116
rect 4249 17085 4261 17088
rect 4295 17116 4307 17119
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 4295 17088 4997 17116
rect 4295 17085 4307 17088
rect 4249 17079 4307 17085
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 1302 17008 1308 17060
rect 1360 17048 1366 17060
rect 3237 17051 3295 17057
rect 3237 17048 3249 17051
rect 1360 17020 3249 17048
rect 1360 17008 1366 17020
rect 3237 17017 3249 17020
rect 3283 17017 3295 17051
rect 3237 17011 3295 17017
rect 4893 17051 4951 17057
rect 4893 17017 4905 17051
rect 4939 17048 4951 17051
rect 5552 17048 5580 17283
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 6273 17323 6331 17329
rect 6273 17289 6285 17323
rect 6319 17320 6331 17323
rect 6362 17320 6368 17332
rect 6319 17292 6368 17320
rect 6319 17289 6331 17292
rect 6273 17283 6331 17289
rect 6362 17280 6368 17292
rect 6420 17280 6426 17332
rect 9582 17280 9588 17332
rect 9640 17280 9646 17332
rect 12158 17320 12164 17332
rect 10704 17292 12164 17320
rect 6454 17212 6460 17264
rect 6512 17252 6518 17264
rect 6512 17224 6960 17252
rect 6512 17212 6518 17224
rect 6178 17144 6184 17196
rect 6236 17144 6242 17196
rect 6362 17144 6368 17196
rect 6420 17184 6426 17196
rect 6932 17193 6960 17224
rect 8202 17212 8208 17264
rect 8260 17252 8266 17264
rect 10704 17252 10732 17292
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12250 17280 12256 17332
rect 12308 17320 12314 17332
rect 12345 17323 12403 17329
rect 12345 17320 12357 17323
rect 12308 17292 12357 17320
rect 12308 17280 12314 17292
rect 12345 17289 12357 17292
rect 12391 17289 12403 17323
rect 12345 17283 12403 17289
rect 13446 17280 13452 17332
rect 13504 17320 13510 17332
rect 13817 17323 13875 17329
rect 13817 17320 13829 17323
rect 13504 17292 13829 17320
rect 13504 17280 13510 17292
rect 13817 17289 13829 17292
rect 13863 17289 13875 17323
rect 15010 17320 15016 17332
rect 13817 17283 13875 17289
rect 14200 17292 15016 17320
rect 13722 17252 13728 17264
rect 8260 17224 10732 17252
rect 12636 17224 13728 17252
rect 8260 17212 8266 17224
rect 6917 17187 6975 17193
rect 6420 17156 6500 17184
rect 6420 17144 6426 17156
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6472 17125 6500 17156
rect 6917 17153 6929 17187
rect 6963 17153 6975 17187
rect 6917 17147 6975 17153
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17184 7251 17187
rect 8757 17187 8815 17193
rect 8757 17184 8769 17187
rect 7239 17156 8769 17184
rect 7239 17153 7251 17156
rect 7193 17147 7251 17153
rect 8757 17153 8769 17156
rect 8803 17153 8815 17187
rect 8757 17147 8815 17153
rect 10870 17144 10876 17196
rect 10928 17144 10934 17196
rect 12636 17193 12664 17224
rect 13722 17212 13728 17224
rect 13780 17212 13786 17264
rect 14200 17196 14228 17292
rect 15010 17280 15016 17292
rect 15068 17280 15074 17332
rect 18322 17280 18328 17332
rect 18380 17280 18386 17332
rect 18601 17323 18659 17329
rect 18601 17289 18613 17323
rect 18647 17320 18659 17323
rect 18782 17320 18788 17332
rect 18647 17292 18788 17320
rect 18647 17289 18659 17292
rect 18601 17283 18659 17289
rect 18782 17280 18788 17292
rect 18840 17280 18846 17332
rect 20254 17280 20260 17332
rect 20312 17280 20318 17332
rect 21453 17323 21511 17329
rect 21453 17289 21465 17323
rect 21499 17320 21511 17323
rect 21542 17320 21548 17332
rect 21499 17292 21548 17320
rect 21499 17289 21511 17292
rect 21453 17283 21511 17289
rect 21542 17280 21548 17292
rect 21600 17280 21606 17332
rect 22830 17320 22836 17332
rect 21652 17292 22836 17320
rect 15470 17252 15476 17264
rect 14292 17224 15476 17252
rect 12621 17187 12679 17193
rect 12621 17153 12633 17187
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12713 17187 12771 17193
rect 12713 17153 12725 17187
rect 12759 17184 12771 17187
rect 12894 17184 12900 17196
rect 12759 17156 12900 17184
rect 12759 17153 12771 17156
rect 12713 17147 12771 17153
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13633 17187 13691 17193
rect 13633 17153 13645 17187
rect 13679 17184 13691 17187
rect 14182 17184 14188 17196
rect 13679 17156 14188 17184
rect 13679 17153 13691 17156
rect 13633 17147 13691 17153
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 14292 17193 14320 17224
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 14366 17144 14372 17196
rect 14424 17144 14430 17196
rect 16390 17184 16396 17196
rect 15764 17156 16396 17184
rect 6457 17119 6515 17125
rect 5960 17088 6408 17116
rect 5960 17076 5966 17088
rect 4939 17020 5580 17048
rect 4939 17017 4951 17020
rect 4893 17011 4951 17017
rect 6270 17008 6276 17060
rect 6328 17008 6334 17060
rect 6380 17048 6408 17088
rect 6457 17085 6469 17119
rect 6503 17085 6515 17119
rect 6457 17079 6515 17085
rect 6549 17119 6607 17125
rect 6549 17085 6561 17119
rect 6595 17085 6607 17119
rect 6549 17079 6607 17085
rect 6564 17048 6592 17079
rect 6822 17076 6828 17128
rect 6880 17076 6886 17128
rect 9306 17076 9312 17128
rect 9364 17076 9370 17128
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 10229 17119 10287 17125
rect 10229 17116 10241 17119
rect 9732 17088 10241 17116
rect 9732 17076 9738 17088
rect 10229 17085 10241 17088
rect 10275 17116 10287 17119
rect 10410 17116 10416 17128
rect 10275 17088 10416 17116
rect 10275 17085 10287 17088
rect 10229 17079 10287 17085
rect 10410 17076 10416 17088
rect 10468 17076 10474 17128
rect 10597 17119 10655 17125
rect 10597 17085 10609 17119
rect 10643 17085 10655 17119
rect 14826 17116 14832 17128
rect 10597 17079 10655 17085
rect 13924 17088 14832 17116
rect 6380 17020 6592 17048
rect 6641 17051 6699 17057
rect 6641 17017 6653 17051
rect 6687 17017 6699 17051
rect 6641 17011 6699 17017
rect 4525 16983 4583 16989
rect 4525 16949 4537 16983
rect 4571 16980 4583 16983
rect 4798 16980 4804 16992
rect 4571 16952 4804 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 6288 16980 6316 17008
rect 6656 16980 6684 17011
rect 6288 16952 6684 16980
rect 6840 16980 6868 17076
rect 7742 17008 7748 17060
rect 7800 17008 7806 17060
rect 10612 17048 10640 17079
rect 8588 17020 9674 17048
rect 8588 16980 8616 17020
rect 6840 16952 8616 16980
rect 8662 16940 8668 16992
rect 8720 16940 8726 16992
rect 9646 16980 9674 17020
rect 10244 17020 10640 17048
rect 10796 17020 11362 17048
rect 10244 16992 10272 17020
rect 9858 16980 9864 16992
rect 9646 16952 9864 16980
rect 9858 16940 9864 16952
rect 9916 16980 9922 16992
rect 9953 16983 10011 16989
rect 9953 16980 9965 16983
rect 9916 16952 9965 16980
rect 9916 16940 9922 16952
rect 9953 16949 9965 16952
rect 9999 16949 10011 16983
rect 9953 16943 10011 16949
rect 10226 16940 10232 16992
rect 10284 16940 10290 16992
rect 10321 16983 10379 16989
rect 10321 16949 10333 16983
rect 10367 16980 10379 16983
rect 10796 16980 10824 17020
rect 12802 17008 12808 17060
rect 12860 17008 12866 17060
rect 13814 17048 13820 17060
rect 13188 17020 13820 17048
rect 13188 16989 13216 17020
rect 13814 17008 13820 17020
rect 13872 17008 13878 17060
rect 13924 16992 13952 17088
rect 14826 17076 14832 17088
rect 14884 17076 14890 17128
rect 15562 17076 15568 17128
rect 15620 17076 15626 17128
rect 15764 17125 15792 17156
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 18138 17144 18144 17196
rect 18196 17193 18202 17196
rect 18196 17187 18224 17193
rect 18212 17153 18224 17187
rect 18340 17184 18368 17280
rect 18509 17255 18567 17261
rect 18509 17221 18521 17255
rect 18555 17252 18567 17255
rect 20272 17252 20300 17280
rect 21652 17252 21680 17292
rect 22830 17280 22836 17292
rect 22888 17320 22894 17332
rect 23017 17323 23075 17329
rect 23017 17320 23029 17323
rect 22888 17292 23029 17320
rect 22888 17280 22894 17292
rect 23017 17289 23029 17292
rect 23063 17289 23075 17323
rect 23017 17283 23075 17289
rect 25222 17280 25228 17332
rect 25280 17320 25286 17332
rect 26602 17320 26608 17332
rect 25280 17292 26608 17320
rect 25280 17280 25286 17292
rect 26602 17280 26608 17292
rect 26660 17280 26666 17332
rect 26712 17292 29040 17320
rect 22278 17252 22284 17264
rect 18555 17224 18644 17252
rect 20272 17224 21680 17252
rect 21744 17224 22284 17252
rect 18555 17221 18567 17224
rect 18509 17215 18567 17221
rect 18340 17156 18460 17184
rect 18196 17147 18224 17153
rect 18196 17144 18202 17147
rect 15749 17119 15807 17125
rect 15749 17085 15761 17119
rect 15795 17085 15807 17119
rect 15749 17079 15807 17085
rect 17586 17076 17592 17128
rect 17644 17116 17650 17128
rect 17681 17119 17739 17125
rect 17681 17116 17693 17119
rect 17644 17088 17693 17116
rect 17644 17076 17650 17088
rect 17681 17085 17693 17088
rect 17727 17085 17739 17119
rect 17681 17079 17739 17085
rect 17862 17076 17868 17128
rect 17920 17116 17926 17128
rect 18049 17119 18107 17125
rect 18049 17116 18061 17119
rect 17920 17088 18061 17116
rect 17920 17076 17926 17088
rect 18049 17085 18061 17088
rect 18095 17116 18107 17119
rect 18322 17116 18328 17128
rect 18095 17088 18328 17116
rect 18095 17085 18107 17088
rect 18049 17079 18107 17085
rect 18322 17076 18328 17088
rect 18380 17076 18386 17128
rect 18432 17125 18460 17156
rect 18616 17128 18644 17224
rect 18690 17144 18696 17196
rect 18748 17144 18754 17196
rect 19245 17187 19303 17193
rect 19245 17153 19257 17187
rect 19291 17184 19303 17187
rect 19794 17184 19800 17196
rect 19291 17156 19800 17184
rect 19291 17153 19303 17156
rect 19245 17147 19303 17153
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 21744 17184 21772 17224
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 22370 17212 22376 17264
rect 22428 17252 22434 17264
rect 26712 17252 26740 17292
rect 22428 17224 26740 17252
rect 22428 17212 22434 17224
rect 26970 17212 26976 17264
rect 27028 17212 27034 17264
rect 29012 17252 29040 17292
rect 29638 17280 29644 17332
rect 29696 17320 29702 17332
rect 29733 17323 29791 17329
rect 29733 17320 29745 17323
rect 29696 17292 29745 17320
rect 29696 17280 29702 17292
rect 29733 17289 29745 17292
rect 29779 17289 29791 17323
rect 29733 17283 29791 17289
rect 31018 17280 31024 17332
rect 31076 17280 31082 17332
rect 32122 17280 32128 17332
rect 32180 17320 32186 17332
rect 33045 17323 33103 17329
rect 33045 17320 33057 17323
rect 32180 17292 33057 17320
rect 32180 17280 32186 17292
rect 33045 17289 33057 17292
rect 33091 17289 33103 17323
rect 33045 17283 33103 17289
rect 29012 17224 30512 17252
rect 20763 17156 21772 17184
rect 22005 17187 22063 17193
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 22005 17153 22017 17187
rect 22051 17184 22063 17187
rect 22554 17184 22560 17196
rect 22051 17156 22560 17184
rect 22051 17153 22063 17156
rect 22005 17147 22063 17153
rect 22554 17144 22560 17156
rect 22612 17184 22618 17196
rect 23014 17184 23020 17196
rect 22612 17156 23020 17184
rect 22612 17144 22618 17156
rect 23014 17144 23020 17156
rect 23072 17144 23078 17196
rect 23569 17187 23627 17193
rect 23569 17184 23581 17187
rect 23492 17156 23581 17184
rect 18417 17119 18475 17125
rect 18417 17085 18429 17119
rect 18463 17085 18475 17119
rect 18417 17079 18475 17085
rect 18506 17076 18512 17128
rect 18564 17076 18570 17128
rect 18598 17076 18604 17128
rect 18656 17076 18662 17128
rect 18782 17076 18788 17128
rect 18840 17116 18846 17128
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 18840 17088 18981 17116
rect 18840 17076 18846 17088
rect 18969 17085 18981 17088
rect 19015 17085 19027 17119
rect 18969 17079 19027 17085
rect 21085 17119 21143 17125
rect 21085 17085 21097 17119
rect 21131 17116 21143 17119
rect 21266 17116 21272 17128
rect 21131 17088 21272 17116
rect 21131 17085 21143 17088
rect 21085 17079 21143 17085
rect 21266 17076 21272 17088
rect 21324 17076 21330 17128
rect 21358 17076 21364 17128
rect 21416 17116 21422 17128
rect 21821 17119 21879 17125
rect 21821 17116 21833 17119
rect 21416 17088 21833 17116
rect 21416 17076 21422 17088
rect 21821 17085 21833 17088
rect 21867 17085 21879 17119
rect 21821 17079 21879 17085
rect 21913 17119 21971 17125
rect 21913 17085 21925 17119
rect 21959 17116 21971 17119
rect 22186 17116 22192 17128
rect 21959 17088 22192 17116
rect 21959 17085 21971 17088
rect 21913 17079 21971 17085
rect 22186 17076 22192 17088
rect 22244 17076 22250 17128
rect 22278 17076 22284 17128
rect 22336 17116 22342 17128
rect 22373 17119 22431 17125
rect 22373 17116 22385 17119
rect 22336 17088 22385 17116
rect 22336 17076 22342 17088
rect 22373 17085 22385 17088
rect 22419 17085 22431 17119
rect 22373 17079 22431 17085
rect 22925 17119 22983 17125
rect 22925 17085 22937 17119
rect 22971 17116 22983 17119
rect 23492 17116 23520 17156
rect 23569 17153 23581 17156
rect 23615 17153 23627 17187
rect 26053 17187 26111 17193
rect 26053 17184 26065 17187
rect 23569 17147 23627 17153
rect 24412 17156 26065 17184
rect 24412 17128 24440 17156
rect 26053 17153 26065 17156
rect 26099 17153 26111 17187
rect 26053 17147 26111 17153
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17184 28043 17187
rect 28626 17184 28632 17196
rect 28031 17156 28632 17184
rect 28031 17153 28043 17156
rect 27985 17147 28043 17153
rect 28626 17144 28632 17156
rect 28684 17144 28690 17196
rect 29457 17187 29515 17193
rect 29457 17153 29469 17187
rect 29503 17153 29515 17187
rect 29457 17147 29515 17153
rect 22971 17088 23520 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 24302 17076 24308 17128
rect 24360 17076 24366 17128
rect 24394 17076 24400 17128
rect 24452 17076 24458 17128
rect 25130 17076 25136 17128
rect 25188 17076 25194 17128
rect 25866 17076 25872 17128
rect 25924 17076 25930 17128
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17085 27767 17119
rect 29472 17116 29500 17147
rect 29549 17119 29607 17125
rect 29549 17116 29561 17119
rect 29472 17088 29561 17116
rect 27709 17079 27767 17085
rect 29549 17085 29561 17088
rect 29595 17085 29607 17119
rect 29549 17079 29607 17085
rect 15289 17051 15347 17057
rect 15289 17017 15301 17051
rect 15335 17048 15347 17051
rect 15654 17048 15660 17060
rect 15335 17020 15660 17048
rect 15335 17017 15347 17020
rect 15289 17011 15347 17017
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 16022 17008 16028 17060
rect 16080 17008 16086 17060
rect 18524 17048 18552 17076
rect 20993 17051 21051 17057
rect 20993 17048 21005 17051
rect 16132 17020 16514 17048
rect 18340 17020 18552 17048
rect 20470 17020 21005 17048
rect 10367 16952 10824 16980
rect 13173 16983 13231 16989
rect 10367 16949 10379 16952
rect 10321 16943 10379 16949
rect 13173 16949 13185 16983
rect 13219 16949 13231 16983
rect 13173 16943 13231 16949
rect 13906 16940 13912 16992
rect 13964 16940 13970 16992
rect 14182 16940 14188 16992
rect 14240 16940 14246 16992
rect 14921 16983 14979 16989
rect 14921 16949 14933 16983
rect 14967 16980 14979 16983
rect 16132 16980 16160 17020
rect 14967 16952 16160 16980
rect 14967 16949 14979 16952
rect 14921 16943 14979 16949
rect 17494 16940 17500 16992
rect 17552 16940 17558 16992
rect 17957 16983 18015 16989
rect 17957 16949 17969 16983
rect 18003 16980 18015 16983
rect 18138 16980 18144 16992
rect 18003 16952 18144 16980
rect 18003 16949 18015 16952
rect 17957 16943 18015 16949
rect 18138 16940 18144 16952
rect 18196 16940 18202 16992
rect 18340 16989 18368 17020
rect 20993 17017 21005 17020
rect 21039 17017 21051 17051
rect 20993 17011 21051 17017
rect 18325 16983 18383 16989
rect 18325 16949 18337 16983
rect 18371 16949 18383 16983
rect 18325 16943 18383 16949
rect 23750 16940 23756 16992
rect 23808 16940 23814 16992
rect 23842 16940 23848 16992
rect 23900 16980 23906 16992
rect 24489 16983 24547 16989
rect 24489 16980 24501 16983
rect 23900 16952 24501 16980
rect 23900 16940 23906 16952
rect 24489 16949 24501 16952
rect 24535 16949 24547 16983
rect 24489 16943 24547 16949
rect 25225 16983 25283 16989
rect 25225 16949 25237 16983
rect 25271 16980 25283 16983
rect 25590 16980 25596 16992
rect 25271 16952 25596 16980
rect 25271 16949 25283 16952
rect 25225 16943 25283 16949
rect 25590 16940 25596 16952
rect 25648 16940 25654 16992
rect 26326 16940 26332 16992
rect 26384 16980 26390 16992
rect 26697 16983 26755 16989
rect 26697 16980 26709 16983
rect 26384 16952 26709 16980
rect 26384 16940 26390 16952
rect 26697 16949 26709 16952
rect 26743 16949 26755 16983
rect 26697 16943 26755 16949
rect 27614 16940 27620 16992
rect 27672 16980 27678 16992
rect 27724 16980 27752 17079
rect 29730 17076 29736 17128
rect 29788 17116 29794 17128
rect 30377 17119 30435 17125
rect 30377 17116 30389 17119
rect 29788 17088 30389 17116
rect 29788 17076 29794 17088
rect 30377 17085 30389 17088
rect 30423 17085 30435 17119
rect 30484 17116 30512 17224
rect 31036 17184 31064 17280
rect 32677 17187 32735 17193
rect 32677 17184 32689 17187
rect 31036 17156 32689 17184
rect 32677 17153 32689 17156
rect 32723 17153 32735 17187
rect 32677 17147 32735 17153
rect 32950 17144 32956 17196
rect 33008 17144 33014 17196
rect 33594 17144 33600 17196
rect 33652 17144 33658 17196
rect 30484 17088 31340 17116
rect 30377 17079 30435 17085
rect 28994 17008 29000 17060
rect 29052 17008 29058 17060
rect 30392 17048 30420 17079
rect 30392 17020 31248 17048
rect 28902 16980 28908 16992
rect 27672 16952 28908 16980
rect 27672 16940 27678 16952
rect 28902 16940 28908 16952
rect 28960 16940 28966 16992
rect 29454 16940 29460 16992
rect 29512 16980 29518 16992
rect 30558 16980 30564 16992
rect 29512 16952 30564 16980
rect 29512 16940 29518 16952
rect 30558 16940 30564 16952
rect 30616 16940 30622 16992
rect 31220 16989 31248 17020
rect 31312 16992 31340 17088
rect 32030 17008 32036 17060
rect 32088 17008 32094 17060
rect 31205 16983 31263 16989
rect 31205 16949 31217 16983
rect 31251 16949 31263 16983
rect 31205 16943 31263 16949
rect 31294 16940 31300 16992
rect 31352 16940 31358 16992
rect 2760 16890 34316 16912
rect 2760 16838 7210 16890
rect 7262 16838 7274 16890
rect 7326 16838 7338 16890
rect 7390 16838 7402 16890
rect 7454 16838 7466 16890
rect 7518 16838 15099 16890
rect 15151 16838 15163 16890
rect 15215 16838 15227 16890
rect 15279 16838 15291 16890
rect 15343 16838 15355 16890
rect 15407 16838 22988 16890
rect 23040 16838 23052 16890
rect 23104 16838 23116 16890
rect 23168 16838 23180 16890
rect 23232 16838 23244 16890
rect 23296 16838 30877 16890
rect 30929 16838 30941 16890
rect 30993 16838 31005 16890
rect 31057 16838 31069 16890
rect 31121 16838 31133 16890
rect 31185 16838 34316 16890
rect 2760 16816 34316 16838
rect 3881 16779 3939 16785
rect 3881 16745 3893 16779
rect 3927 16745 3939 16779
rect 3881 16739 3939 16745
rect 3789 16643 3847 16649
rect 3789 16609 3801 16643
rect 3835 16640 3847 16643
rect 3896 16640 3924 16739
rect 4522 16736 4528 16788
rect 4580 16776 4586 16788
rect 4709 16779 4767 16785
rect 4709 16776 4721 16779
rect 4580 16748 4721 16776
rect 4580 16736 4586 16748
rect 4709 16745 4721 16748
rect 4755 16745 4767 16779
rect 4709 16739 4767 16745
rect 4798 16736 4804 16788
rect 4856 16736 4862 16788
rect 5258 16736 5264 16788
rect 5316 16736 5322 16788
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 5537 16779 5595 16785
rect 5537 16776 5549 16779
rect 5408 16748 5549 16776
rect 5408 16736 5414 16748
rect 5537 16745 5549 16748
rect 5583 16745 5595 16779
rect 5537 16739 5595 16745
rect 6454 16736 6460 16788
rect 6512 16776 6518 16788
rect 7009 16779 7067 16785
rect 7009 16776 7021 16779
rect 6512 16748 7021 16776
rect 6512 16736 6518 16748
rect 7009 16745 7021 16748
rect 7055 16745 7067 16779
rect 7009 16739 7067 16745
rect 7742 16736 7748 16788
rect 7800 16736 7806 16788
rect 8941 16779 8999 16785
rect 8941 16745 8953 16779
rect 8987 16776 8999 16779
rect 9306 16776 9312 16788
rect 8987 16748 9312 16776
rect 8987 16745 8999 16748
rect 8941 16739 8999 16745
rect 9306 16736 9312 16748
rect 9364 16736 9370 16788
rect 10873 16779 10931 16785
rect 10873 16745 10885 16779
rect 10919 16776 10931 16779
rect 11146 16776 11152 16788
rect 10919 16748 11152 16776
rect 10919 16745 10931 16748
rect 10873 16739 10931 16745
rect 11146 16736 11152 16748
rect 11204 16736 11210 16788
rect 15838 16776 15844 16788
rect 12176 16748 15844 16776
rect 3835 16612 3924 16640
rect 3835 16609 3847 16612
rect 3789 16603 3847 16609
rect 4246 16600 4252 16652
rect 4304 16600 4310 16652
rect 4816 16640 4844 16736
rect 5276 16708 5304 16736
rect 12176 16720 12204 16748
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 15930 16736 15936 16788
rect 15988 16736 15994 16788
rect 16114 16736 16120 16788
rect 16172 16736 16178 16788
rect 16301 16779 16359 16785
rect 16301 16745 16313 16779
rect 16347 16776 16359 16779
rect 16574 16776 16580 16788
rect 16347 16748 16580 16776
rect 16347 16745 16359 16748
rect 16301 16739 16359 16745
rect 16574 16736 16580 16748
rect 16632 16736 16638 16788
rect 18598 16776 18604 16788
rect 18064 16748 18604 16776
rect 9953 16711 10011 16717
rect 9953 16708 9965 16711
rect 5276 16680 5488 16708
rect 5460 16649 5488 16680
rect 6104 16680 9965 16708
rect 6104 16652 6132 16680
rect 9953 16677 9965 16680
rect 9999 16708 10011 16711
rect 11054 16708 11060 16720
rect 9999 16680 11060 16708
rect 9999 16677 10011 16680
rect 9953 16671 10011 16677
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 11974 16668 11980 16720
rect 12032 16668 12038 16720
rect 12158 16668 12164 16720
rect 12216 16668 12222 16720
rect 13998 16668 14004 16720
rect 14056 16668 14062 16720
rect 15473 16711 15531 16717
rect 15473 16677 15485 16711
rect 15519 16708 15531 16711
rect 15562 16708 15568 16720
rect 15519 16680 15568 16708
rect 15519 16677 15531 16680
rect 15473 16671 15531 16677
rect 5261 16643 5319 16649
rect 5261 16640 5273 16643
rect 4816 16612 5273 16640
rect 5261 16609 5273 16612
rect 5307 16609 5319 16643
rect 5261 16603 5319 16609
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16609 5503 16643
rect 5445 16603 5503 16609
rect 5721 16643 5779 16649
rect 5721 16609 5733 16643
rect 5767 16640 5779 16643
rect 6086 16640 6092 16652
rect 5767 16612 6092 16640
rect 5767 16609 5779 16612
rect 5721 16603 5779 16609
rect 6086 16600 6092 16612
rect 6144 16600 6150 16652
rect 7653 16643 7711 16649
rect 7653 16609 7665 16643
rect 7699 16640 7711 16643
rect 8202 16640 8208 16652
rect 7699 16612 8208 16640
rect 7699 16609 7711 16612
rect 7653 16603 7711 16609
rect 8202 16600 8208 16612
rect 8260 16600 8266 16652
rect 8478 16600 8484 16652
rect 8536 16600 8542 16652
rect 8573 16643 8631 16649
rect 8573 16609 8585 16643
rect 8619 16609 8631 16643
rect 8573 16603 8631 16609
rect 4338 16532 4344 16584
rect 4396 16532 4402 16584
rect 4522 16532 4528 16584
rect 4580 16532 4586 16584
rect 8294 16532 8300 16584
rect 8352 16532 8358 16584
rect 8588 16572 8616 16603
rect 8662 16600 8668 16652
rect 8720 16640 8726 16652
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8720 16612 9045 16640
rect 8720 16600 8726 16612
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9033 16603 9091 16609
rect 9140 16612 9689 16640
rect 9140 16584 9168 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16640 10379 16643
rect 12713 16643 12771 16649
rect 10367 16612 11008 16640
rect 10367 16609 10379 16612
rect 10321 16603 10379 16609
rect 9122 16572 9128 16584
rect 8588 16544 9128 16572
rect 9122 16532 9128 16544
rect 9180 16532 9186 16584
rect 10980 16581 11008 16612
rect 12713 16609 12725 16643
rect 12759 16640 12771 16643
rect 13078 16640 13084 16652
rect 12759 16612 13084 16640
rect 12759 16609 12771 16612
rect 12713 16603 12771 16609
rect 13078 16600 13084 16612
rect 13136 16640 13142 16652
rect 13173 16643 13231 16649
rect 13173 16640 13185 16643
rect 13136 16612 13185 16640
rect 13136 16600 13142 16612
rect 13173 16609 13185 16612
rect 13219 16609 13231 16643
rect 13173 16603 13231 16609
rect 10965 16575 11023 16581
rect 10965 16541 10977 16575
rect 11011 16541 11023 16575
rect 10965 16535 11023 16541
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16572 12495 16575
rect 12483 16544 13124 16572
rect 12483 16541 12495 16544
rect 12437 16535 12495 16541
rect 13096 16504 13124 16544
rect 13446 16532 13452 16584
rect 13504 16532 13510 16584
rect 13538 16532 13544 16584
rect 13596 16572 13602 16584
rect 15488 16572 15516 16671
rect 15562 16668 15568 16680
rect 15620 16708 15626 16720
rect 16132 16708 16160 16736
rect 15620 16680 16160 16708
rect 15620 16668 15626 16680
rect 16482 16668 16488 16720
rect 16540 16708 16546 16720
rect 18064 16708 18092 16748
rect 18598 16736 18604 16748
rect 18656 16736 18662 16788
rect 21634 16776 21640 16788
rect 20180 16748 21640 16776
rect 20180 16717 20208 16748
rect 21634 16736 21640 16748
rect 21692 16736 21698 16788
rect 22370 16736 22376 16788
rect 22428 16736 22434 16788
rect 22830 16736 22836 16788
rect 22888 16736 22894 16788
rect 22925 16779 22983 16785
rect 22925 16745 22937 16779
rect 22971 16776 22983 16779
rect 23842 16776 23848 16788
rect 22971 16748 23848 16776
rect 22971 16745 22983 16748
rect 22925 16739 22983 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 23937 16779 23995 16785
rect 23937 16745 23949 16779
rect 23983 16776 23995 16779
rect 24210 16776 24216 16788
rect 23983 16748 24216 16776
rect 23983 16745 23995 16748
rect 23937 16739 23995 16745
rect 24210 16736 24216 16748
rect 24268 16736 24274 16788
rect 24302 16736 24308 16788
rect 24360 16736 24366 16788
rect 25866 16736 25872 16788
rect 25924 16776 25930 16788
rect 26053 16779 26111 16785
rect 26053 16776 26065 16779
rect 25924 16748 26065 16776
rect 25924 16736 25930 16748
rect 26053 16745 26065 16748
rect 26099 16745 26111 16779
rect 28166 16776 28172 16788
rect 26053 16739 26111 16745
rect 28092 16748 28172 16776
rect 16540 16680 18092 16708
rect 18141 16711 18199 16717
rect 16540 16668 16546 16680
rect 18141 16677 18153 16711
rect 18187 16708 18199 16711
rect 20165 16711 20223 16717
rect 20165 16708 20177 16711
rect 18187 16680 20177 16708
rect 18187 16677 18199 16680
rect 18141 16671 18199 16677
rect 20165 16677 20177 16680
rect 20211 16677 20223 16711
rect 20806 16708 20812 16720
rect 20165 16671 20223 16677
rect 20640 16680 20812 16708
rect 15841 16643 15899 16649
rect 15841 16609 15853 16643
rect 15887 16640 15899 16643
rect 15887 16612 16804 16640
rect 15887 16609 15899 16612
rect 15841 16603 15899 16609
rect 16776 16584 16804 16612
rect 16942 16600 16948 16652
rect 17000 16600 17006 16652
rect 17586 16600 17592 16652
rect 17644 16600 17650 16652
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 20640 16649 20668 16680
rect 20806 16668 20812 16680
rect 20864 16668 20870 16720
rect 24320 16708 24348 16736
rect 23216 16680 24348 16708
rect 20441 16643 20499 16649
rect 20441 16640 20453 16643
rect 19392 16612 20453 16640
rect 19392 16600 19398 16612
rect 20441 16609 20453 16612
rect 20487 16609 20499 16643
rect 20441 16603 20499 16609
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16609 20683 16643
rect 20625 16603 20683 16609
rect 22002 16600 22008 16652
rect 22060 16600 22066 16652
rect 23216 16630 23244 16680
rect 25038 16668 25044 16720
rect 25096 16668 25102 16720
rect 25976 16680 27660 16708
rect 23216 16602 23336 16630
rect 13596 16544 15516 16572
rect 13596 16532 13602 16544
rect 15654 16532 15660 16584
rect 15712 16532 15718 16584
rect 16758 16532 16764 16584
rect 16816 16532 16822 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20732 16544 20913 16572
rect 13170 16504 13176 16516
rect 13096 16476 13176 16504
rect 13170 16464 13176 16476
rect 13228 16464 13234 16516
rect 14844 16476 16896 16504
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16436 3203 16439
rect 3234 16436 3240 16448
rect 3191 16408 3240 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 3234 16396 3240 16408
rect 3292 16396 3298 16448
rect 7926 16396 7932 16448
rect 7984 16436 7990 16448
rect 14844 16436 14872 16476
rect 7984 16408 14872 16436
rect 7984 16396 7990 16408
rect 14918 16396 14924 16448
rect 14976 16396 14982 16448
rect 16482 16396 16488 16448
rect 16540 16436 16546 16448
rect 16761 16439 16819 16445
rect 16761 16436 16773 16439
rect 16540 16408 16773 16436
rect 16540 16396 16546 16408
rect 16761 16405 16773 16408
rect 16807 16405 16819 16439
rect 16868 16436 16896 16476
rect 20732 16448 20760 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 22741 16575 22799 16581
rect 22741 16541 22753 16575
rect 22787 16572 22799 16575
rect 22787 16544 23244 16572
rect 22787 16541 22799 16544
rect 22741 16535 22799 16541
rect 18138 16436 18144 16448
rect 16868 16408 18144 16436
rect 16761 16399 16819 16405
rect 18138 16396 18144 16408
rect 18196 16396 18202 16448
rect 18414 16396 18420 16448
rect 18472 16436 18478 16448
rect 18693 16439 18751 16445
rect 18693 16436 18705 16439
rect 18472 16408 18705 16436
rect 18472 16396 18478 16408
rect 18693 16405 18705 16408
rect 18739 16436 18751 16439
rect 18782 16436 18788 16448
rect 18739 16408 18788 16436
rect 18739 16405 18751 16408
rect 18693 16399 18751 16405
rect 18782 16396 18788 16408
rect 18840 16396 18846 16448
rect 20346 16396 20352 16448
rect 20404 16396 20410 16448
rect 20714 16396 20720 16448
rect 20772 16396 20778 16448
rect 22554 16396 22560 16448
rect 22612 16436 22618 16448
rect 22830 16436 22836 16448
rect 22612 16408 22836 16436
rect 22612 16396 22618 16408
rect 22830 16396 22836 16408
rect 22888 16396 22894 16448
rect 23216 16436 23244 16544
rect 23308 16513 23336 16602
rect 23474 16600 23480 16652
rect 23532 16640 23538 16652
rect 23842 16640 23848 16652
rect 23532 16612 23848 16640
rect 23532 16600 23538 16612
rect 23842 16600 23848 16612
rect 23900 16600 23906 16652
rect 24167 16643 24225 16649
rect 24167 16640 24179 16643
rect 23952 16612 24179 16640
rect 23382 16532 23388 16584
rect 23440 16572 23446 16584
rect 23952 16572 23980 16612
rect 24167 16609 24179 16612
rect 24213 16640 24225 16643
rect 24394 16640 24400 16652
rect 24213 16612 24400 16640
rect 24213 16609 24225 16612
rect 24167 16603 24225 16609
rect 24394 16600 24400 16612
rect 24452 16600 24458 16652
rect 25590 16600 25596 16652
rect 25648 16600 25654 16652
rect 25976 16649 26004 16680
rect 27632 16652 27660 16680
rect 25961 16643 26019 16649
rect 25961 16609 25973 16643
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 26237 16643 26295 16649
rect 26237 16609 26249 16643
rect 26283 16609 26295 16643
rect 26237 16603 26295 16609
rect 23440 16544 23980 16572
rect 26252 16572 26280 16603
rect 26326 16600 26332 16652
rect 26384 16600 26390 16652
rect 26418 16600 26424 16652
rect 26476 16600 26482 16652
rect 26510 16600 26516 16652
rect 26568 16600 26574 16652
rect 26602 16600 26608 16652
rect 26660 16600 26666 16652
rect 27065 16643 27123 16649
rect 27065 16609 27077 16643
rect 27111 16609 27123 16643
rect 27065 16603 27123 16609
rect 27157 16643 27215 16649
rect 27157 16609 27169 16643
rect 27203 16640 27215 16643
rect 27522 16640 27528 16652
rect 27203 16612 27528 16640
rect 27203 16609 27215 16612
rect 27157 16603 27215 16609
rect 26528 16572 26556 16600
rect 26252 16544 26556 16572
rect 27080 16572 27108 16603
rect 27522 16600 27528 16612
rect 27580 16600 27586 16652
rect 27614 16600 27620 16652
rect 27672 16600 27678 16652
rect 27706 16600 27712 16652
rect 27764 16600 27770 16652
rect 27801 16643 27859 16649
rect 27801 16609 27813 16643
rect 27847 16640 27859 16643
rect 28092 16640 28120 16748
rect 28166 16736 28172 16748
rect 28224 16736 28230 16788
rect 28350 16736 28356 16788
rect 28408 16776 28414 16788
rect 28813 16779 28871 16785
rect 28813 16776 28825 16779
rect 28408 16748 28825 16776
rect 28408 16736 28414 16748
rect 28813 16745 28825 16748
rect 28859 16745 28871 16779
rect 28813 16739 28871 16745
rect 29546 16736 29552 16788
rect 29604 16736 29610 16788
rect 29730 16736 29736 16788
rect 29788 16736 29794 16788
rect 29822 16736 29828 16788
rect 29880 16736 29886 16788
rect 29917 16779 29975 16785
rect 29917 16745 29929 16779
rect 29963 16776 29975 16779
rect 30098 16776 30104 16788
rect 29963 16748 30104 16776
rect 29963 16745 29975 16748
rect 29917 16739 29975 16745
rect 30098 16736 30104 16748
rect 30156 16776 30162 16788
rect 30351 16779 30409 16785
rect 30351 16776 30363 16779
rect 30156 16748 30363 16776
rect 30156 16736 30162 16748
rect 30351 16745 30363 16748
rect 30397 16745 30409 16779
rect 30351 16739 30409 16745
rect 30650 16736 30656 16788
rect 30708 16776 30714 16788
rect 30751 16779 30809 16785
rect 30751 16776 30763 16779
rect 30708 16748 30763 16776
rect 30708 16736 30714 16748
rect 30751 16745 30763 16748
rect 30797 16745 30809 16779
rect 30751 16739 30809 16745
rect 31294 16736 31300 16788
rect 31352 16776 31358 16788
rect 31352 16748 32260 16776
rect 31352 16736 31358 16748
rect 29564 16708 29592 16736
rect 30190 16708 30196 16720
rect 28184 16680 29592 16708
rect 29656 16680 30196 16708
rect 28184 16649 28212 16680
rect 27847 16612 28120 16640
rect 28169 16643 28227 16649
rect 27847 16609 27859 16612
rect 27801 16603 27859 16609
rect 28169 16609 28181 16643
rect 28215 16609 28227 16643
rect 28169 16603 28227 16609
rect 28353 16643 28411 16649
rect 28353 16609 28365 16643
rect 28399 16640 28411 16643
rect 28399 16612 28672 16640
rect 28399 16609 28411 16612
rect 28353 16603 28411 16609
rect 27724 16572 27752 16600
rect 27080 16544 27752 16572
rect 28445 16575 28503 16581
rect 23440 16532 23446 16544
rect 23293 16507 23351 16513
rect 23293 16473 23305 16507
rect 23339 16473 23351 16507
rect 23293 16467 23351 16473
rect 23566 16464 23572 16516
rect 23624 16464 23630 16516
rect 26326 16464 26332 16516
rect 26384 16504 26390 16516
rect 27080 16504 27108 16544
rect 28445 16541 28457 16575
rect 28491 16572 28503 16575
rect 28534 16572 28540 16584
rect 28491 16544 28540 16572
rect 28491 16541 28503 16544
rect 28445 16535 28503 16541
rect 28534 16532 28540 16544
rect 28592 16532 28598 16584
rect 28644 16572 28672 16612
rect 28718 16600 28724 16652
rect 28776 16600 28782 16652
rect 29656 16640 29684 16680
rect 30190 16668 30196 16680
rect 30248 16668 30254 16720
rect 30558 16668 30564 16720
rect 30616 16708 30622 16720
rect 31849 16711 31907 16717
rect 31849 16708 31861 16711
rect 30616 16680 31616 16708
rect 30616 16668 30622 16680
rect 28828 16612 29684 16640
rect 28828 16572 28856 16612
rect 29730 16600 29736 16652
rect 29788 16600 29794 16652
rect 29914 16600 29920 16652
rect 29972 16640 29978 16652
rect 30101 16643 30159 16649
rect 30101 16640 30113 16643
rect 29972 16612 30113 16640
rect 29972 16600 29978 16612
rect 30101 16609 30113 16612
rect 30147 16609 30159 16643
rect 30208 16640 30236 16668
rect 30653 16643 30711 16649
rect 30653 16640 30665 16643
rect 30208 16612 30665 16640
rect 30101 16603 30159 16609
rect 30653 16609 30665 16612
rect 30699 16609 30711 16643
rect 30653 16603 30711 16609
rect 30742 16600 30748 16652
rect 30800 16640 30806 16652
rect 30837 16643 30895 16649
rect 30837 16640 30849 16643
rect 30800 16612 30849 16640
rect 30800 16600 30806 16612
rect 30837 16609 30849 16612
rect 30883 16609 30895 16643
rect 30837 16603 30895 16609
rect 30929 16643 30987 16649
rect 30929 16609 30941 16643
rect 30975 16640 30987 16643
rect 31021 16643 31079 16649
rect 31021 16640 31033 16643
rect 30975 16612 31033 16640
rect 30975 16609 30987 16612
rect 30929 16603 30987 16609
rect 31021 16609 31033 16612
rect 31067 16609 31079 16643
rect 31021 16603 31079 16609
rect 28644 16544 28856 16572
rect 29178 16532 29184 16584
rect 29236 16532 29242 16584
rect 29549 16575 29607 16581
rect 29549 16541 29561 16575
rect 29595 16572 29607 16575
rect 29748 16572 29776 16600
rect 30466 16572 30472 16584
rect 29595 16544 29776 16572
rect 29840 16544 30472 16572
rect 29595 16541 29607 16544
rect 29549 16535 29607 16541
rect 26384 16476 27108 16504
rect 27801 16507 27859 16513
rect 26384 16464 26390 16476
rect 27801 16473 27813 16507
rect 27847 16504 27859 16507
rect 27890 16504 27896 16516
rect 27847 16476 27896 16504
rect 27847 16473 27859 16476
rect 27801 16467 27859 16473
rect 27890 16464 27896 16476
rect 27948 16464 27954 16516
rect 27985 16507 28043 16513
rect 27985 16473 27997 16507
rect 28031 16504 28043 16507
rect 29196 16504 29224 16532
rect 28031 16476 29224 16504
rect 28031 16473 28043 16476
rect 27985 16467 28043 16473
rect 29638 16464 29644 16516
rect 29696 16504 29702 16516
rect 29840 16504 29868 16544
rect 30466 16532 30472 16544
rect 30524 16532 30530 16584
rect 31588 16572 31616 16680
rect 31680 16680 31861 16708
rect 31680 16649 31708 16680
rect 31849 16677 31861 16680
rect 31895 16677 31907 16711
rect 31849 16671 31907 16677
rect 32232 16649 32260 16748
rect 31665 16643 31723 16649
rect 31665 16609 31677 16643
rect 31711 16609 31723 16643
rect 31665 16603 31723 16609
rect 31757 16643 31815 16649
rect 31757 16609 31769 16643
rect 31803 16609 31815 16643
rect 31757 16603 31815 16609
rect 31941 16643 31999 16649
rect 31941 16609 31953 16643
rect 31987 16609 31999 16643
rect 31941 16603 31999 16609
rect 32217 16643 32275 16649
rect 32217 16609 32229 16643
rect 32263 16609 32275 16643
rect 32217 16603 32275 16609
rect 31772 16572 31800 16603
rect 31588 16544 31800 16572
rect 29696 16476 29868 16504
rect 29696 16464 29702 16476
rect 30190 16464 30196 16516
rect 30248 16464 30254 16516
rect 30484 16504 30512 16532
rect 31956 16504 31984 16603
rect 33042 16532 33048 16584
rect 33100 16532 33106 16584
rect 30484 16476 31984 16504
rect 23584 16436 23612 16464
rect 23216 16408 23612 16436
rect 28718 16396 28724 16448
rect 28776 16436 28782 16448
rect 29822 16436 29828 16448
rect 28776 16408 29828 16436
rect 28776 16396 28782 16408
rect 29822 16396 29828 16408
rect 29880 16436 29886 16448
rect 30377 16439 30435 16445
rect 30377 16436 30389 16439
rect 29880 16408 30389 16436
rect 29880 16396 29886 16408
rect 30377 16405 30389 16408
rect 30423 16405 30435 16439
rect 30377 16399 30435 16405
rect 2760 16346 34316 16368
rect 2760 16294 6550 16346
rect 6602 16294 6614 16346
rect 6666 16294 6678 16346
rect 6730 16294 6742 16346
rect 6794 16294 6806 16346
rect 6858 16294 14439 16346
rect 14491 16294 14503 16346
rect 14555 16294 14567 16346
rect 14619 16294 14631 16346
rect 14683 16294 14695 16346
rect 14747 16294 22328 16346
rect 22380 16294 22392 16346
rect 22444 16294 22456 16346
rect 22508 16294 22520 16346
rect 22572 16294 22584 16346
rect 22636 16294 30217 16346
rect 30269 16294 30281 16346
rect 30333 16294 30345 16346
rect 30397 16294 30409 16346
rect 30461 16294 30473 16346
rect 30525 16294 34316 16346
rect 2760 16272 34316 16294
rect 4338 16192 4344 16244
rect 4396 16232 4402 16244
rect 4801 16235 4859 16241
rect 4801 16232 4813 16235
rect 4396 16204 4813 16232
rect 4396 16192 4402 16204
rect 4801 16201 4813 16204
rect 4847 16201 4859 16235
rect 4801 16195 4859 16201
rect 6362 16192 6368 16244
rect 6420 16232 6426 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 6420 16204 8217 16232
rect 6420 16192 6426 16204
rect 8205 16201 8217 16204
rect 8251 16232 8263 16235
rect 8251 16204 12434 16232
rect 8251 16201 8263 16204
rect 8205 16195 8263 16201
rect 11054 16124 11060 16176
rect 11112 16124 11118 16176
rect 12406 16164 12434 16204
rect 13170 16192 13176 16244
rect 13228 16192 13234 16244
rect 13998 16192 14004 16244
rect 14056 16192 14062 16244
rect 16022 16192 16028 16244
rect 16080 16192 16086 16244
rect 16758 16192 16764 16244
rect 16816 16232 16822 16244
rect 17678 16232 17684 16244
rect 16816 16204 17684 16232
rect 16816 16192 16822 16204
rect 17678 16192 17684 16204
rect 17736 16192 17742 16244
rect 23566 16192 23572 16244
rect 23624 16232 23630 16244
rect 24578 16232 24584 16244
rect 23624 16204 24584 16232
rect 23624 16192 23630 16204
rect 24578 16192 24584 16204
rect 24636 16232 24642 16244
rect 24636 16204 25004 16232
rect 24636 16192 24642 16204
rect 14553 16167 14611 16173
rect 14553 16164 14565 16167
rect 12406 16136 14565 16164
rect 14553 16133 14565 16136
rect 14599 16164 14611 16167
rect 15654 16164 15660 16176
rect 14599 16136 15660 16164
rect 14599 16133 14611 16136
rect 14553 16127 14611 16133
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 20717 16167 20775 16173
rect 20717 16133 20729 16167
rect 20763 16164 20775 16167
rect 20806 16164 20812 16176
rect 20763 16136 20812 16164
rect 20763 16133 20775 16136
rect 20717 16127 20775 16133
rect 20806 16124 20812 16136
rect 20864 16124 20870 16176
rect 4062 16096 4068 16108
rect 3068 16068 4068 16096
rect 3068 16040 3096 16068
rect 4062 16056 4068 16068
rect 4120 16056 4126 16108
rect 5258 16096 5264 16108
rect 5092 16068 5264 16096
rect 3050 15988 3056 16040
rect 3108 15988 3114 16040
rect 5092 16037 5120 16068
rect 5258 16056 5264 16068
rect 5316 16056 5322 16108
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 6512 16068 7205 16096
rect 6512 16056 6518 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 11072 16096 11100 16124
rect 11072 16068 11376 16096
rect 7193 16059 7251 16065
rect 11348 16040 11376 16068
rect 13078 16056 13084 16108
rect 13136 16056 13142 16108
rect 13814 16056 13820 16108
rect 13872 16056 13878 16108
rect 15013 16099 15071 16105
rect 15013 16065 15025 16099
rect 15059 16096 15071 16099
rect 15059 16068 16344 16096
rect 15059 16065 15071 16068
rect 15013 16059 15071 16065
rect 5077 16031 5135 16037
rect 5077 15997 5089 16031
rect 5123 15997 5135 16031
rect 5077 15991 5135 15997
rect 7926 15988 7932 16040
rect 7984 15988 7990 16040
rect 10413 16031 10471 16037
rect 10413 15997 10425 16031
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 3234 15920 3240 15972
rect 3292 15960 3298 15972
rect 3329 15963 3387 15969
rect 3329 15960 3341 15963
rect 3292 15932 3341 15960
rect 3292 15920 3298 15932
rect 3329 15929 3341 15932
rect 3375 15929 3387 15963
rect 4985 15963 5043 15969
rect 4985 15960 4997 15963
rect 4554 15932 4997 15960
rect 3329 15923 3387 15929
rect 4985 15929 4997 15932
rect 5031 15929 5043 15963
rect 4985 15923 5043 15929
rect 5902 15920 5908 15972
rect 5960 15920 5966 15972
rect 6914 15920 6920 15972
rect 6972 15920 6978 15972
rect 9674 15920 9680 15972
rect 9732 15920 9738 15972
rect 10134 15920 10140 15972
rect 10192 15920 10198 15972
rect 10428 15960 10456 15991
rect 10502 15988 10508 16040
rect 10560 16028 10566 16040
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10560 16000 11161 16028
rect 10560 15988 10566 16000
rect 11149 15997 11161 16000
rect 11195 15997 11207 16031
rect 11149 15991 11207 15997
rect 11330 15988 11336 16040
rect 11388 15988 11394 16040
rect 13096 15960 13124 16056
rect 13906 15988 13912 16040
rect 13964 15988 13970 16040
rect 10244 15932 11284 15960
rect 10244 15904 10272 15932
rect 5442 15852 5448 15904
rect 5500 15852 5506 15904
rect 5626 15852 5632 15904
rect 5684 15892 5690 15904
rect 6270 15892 6276 15904
rect 5684 15864 6276 15892
rect 5684 15852 5690 15864
rect 6270 15852 6276 15864
rect 6328 15892 6334 15904
rect 7285 15895 7343 15901
rect 7285 15892 7297 15895
rect 6328 15864 7297 15892
rect 6328 15852 6334 15864
rect 7285 15861 7297 15864
rect 7331 15861 7343 15895
rect 7285 15855 7343 15861
rect 8665 15895 8723 15901
rect 8665 15861 8677 15895
rect 8711 15892 8723 15895
rect 9766 15892 9772 15904
rect 8711 15864 9772 15892
rect 8711 15861 8723 15864
rect 8665 15855 8723 15861
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 10226 15852 10232 15904
rect 10284 15852 10290 15904
rect 10594 15852 10600 15904
rect 10652 15852 10658 15904
rect 11256 15892 11284 15932
rect 12406 15932 13124 15960
rect 12406 15892 12434 15932
rect 13170 15920 13176 15972
rect 13228 15960 13234 15972
rect 13924 15960 13952 15988
rect 13228 15932 13952 15960
rect 13228 15920 13234 15932
rect 11256 15864 12434 15892
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 15028 15892 15056 16059
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 16028 15163 16031
rect 16316 16028 16344 16068
rect 16574 16056 16580 16108
rect 16632 16056 16638 16108
rect 17405 16099 17463 16105
rect 17405 16065 17417 16099
rect 17451 16096 17463 16099
rect 17494 16096 17500 16108
rect 17451 16068 17500 16096
rect 17451 16065 17463 16068
rect 17405 16059 17463 16065
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 17681 16099 17739 16105
rect 17681 16065 17693 16099
rect 17727 16096 17739 16099
rect 18414 16096 18420 16108
rect 17727 16068 18420 16096
rect 17727 16065 17739 16068
rect 17681 16059 17739 16065
rect 18414 16056 18420 16068
rect 18472 16056 18478 16108
rect 21910 16056 21916 16108
rect 21968 16096 21974 16108
rect 22741 16099 22799 16105
rect 22741 16096 22753 16099
rect 21968 16068 22753 16096
rect 21968 16056 21974 16068
rect 22741 16065 22753 16068
rect 22787 16065 22799 16099
rect 22741 16059 22799 16065
rect 23017 16099 23075 16105
rect 23017 16065 23029 16099
rect 23063 16096 23075 16099
rect 23750 16096 23756 16108
rect 23063 16068 23756 16096
rect 23063 16065 23075 16068
rect 23017 16059 23075 16065
rect 23750 16056 23756 16068
rect 23808 16056 23814 16108
rect 24976 16096 25004 16204
rect 25038 16192 25044 16244
rect 25096 16232 25102 16244
rect 25133 16235 25191 16241
rect 25133 16232 25145 16235
rect 25096 16204 25145 16232
rect 25096 16192 25102 16204
rect 25133 16201 25145 16204
rect 25179 16201 25191 16235
rect 25133 16195 25191 16201
rect 28813 16235 28871 16241
rect 28813 16201 28825 16235
rect 28859 16232 28871 16235
rect 28902 16232 28908 16244
rect 28859 16204 28908 16232
rect 28859 16201 28871 16204
rect 28813 16195 28871 16201
rect 28902 16192 28908 16204
rect 28960 16192 28966 16244
rect 29457 16235 29515 16241
rect 29457 16201 29469 16235
rect 29503 16232 29515 16235
rect 29914 16232 29920 16244
rect 29503 16204 29920 16232
rect 29503 16201 29515 16204
rect 29457 16195 29515 16201
rect 29914 16192 29920 16204
rect 29972 16192 29978 16244
rect 32030 16192 32036 16244
rect 32088 16192 32094 16244
rect 26050 16124 26056 16176
rect 26108 16164 26114 16176
rect 26421 16167 26479 16173
rect 26421 16164 26433 16167
rect 26108 16136 26433 16164
rect 26108 16124 26114 16136
rect 26421 16133 26433 16136
rect 26467 16164 26479 16167
rect 28442 16164 28448 16176
rect 26467 16136 28448 16164
rect 26467 16133 26479 16136
rect 26421 16127 26479 16133
rect 28442 16124 28448 16136
rect 28500 16164 28506 16176
rect 29733 16167 29791 16173
rect 28500 16136 28994 16164
rect 28500 16124 28506 16136
rect 26513 16099 26571 16105
rect 26513 16096 26525 16099
rect 24976 16068 26525 16096
rect 26513 16065 26525 16068
rect 26559 16096 26571 16099
rect 28966 16096 28994 16136
rect 29733 16133 29745 16167
rect 29779 16164 29791 16167
rect 29779 16136 30236 16164
rect 29779 16133 29791 16136
rect 29733 16127 29791 16133
rect 29638 16096 29644 16108
rect 26559 16068 27200 16096
rect 26559 16065 26571 16068
rect 26513 16059 26571 16065
rect 17034 16028 17040 16040
rect 15151 16000 16252 16028
rect 16316 16000 17040 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 16224 15904 16252 16000
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 19242 15988 19248 16040
rect 19300 16028 19306 16040
rect 19613 16031 19671 16037
rect 19613 16028 19625 16031
rect 19300 16000 19625 16028
rect 19300 15988 19306 16000
rect 19613 15997 19625 16000
rect 19659 15997 19671 16031
rect 19613 15991 19671 15997
rect 19794 15988 19800 16040
rect 19852 16028 19858 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19852 16000 19901 16028
rect 19852 15988 19858 16000
rect 19889 15997 19901 16000
rect 19935 15997 19947 16031
rect 19889 15991 19947 15997
rect 20346 15988 20352 16040
rect 20404 15988 20410 16040
rect 20438 15988 20444 16040
rect 20496 16028 20502 16040
rect 20533 16031 20591 16037
rect 20533 16028 20545 16031
rect 20496 16000 20545 16028
rect 20496 15988 20502 16000
rect 20533 15997 20545 16000
rect 20579 15997 20591 16031
rect 20533 15991 20591 15997
rect 20717 16031 20775 16037
rect 20717 15997 20729 16031
rect 20763 15997 20775 16031
rect 20717 15991 20775 15997
rect 16758 15920 16764 15972
rect 16816 15960 16822 15972
rect 17957 15963 18015 15969
rect 17957 15960 17969 15963
rect 16816 15932 17969 15960
rect 16816 15920 16822 15932
rect 17957 15929 17969 15932
rect 18003 15929 18015 15963
rect 20364 15960 20392 15988
rect 19182 15932 20392 15960
rect 17957 15923 18015 15929
rect 13044 15864 15056 15892
rect 15197 15895 15255 15901
rect 13044 15852 13050 15864
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15470 15892 15476 15904
rect 15243 15864 15476 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16206 15852 16212 15904
rect 16264 15852 16270 15904
rect 19426 15852 19432 15904
rect 19484 15852 19490 15904
rect 19886 15852 19892 15904
rect 19944 15892 19950 15904
rect 20732 15892 20760 15991
rect 20898 15988 20904 16040
rect 20956 15988 20962 16040
rect 24946 15988 24952 16040
rect 25004 16028 25010 16040
rect 25225 16031 25283 16037
rect 25225 16028 25237 16031
rect 25004 16000 25237 16028
rect 25004 15988 25010 16000
rect 25225 15997 25237 16000
rect 25271 15997 25283 16031
rect 26694 16028 26700 16040
rect 25225 15991 25283 15997
rect 26068 16000 26700 16028
rect 23750 15920 23756 15972
rect 23808 15920 23814 15972
rect 24394 15920 24400 15972
rect 24452 15960 24458 15972
rect 26068 15969 26096 16000
rect 26694 15988 26700 16000
rect 26752 15988 26758 16040
rect 26053 15963 26111 15969
rect 26053 15960 26065 15963
rect 24452 15932 26065 15960
rect 24452 15920 24458 15932
rect 26053 15929 26065 15932
rect 26099 15929 26111 15963
rect 26053 15923 26111 15929
rect 26237 15963 26295 15969
rect 26237 15929 26249 15963
rect 26283 15960 26295 15963
rect 26326 15960 26332 15972
rect 26283 15932 26332 15960
rect 26283 15929 26295 15932
rect 26237 15923 26295 15929
rect 26326 15920 26332 15932
rect 26384 15920 26390 15972
rect 27172 15960 27200 16068
rect 27264 16068 28764 16096
rect 28966 16068 29644 16096
rect 27264 16037 27292 16068
rect 28736 16040 28764 16068
rect 29638 16056 29644 16068
rect 29696 16056 29702 16108
rect 29914 16056 29920 16108
rect 29972 16056 29978 16108
rect 30208 16105 30236 16136
rect 30193 16099 30251 16105
rect 30193 16065 30205 16099
rect 30239 16065 30251 16099
rect 33134 16096 33140 16108
rect 30193 16059 30251 16065
rect 32140 16068 33140 16096
rect 27249 16031 27307 16037
rect 27249 15997 27261 16031
rect 27295 15997 27307 16031
rect 27249 15991 27307 15997
rect 27338 15988 27344 16040
rect 27396 15988 27402 16040
rect 28718 15988 28724 16040
rect 28776 15988 28782 16040
rect 28810 15988 28816 16040
rect 28868 16028 28874 16040
rect 29365 16031 29423 16037
rect 29365 16028 29377 16031
rect 28868 16000 29377 16028
rect 28868 15988 28874 16000
rect 29365 15997 29377 16000
rect 29411 16028 29423 16031
rect 29932 16028 29960 16056
rect 30009 16031 30067 16037
rect 30009 16028 30021 16031
rect 29411 16000 29868 16028
rect 29932 16000 30021 16028
rect 29411 15997 29423 16000
rect 29365 15991 29423 15997
rect 29641 15963 29699 15969
rect 27172 15932 28994 15960
rect 21174 15892 21180 15904
rect 19944 15864 21180 15892
rect 19944 15852 19950 15864
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 21450 15852 21456 15904
rect 21508 15892 21514 15904
rect 21634 15892 21640 15904
rect 21508 15864 21640 15892
rect 21508 15852 21514 15864
rect 21634 15852 21640 15864
rect 21692 15892 21698 15904
rect 22189 15895 22247 15901
rect 22189 15892 22201 15895
rect 21692 15864 22201 15892
rect 21692 15852 21698 15864
rect 22189 15861 22201 15864
rect 22235 15892 22247 15895
rect 24026 15892 24032 15904
rect 22235 15864 24032 15892
rect 22235 15861 22247 15864
rect 22189 15855 22247 15861
rect 24026 15852 24032 15864
rect 24084 15852 24090 15904
rect 24489 15895 24547 15901
rect 24489 15861 24501 15895
rect 24535 15892 24547 15895
rect 25130 15892 25136 15904
rect 24535 15864 25136 15892
rect 24535 15861 24547 15864
rect 24489 15855 24547 15861
rect 25130 15852 25136 15864
rect 25188 15892 25194 15904
rect 26142 15892 26148 15904
rect 25188 15864 26148 15892
rect 25188 15852 25194 15864
rect 26142 15852 26148 15864
rect 26200 15852 26206 15904
rect 28810 15852 28816 15904
rect 28868 15892 28874 15904
rect 28966 15892 28994 15932
rect 29641 15929 29653 15963
rect 29687 15960 29699 15963
rect 29733 15963 29791 15969
rect 29733 15960 29745 15963
rect 29687 15932 29745 15960
rect 29687 15929 29699 15932
rect 29641 15923 29699 15929
rect 29733 15929 29745 15932
rect 29779 15929 29791 15963
rect 29840 15960 29868 16000
rect 30009 15997 30021 16000
rect 30055 15997 30067 16031
rect 30009 15991 30067 15997
rect 31849 16031 31907 16037
rect 31849 15997 31861 16031
rect 31895 16028 31907 16031
rect 31938 16028 31944 16040
rect 31895 16000 31944 16028
rect 31895 15997 31907 16000
rect 31849 15991 31907 15997
rect 31938 15988 31944 16000
rect 31996 15988 32002 16040
rect 32030 15988 32036 16040
rect 32088 16028 32094 16040
rect 32140 16037 32168 16068
rect 33134 16056 33140 16068
rect 33192 16056 33198 16108
rect 32125 16031 32183 16037
rect 32125 16028 32137 16031
rect 32088 16000 32137 16028
rect 32088 15988 32094 16000
rect 32125 15997 32137 16000
rect 32171 15997 32183 16031
rect 32125 15991 32183 15997
rect 32769 16031 32827 16037
rect 32769 15997 32781 16031
rect 32815 16028 32827 16031
rect 33594 16028 33600 16040
rect 32815 16000 33600 16028
rect 32815 15997 32827 16000
rect 32769 15991 32827 15997
rect 33594 15988 33600 16000
rect 33652 15988 33658 16040
rect 29917 15963 29975 15969
rect 29917 15960 29929 15963
rect 29840 15932 29929 15960
rect 29733 15923 29791 15929
rect 29917 15929 29929 15932
rect 29963 15960 29975 15963
rect 33781 15963 33839 15969
rect 29963 15932 31708 15960
rect 29963 15929 29975 15932
rect 29917 15923 29975 15929
rect 29362 15892 29368 15904
rect 28868 15864 29368 15892
rect 28868 15852 28874 15864
rect 29362 15852 29368 15864
rect 29420 15852 29426 15904
rect 30558 15852 30564 15904
rect 30616 15892 30622 15904
rect 31680 15901 31708 15932
rect 33781 15929 33793 15963
rect 33827 15960 33839 15963
rect 34882 15960 34888 15972
rect 33827 15932 34888 15960
rect 33827 15929 33839 15932
rect 33781 15923 33839 15929
rect 34882 15920 34888 15932
rect 34940 15920 34946 15972
rect 30837 15895 30895 15901
rect 30837 15892 30849 15895
rect 30616 15864 30849 15892
rect 30616 15852 30622 15864
rect 30837 15861 30849 15864
rect 30883 15861 30895 15895
rect 30837 15855 30895 15861
rect 31665 15895 31723 15901
rect 31665 15861 31677 15895
rect 31711 15861 31723 15895
rect 31665 15855 31723 15861
rect 32398 15852 32404 15904
rect 32456 15852 32462 15904
rect 2760 15802 34316 15824
rect 2760 15750 7210 15802
rect 7262 15750 7274 15802
rect 7326 15750 7338 15802
rect 7390 15750 7402 15802
rect 7454 15750 7466 15802
rect 7518 15750 15099 15802
rect 15151 15750 15163 15802
rect 15215 15750 15227 15802
rect 15279 15750 15291 15802
rect 15343 15750 15355 15802
rect 15407 15750 22988 15802
rect 23040 15750 23052 15802
rect 23104 15750 23116 15802
rect 23168 15750 23180 15802
rect 23232 15750 23244 15802
rect 23296 15750 30877 15802
rect 30929 15750 30941 15802
rect 30993 15750 31005 15802
rect 31057 15750 31069 15802
rect 31121 15750 31133 15802
rect 31185 15750 34316 15802
rect 2760 15728 34316 15750
rect 4246 15648 4252 15700
rect 4304 15688 4310 15700
rect 4893 15691 4951 15697
rect 4893 15688 4905 15691
rect 4304 15660 4905 15688
rect 4304 15648 4310 15660
rect 4893 15657 4905 15660
rect 4939 15657 4951 15691
rect 4893 15651 4951 15657
rect 1302 15580 1308 15632
rect 1360 15620 1366 15632
rect 3237 15623 3295 15629
rect 3237 15620 3249 15623
rect 1360 15592 3249 15620
rect 1360 15580 1366 15592
rect 3237 15589 3249 15592
rect 3283 15589 3295 15623
rect 3237 15583 3295 15589
rect 4706 15580 4712 15632
rect 4764 15580 4770 15632
rect 4338 15512 4344 15564
rect 4396 15512 4402 15564
rect 4908 15484 4936 15651
rect 5442 15648 5448 15700
rect 5500 15648 5506 15700
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7009 15691 7067 15697
rect 7009 15688 7021 15691
rect 6972 15660 7021 15688
rect 6972 15648 6978 15660
rect 7009 15657 7021 15660
rect 7055 15657 7067 15691
rect 7558 15688 7564 15700
rect 7009 15651 7067 15657
rect 7116 15660 7564 15688
rect 5460 15561 5488 15648
rect 5810 15580 5816 15632
rect 5868 15620 5874 15632
rect 7116 15620 7144 15660
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 7926 15648 7932 15700
rect 7984 15688 7990 15700
rect 8021 15691 8079 15697
rect 8021 15688 8033 15691
rect 7984 15660 8033 15688
rect 7984 15648 7990 15660
rect 8021 15657 8033 15660
rect 8067 15657 8079 15691
rect 8021 15651 8079 15657
rect 9033 15691 9091 15697
rect 9033 15657 9045 15691
rect 9079 15688 9091 15691
rect 9122 15688 9128 15700
rect 9079 15660 9128 15688
rect 9079 15657 9091 15660
rect 9033 15651 9091 15657
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9674 15648 9680 15700
rect 9732 15648 9738 15700
rect 10134 15648 10140 15700
rect 10192 15688 10198 15700
rect 10229 15691 10287 15697
rect 10229 15688 10241 15691
rect 10192 15660 10241 15688
rect 10192 15648 10198 15660
rect 10229 15657 10241 15660
rect 10275 15657 10287 15691
rect 10229 15651 10287 15657
rect 11330 15648 11336 15700
rect 11388 15688 11394 15700
rect 11517 15691 11575 15697
rect 11517 15688 11529 15691
rect 11388 15660 11529 15688
rect 11388 15648 11394 15660
rect 11517 15657 11529 15660
rect 11563 15657 11575 15691
rect 11517 15651 11575 15657
rect 11974 15648 11980 15700
rect 12032 15648 12038 15700
rect 13630 15688 13636 15700
rect 12406 15660 13636 15688
rect 5868 15592 7144 15620
rect 7469 15623 7527 15629
rect 5868 15580 5874 15592
rect 7469 15589 7481 15623
rect 7515 15620 7527 15623
rect 7742 15620 7748 15632
rect 7515 15592 7748 15620
rect 7515 15589 7527 15592
rect 7469 15583 7527 15589
rect 7742 15580 7748 15592
rect 7800 15580 7806 15632
rect 9692 15620 9720 15648
rect 10689 15623 10747 15629
rect 10689 15620 10701 15623
rect 9692 15592 10701 15620
rect 10689 15589 10701 15592
rect 10735 15589 10747 15623
rect 10689 15583 10747 15589
rect 11146 15580 11152 15632
rect 11204 15580 11210 15632
rect 12406 15620 12434 15660
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 14093 15691 14151 15697
rect 14093 15657 14105 15691
rect 14139 15688 14151 15691
rect 15746 15688 15752 15700
rect 14139 15660 15752 15688
rect 14139 15657 14151 15660
rect 14093 15651 14151 15657
rect 15746 15648 15752 15660
rect 15804 15688 15810 15700
rect 17313 15691 17371 15697
rect 17313 15688 17325 15691
rect 15804 15660 17325 15688
rect 15804 15648 15810 15660
rect 17313 15657 17325 15660
rect 17359 15657 17371 15691
rect 17313 15651 17371 15657
rect 18138 15648 18144 15700
rect 18196 15688 18202 15700
rect 18693 15691 18751 15697
rect 18693 15688 18705 15691
rect 18196 15660 18705 15688
rect 18196 15648 18202 15660
rect 18693 15657 18705 15660
rect 18739 15688 18751 15691
rect 19242 15688 19248 15700
rect 18739 15660 19248 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 19242 15648 19248 15660
rect 19300 15648 19306 15700
rect 20530 15648 20536 15700
rect 20588 15648 20594 15700
rect 20714 15648 20720 15700
rect 20772 15688 20778 15700
rect 20901 15691 20959 15697
rect 20901 15688 20913 15691
rect 20772 15660 20913 15688
rect 20772 15648 20778 15660
rect 20901 15657 20913 15660
rect 20947 15657 20959 15691
rect 20901 15651 20959 15657
rect 22002 15648 22008 15700
rect 22060 15688 22066 15700
rect 23569 15691 23627 15697
rect 23569 15688 23581 15691
rect 22060 15660 23581 15688
rect 22060 15648 22066 15660
rect 23569 15657 23581 15660
rect 23615 15657 23627 15691
rect 23569 15651 23627 15657
rect 23750 15648 23756 15700
rect 23808 15688 23814 15700
rect 23845 15691 23903 15697
rect 23845 15688 23857 15691
rect 23808 15660 23857 15688
rect 23808 15648 23814 15660
rect 23845 15657 23857 15660
rect 23891 15657 23903 15691
rect 23845 15651 23903 15657
rect 24026 15648 24032 15700
rect 24084 15688 24090 15700
rect 27157 15691 27215 15697
rect 27157 15688 27169 15691
rect 24084 15660 27169 15688
rect 24084 15648 24090 15660
rect 27157 15657 27169 15660
rect 27203 15688 27215 15691
rect 27338 15688 27344 15700
rect 27203 15660 27344 15688
rect 27203 15657 27215 15660
rect 27157 15651 27215 15657
rect 27338 15648 27344 15660
rect 27396 15688 27402 15700
rect 32398 15688 32404 15700
rect 27396 15660 32404 15688
rect 27396 15648 27402 15660
rect 13170 15620 13176 15632
rect 11992 15592 12434 15620
rect 13004 15592 13176 15620
rect 5445 15555 5503 15561
rect 5445 15521 5457 15555
rect 5491 15521 5503 15555
rect 5445 15515 5503 15521
rect 5626 15512 5632 15564
rect 5684 15512 5690 15564
rect 5905 15555 5963 15561
rect 5905 15521 5917 15555
rect 5951 15521 5963 15555
rect 5905 15515 5963 15521
rect 5997 15555 6055 15561
rect 5997 15521 6009 15555
rect 6043 15552 6055 15555
rect 6270 15552 6276 15564
rect 6043 15524 6276 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 5920 15484 5948 15515
rect 6270 15512 6276 15524
rect 6328 15512 6334 15564
rect 8205 15555 8263 15561
rect 8205 15552 8217 15555
rect 7668 15524 8217 15552
rect 6365 15487 6423 15493
rect 6365 15484 6377 15487
rect 4908 15456 5948 15484
rect 6196 15456 6377 15484
rect 5718 15376 5724 15428
rect 5776 15376 5782 15428
rect 6196 15425 6224 15456
rect 6365 15453 6377 15456
rect 6411 15453 6423 15487
rect 6365 15447 6423 15453
rect 7668 15425 7696 15524
rect 8205 15521 8217 15524
rect 8251 15521 8263 15555
rect 8205 15515 8263 15521
rect 8389 15555 8447 15561
rect 8389 15521 8401 15555
rect 8435 15552 8447 15555
rect 9125 15555 9183 15561
rect 8435 15524 9076 15552
rect 8435 15521 8447 15524
rect 8389 15515 8447 15521
rect 9048 15496 9076 15524
rect 9125 15521 9137 15555
rect 9171 15552 9183 15555
rect 9766 15552 9772 15564
rect 9171 15524 9772 15552
rect 9171 15521 9183 15524
rect 9125 15515 9183 15521
rect 9766 15512 9772 15524
rect 9824 15552 9830 15564
rect 10318 15552 10324 15564
rect 9824 15524 10324 15552
rect 9824 15512 9830 15524
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 10597 15555 10655 15561
rect 10597 15521 10609 15555
rect 10643 15521 10655 15555
rect 10597 15515 10655 15521
rect 11057 15555 11115 15561
rect 11057 15521 11069 15555
rect 11103 15552 11115 15555
rect 11164 15552 11192 15580
rect 11103 15524 11192 15552
rect 11103 15521 11115 15524
rect 11057 15515 11115 15521
rect 8846 15444 8852 15496
rect 8904 15444 8910 15496
rect 9030 15444 9036 15496
rect 9088 15444 9094 15496
rect 9585 15487 9643 15493
rect 9585 15484 9597 15487
rect 9508 15456 9597 15484
rect 9508 15425 9536 15456
rect 9585 15453 9597 15456
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 10410 15444 10416 15496
rect 10468 15484 10474 15496
rect 10612 15484 10640 15515
rect 10468 15456 10640 15484
rect 10468 15444 10474 15456
rect 6181 15419 6239 15425
rect 6181 15385 6193 15419
rect 6227 15385 6239 15419
rect 6181 15379 6239 15385
rect 7101 15419 7159 15425
rect 7101 15385 7113 15419
rect 7147 15385 7159 15419
rect 7653 15419 7711 15425
rect 7653 15416 7665 15419
rect 7101 15379 7159 15385
rect 7392 15388 7665 15416
rect 5736 15348 5764 15376
rect 6362 15348 6368 15360
rect 5736 15320 6368 15348
rect 6362 15308 6368 15320
rect 6420 15348 6426 15360
rect 7006 15348 7012 15360
rect 6420 15320 7012 15348
rect 6420 15308 6426 15320
rect 7006 15308 7012 15320
rect 7064 15348 7070 15360
rect 7116 15348 7144 15379
rect 7392 15360 7420 15388
rect 7653 15385 7665 15388
rect 7699 15385 7711 15419
rect 7653 15379 7711 15385
rect 9493 15419 9551 15425
rect 9493 15385 9505 15419
rect 9539 15385 9551 15419
rect 11514 15416 11520 15428
rect 9493 15379 9551 15385
rect 11072 15388 11520 15416
rect 11072 15360 11100 15388
rect 11514 15376 11520 15388
rect 11572 15416 11578 15428
rect 11992 15416 12020 15592
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15552 12127 15555
rect 13004 15552 13032 15592
rect 13170 15580 13176 15592
rect 13228 15580 13234 15632
rect 13722 15580 13728 15632
rect 13780 15620 13786 15632
rect 14734 15620 14740 15632
rect 13780 15592 14740 15620
rect 13780 15580 13786 15592
rect 14734 15580 14740 15592
rect 14792 15580 14798 15632
rect 15470 15580 15476 15632
rect 15528 15580 15534 15632
rect 16577 15623 16635 15629
rect 16132 15592 16528 15620
rect 12115 15524 13032 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 12084 15484 12112 15515
rect 13078 15512 13084 15564
rect 13136 15512 13142 15564
rect 13188 15552 13216 15580
rect 16132 15564 16160 15592
rect 13333 15555 13391 15561
rect 13333 15552 13345 15555
rect 13188 15524 13345 15552
rect 13333 15521 13345 15524
rect 13379 15521 13391 15555
rect 13333 15515 13391 15521
rect 16114 15512 16120 15564
rect 16172 15512 16178 15564
rect 16500 15561 16528 15592
rect 16577 15589 16589 15623
rect 16623 15620 16635 15623
rect 17402 15620 17408 15632
rect 16623 15592 17408 15620
rect 16623 15589 16635 15592
rect 16577 15583 16635 15589
rect 17402 15580 17408 15592
rect 17460 15580 17466 15632
rect 17678 15620 17684 15632
rect 17512 15592 17684 15620
rect 16301 15555 16359 15561
rect 16301 15521 16313 15555
rect 16347 15521 16359 15555
rect 16301 15515 16359 15521
rect 16485 15555 16543 15561
rect 16485 15521 16497 15555
rect 16531 15521 16543 15555
rect 16485 15515 16543 15521
rect 16669 15555 16727 15561
rect 16669 15521 16681 15555
rect 16715 15552 16727 15555
rect 17512 15552 17540 15592
rect 17678 15580 17684 15592
rect 17736 15580 17742 15632
rect 20548 15620 20576 15648
rect 19306 15592 20576 15620
rect 16715 15524 17540 15552
rect 17589 15555 17647 15561
rect 16715 15521 16727 15524
rect 16669 15515 16727 15521
rect 17589 15521 17601 15555
rect 17635 15552 17647 15555
rect 18046 15552 18052 15564
rect 17635 15524 18052 15552
rect 17635 15521 17647 15524
rect 17589 15515 17647 15521
rect 12158 15484 12164 15496
rect 12084 15456 12164 15484
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 12802 15444 12808 15496
rect 12860 15444 12866 15496
rect 13096 15484 13124 15512
rect 13906 15484 13912 15496
rect 13096 15456 13912 15484
rect 13906 15444 13912 15456
rect 13964 15484 13970 15496
rect 14185 15487 14243 15493
rect 14185 15484 14197 15487
rect 13964 15456 14197 15484
rect 13964 15444 13970 15456
rect 14185 15453 14197 15456
rect 14231 15453 14243 15487
rect 14461 15487 14519 15493
rect 14461 15484 14473 15487
rect 14185 15447 14243 15453
rect 14292 15456 14473 15484
rect 12437 15419 12495 15425
rect 12437 15416 12449 15419
rect 11572 15388 12449 15416
rect 11572 15376 11578 15388
rect 12437 15385 12449 15388
rect 12483 15385 12495 15419
rect 12437 15379 12495 15385
rect 12820 15416 12848 15444
rect 13446 15416 13452 15428
rect 12820 15388 13452 15416
rect 7064 15320 7144 15348
rect 7064 15308 7070 15320
rect 7374 15308 7380 15360
rect 7432 15308 7438 15360
rect 7469 15351 7527 15357
rect 7469 15317 7481 15351
rect 7515 15348 7527 15351
rect 8018 15348 8024 15360
rect 7515 15320 8024 15348
rect 7515 15317 7527 15320
rect 7469 15311 7527 15317
rect 8018 15308 8024 15320
rect 8076 15348 8082 15360
rect 11054 15348 11060 15360
rect 8076 15320 11060 15348
rect 8076 15308 8082 15320
rect 11054 15308 11060 15320
rect 11112 15308 11118 15360
rect 11146 15308 11152 15360
rect 11204 15348 11210 15360
rect 12820 15348 12848 15388
rect 13446 15376 13452 15388
rect 13504 15376 13510 15428
rect 14292 15360 14320 15456
rect 14461 15453 14473 15456
rect 14507 15453 14519 15487
rect 14461 15447 14519 15453
rect 15838 15444 15844 15496
rect 15896 15444 15902 15496
rect 16316 15484 16344 15515
rect 18046 15512 18052 15524
rect 18104 15512 18110 15564
rect 18874 15512 18880 15564
rect 18932 15552 18938 15564
rect 19306 15552 19334 15592
rect 26694 15580 26700 15632
rect 26752 15620 26758 15632
rect 26752 15592 27568 15620
rect 26752 15580 26758 15592
rect 20533 15555 20591 15561
rect 20533 15552 20545 15555
rect 18932 15524 19334 15552
rect 19444 15524 20545 15552
rect 18932 15512 18938 15524
rect 19444 15496 19472 15524
rect 20533 15521 20545 15524
rect 20579 15521 20591 15555
rect 20533 15515 20591 15521
rect 22186 15512 22192 15564
rect 22244 15552 22250 15564
rect 22373 15555 22431 15561
rect 22373 15552 22385 15555
rect 22244 15524 22385 15552
rect 22244 15512 22250 15524
rect 22373 15521 22385 15524
rect 22419 15521 22431 15555
rect 22373 15515 22431 15521
rect 23201 15555 23259 15561
rect 23201 15521 23213 15555
rect 23247 15552 23259 15555
rect 23474 15552 23480 15564
rect 23247 15524 23480 15552
rect 23247 15521 23259 15524
rect 23201 15515 23259 15521
rect 23474 15512 23480 15524
rect 23532 15512 23538 15564
rect 23661 15555 23719 15561
rect 23661 15521 23673 15555
rect 23707 15552 23719 15555
rect 23750 15552 23756 15564
rect 23707 15524 23756 15552
rect 23707 15521 23719 15524
rect 23661 15515 23719 15521
rect 23750 15512 23756 15524
rect 23808 15512 23814 15564
rect 27430 15512 27436 15564
rect 27488 15512 27494 15564
rect 27540 15561 27568 15592
rect 27982 15580 27988 15632
rect 28040 15580 28046 15632
rect 28721 15623 28779 15629
rect 28721 15589 28733 15623
rect 28767 15620 28779 15623
rect 28994 15620 29000 15632
rect 28767 15592 29000 15620
rect 28767 15589 28779 15592
rect 28721 15583 28779 15589
rect 28994 15580 29000 15592
rect 29052 15580 29058 15632
rect 30285 15623 30343 15629
rect 30285 15589 30297 15623
rect 30331 15620 30343 15623
rect 30558 15620 30564 15632
rect 30331 15592 30564 15620
rect 30331 15589 30343 15592
rect 30285 15583 30343 15589
rect 30558 15580 30564 15592
rect 30616 15580 30622 15632
rect 31294 15580 31300 15632
rect 31352 15580 31358 15632
rect 31864 15629 31892 15660
rect 32398 15648 32404 15660
rect 32456 15648 32462 15700
rect 32950 15648 32956 15700
rect 33008 15688 33014 15700
rect 33137 15691 33195 15697
rect 33137 15688 33149 15691
rect 33008 15660 33149 15688
rect 33008 15648 33014 15660
rect 33137 15657 33149 15660
rect 33183 15657 33195 15691
rect 33137 15651 33195 15657
rect 31849 15623 31907 15629
rect 31849 15589 31861 15623
rect 31895 15620 31907 15623
rect 31895 15592 31929 15620
rect 31895 15589 31907 15592
rect 31849 15583 31907 15589
rect 27525 15555 27583 15561
rect 27525 15521 27537 15555
rect 27571 15521 27583 15555
rect 28000 15552 28028 15580
rect 28077 15555 28135 15561
rect 28077 15552 28089 15555
rect 28000 15524 28089 15552
rect 27525 15515 27583 15521
rect 28077 15521 28089 15524
rect 28123 15552 28135 15555
rect 28626 15552 28632 15564
rect 28123 15524 28632 15552
rect 28123 15521 28135 15524
rect 28077 15515 28135 15521
rect 28626 15512 28632 15524
rect 28684 15512 28690 15564
rect 29181 15555 29239 15561
rect 29181 15521 29193 15555
rect 29227 15552 29239 15555
rect 29914 15552 29920 15564
rect 29227 15524 29920 15552
rect 29227 15521 29239 15524
rect 29181 15515 29239 15521
rect 16945 15487 17003 15493
rect 16945 15484 16957 15487
rect 16316 15456 16957 15484
rect 16945 15453 16957 15456
rect 16991 15453 17003 15487
rect 16945 15447 17003 15453
rect 17034 15444 17040 15496
rect 17092 15484 17098 15496
rect 17129 15487 17187 15493
rect 17129 15484 17141 15487
rect 17092 15456 17141 15484
rect 17092 15444 17098 15456
rect 17129 15453 17141 15456
rect 17175 15453 17187 15487
rect 17129 15447 17187 15453
rect 17218 15444 17224 15496
rect 17276 15444 17282 15496
rect 17497 15487 17555 15493
rect 17497 15453 17509 15487
rect 17543 15453 17555 15487
rect 17497 15447 17555 15453
rect 15856 15416 15884 15444
rect 17512 15416 17540 15447
rect 19334 15444 19340 15496
rect 19392 15444 19398 15496
rect 19426 15444 19432 15496
rect 19484 15444 19490 15496
rect 20162 15444 20168 15496
rect 20220 15484 20226 15496
rect 20622 15484 20628 15496
rect 20220 15456 20628 15484
rect 20220 15444 20226 15456
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 20898 15444 20904 15496
rect 20956 15484 20962 15496
rect 21453 15487 21511 15493
rect 21453 15484 21465 15487
rect 20956 15456 21465 15484
rect 20956 15444 20962 15456
rect 21453 15453 21465 15456
rect 21499 15453 21511 15487
rect 21453 15447 21511 15453
rect 27890 15444 27896 15496
rect 27948 15484 27954 15496
rect 28902 15484 28908 15496
rect 27948 15456 28908 15484
rect 27948 15444 27954 15456
rect 28902 15444 28908 15456
rect 28960 15444 28966 15496
rect 19886 15416 19892 15428
rect 15856 15388 16988 15416
rect 17512 15388 19892 15416
rect 11204 15320 12848 15348
rect 11204 15308 11210 15320
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 13265 15351 13323 15357
rect 13265 15348 13277 15351
rect 13228 15320 13277 15348
rect 13228 15308 13234 15320
rect 13265 15317 13277 15320
rect 13311 15317 13323 15351
rect 13265 15311 13323 15317
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 15933 15351 15991 15357
rect 15933 15317 15945 15351
rect 15979 15348 15991 15351
rect 16482 15348 16488 15360
rect 15979 15320 16488 15348
rect 15979 15317 15991 15320
rect 15933 15311 15991 15317
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 16758 15308 16764 15360
rect 16816 15348 16822 15360
rect 16853 15351 16911 15357
rect 16853 15348 16865 15351
rect 16816 15320 16865 15348
rect 16816 15308 16822 15320
rect 16853 15317 16865 15320
rect 16899 15317 16911 15351
rect 16960 15348 16988 15388
rect 19886 15376 19892 15388
rect 19944 15376 19950 15428
rect 26602 15376 26608 15428
rect 26660 15416 26666 15428
rect 26970 15416 26976 15428
rect 26660 15388 26976 15416
rect 26660 15376 26666 15388
rect 26970 15376 26976 15388
rect 27028 15416 27034 15428
rect 29196 15416 29224 15515
rect 29914 15512 29920 15524
rect 29972 15512 29978 15564
rect 30009 15487 30067 15493
rect 30009 15453 30021 15487
rect 30055 15453 30067 15487
rect 30009 15447 30067 15453
rect 27028 15388 29224 15416
rect 27028 15376 27034 15388
rect 18049 15351 18107 15357
rect 18049 15348 18061 15351
rect 16960 15320 18061 15348
rect 16853 15311 16911 15317
rect 18049 15317 18061 15320
rect 18095 15348 18107 15351
rect 18874 15348 18880 15360
rect 18095 15320 18880 15348
rect 18095 15317 18107 15320
rect 18049 15311 18107 15317
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 19978 15308 19984 15360
rect 20036 15308 20042 15360
rect 21818 15308 21824 15360
rect 21876 15308 21882 15360
rect 23017 15351 23075 15357
rect 23017 15317 23029 15351
rect 23063 15348 23075 15351
rect 23382 15348 23388 15360
rect 23063 15320 23388 15348
rect 23063 15317 23075 15320
rect 23017 15311 23075 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 27154 15308 27160 15360
rect 27212 15348 27218 15360
rect 27709 15351 27767 15357
rect 27709 15348 27721 15351
rect 27212 15320 27721 15348
rect 27212 15308 27218 15320
rect 27709 15317 27721 15320
rect 27755 15317 27767 15351
rect 27709 15311 27767 15317
rect 28074 15308 28080 15360
rect 28132 15348 28138 15360
rect 28169 15351 28227 15357
rect 28169 15348 28181 15351
rect 28132 15320 28181 15348
rect 28132 15308 28138 15320
rect 28169 15317 28181 15320
rect 28215 15317 28227 15351
rect 30024 15348 30052 15447
rect 31757 15419 31815 15425
rect 31757 15385 31769 15419
rect 31803 15416 31815 15419
rect 31938 15416 31944 15428
rect 31803 15388 31944 15416
rect 31803 15385 31815 15388
rect 31757 15379 31815 15385
rect 31938 15376 31944 15388
rect 31996 15376 32002 15428
rect 31846 15348 31852 15360
rect 30024 15320 31852 15348
rect 28169 15311 28227 15317
rect 31846 15308 31852 15320
rect 31904 15348 31910 15360
rect 32968 15348 32996 15648
rect 33134 15512 33140 15564
rect 33192 15552 33198 15564
rect 33781 15555 33839 15561
rect 33781 15552 33793 15555
rect 33192 15524 33793 15552
rect 33192 15512 33198 15524
rect 33781 15521 33793 15524
rect 33827 15521 33839 15555
rect 33781 15515 33839 15521
rect 31904 15320 32996 15348
rect 31904 15308 31910 15320
rect 33870 15308 33876 15360
rect 33928 15308 33934 15360
rect 2760 15258 34316 15280
rect 2760 15206 6550 15258
rect 6602 15206 6614 15258
rect 6666 15206 6678 15258
rect 6730 15206 6742 15258
rect 6794 15206 6806 15258
rect 6858 15206 14439 15258
rect 14491 15206 14503 15258
rect 14555 15206 14567 15258
rect 14619 15206 14631 15258
rect 14683 15206 14695 15258
rect 14747 15206 22328 15258
rect 22380 15206 22392 15258
rect 22444 15206 22456 15258
rect 22508 15206 22520 15258
rect 22572 15206 22584 15258
rect 22636 15206 30217 15258
rect 30269 15206 30281 15258
rect 30333 15206 30345 15258
rect 30397 15206 30409 15258
rect 30461 15206 30473 15258
rect 30525 15206 34316 15258
rect 2760 15184 34316 15206
rect 4893 15147 4951 15153
rect 4893 15113 4905 15147
rect 4939 15144 4951 15147
rect 5258 15144 5264 15156
rect 4939 15116 5264 15144
rect 4939 15113 4951 15116
rect 4893 15107 4951 15113
rect 5258 15104 5264 15116
rect 5316 15144 5322 15156
rect 5810 15144 5816 15156
rect 5316 15116 5816 15144
rect 5316 15104 5322 15116
rect 5810 15104 5816 15116
rect 5868 15104 5874 15156
rect 5902 15104 5908 15156
rect 5960 15144 5966 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5960 15116 6009 15144
rect 5960 15104 5966 15116
rect 5997 15113 6009 15116
rect 6043 15113 6055 15147
rect 5997 15107 6055 15113
rect 6270 15104 6276 15156
rect 6328 15144 6334 15156
rect 6365 15147 6423 15153
rect 6365 15144 6377 15147
rect 6328 15116 6377 15144
rect 6328 15104 6334 15116
rect 6365 15113 6377 15116
rect 6411 15113 6423 15147
rect 6365 15107 6423 15113
rect 6825 15147 6883 15153
rect 6825 15113 6837 15147
rect 6871 15144 6883 15147
rect 7006 15144 7012 15156
rect 6871 15116 7012 15144
rect 6871 15113 6883 15116
rect 6825 15107 6883 15113
rect 7006 15104 7012 15116
rect 7064 15144 7070 15156
rect 7064 15116 7696 15144
rect 7064 15104 7070 15116
rect 3789 15079 3847 15085
rect 3789 15076 3801 15079
rect 3712 15048 3801 15076
rect 3712 15017 3740 15048
rect 3789 15045 3801 15048
rect 3835 15045 3847 15079
rect 5074 15076 5080 15088
rect 3789 15039 3847 15045
rect 4356 15048 5080 15076
rect 4356 15020 4384 15048
rect 5074 15036 5080 15048
rect 5132 15076 5138 15088
rect 5169 15079 5227 15085
rect 5169 15076 5181 15079
rect 5132 15048 5181 15076
rect 5132 15036 5138 15048
rect 5169 15045 5181 15048
rect 5215 15045 5227 15079
rect 5169 15039 5227 15045
rect 5718 15036 5724 15088
rect 5776 15076 5782 15088
rect 5776 15048 7039 15076
rect 5776 15036 5782 15048
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 4338 14968 4344 15020
rect 4396 14968 4402 15020
rect 4430 14968 4436 15020
rect 4488 14968 4494 15020
rect 5350 14968 5356 15020
rect 5408 14968 5414 15020
rect 7011 15008 7039 15048
rect 7668 15008 7696 15116
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8202 15144 8208 15156
rect 7892 15116 8208 15144
rect 7892 15104 7898 15116
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 10410 15144 10416 15156
rect 8352 15116 10416 15144
rect 8352 15104 8358 15116
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 11054 15104 11060 15156
rect 11112 15104 11118 15156
rect 14826 15104 14832 15156
rect 14884 15104 14890 15156
rect 17862 15144 17868 15156
rect 16868 15116 17868 15144
rect 7742 15036 7748 15088
rect 7800 15076 7806 15088
rect 11330 15076 11336 15088
rect 7800 15048 11336 15076
rect 7800 15036 7806 15048
rect 11330 15036 11336 15048
rect 11388 15036 11394 15088
rect 16758 15076 16764 15088
rect 15212 15048 16764 15076
rect 7011 14980 7512 15008
rect 7668 14980 8892 15008
rect 4249 14943 4307 14949
rect 4249 14909 4261 14943
rect 4295 14940 4307 14943
rect 4448 14940 4476 14968
rect 4295 14912 4476 14940
rect 4295 14909 4307 14912
rect 4249 14903 4307 14909
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 5368 14940 5396 14968
rect 5905 14943 5963 14949
rect 5905 14940 5917 14943
rect 5224 14912 5917 14940
rect 5224 14900 5230 14912
rect 5905 14909 5917 14912
rect 5951 14909 5963 14943
rect 5905 14903 5963 14909
rect 6270 14900 6276 14952
rect 6328 14940 6334 14952
rect 7484 14949 7512 14980
rect 7055 14943 7113 14949
rect 7055 14940 7067 14943
rect 6328 14912 7067 14940
rect 6328 14900 6334 14912
rect 7055 14909 7067 14912
rect 7101 14909 7113 14943
rect 7055 14903 7113 14909
rect 7193 14943 7251 14949
rect 7193 14909 7205 14943
rect 7239 14940 7251 14943
rect 7469 14943 7527 14949
rect 7300 14940 7420 14942
rect 7239 14914 7420 14940
rect 7239 14912 7328 14914
rect 7239 14909 7251 14912
rect 7193 14903 7251 14909
rect 7285 14875 7343 14881
rect 7285 14841 7297 14875
rect 7331 14841 7343 14875
rect 7392 14872 7420 14914
rect 7469 14909 7481 14943
rect 7515 14940 7527 14943
rect 7515 14912 8616 14940
rect 7515 14909 7527 14912
rect 7469 14903 7527 14909
rect 7558 14872 7564 14884
rect 7392 14844 7564 14872
rect 7285 14835 7343 14841
rect 3053 14807 3111 14813
rect 3053 14804 3065 14807
rect 2700 14776 3065 14804
rect 2700 14600 2728 14776
rect 3053 14773 3065 14776
rect 3099 14773 3111 14807
rect 3053 14767 3111 14773
rect 4154 14764 4160 14816
rect 4212 14764 4218 14816
rect 6914 14764 6920 14816
rect 6972 14764 6978 14816
rect 7300 14804 7328 14835
rect 7558 14832 7564 14844
rect 7616 14872 7622 14884
rect 8021 14875 8079 14881
rect 8021 14872 8033 14875
rect 7616 14844 8033 14872
rect 7616 14832 7622 14844
rect 8021 14841 8033 14844
rect 8067 14841 8079 14875
rect 8588 14872 8616 14912
rect 8662 14900 8668 14952
rect 8720 14900 8726 14952
rect 8754 14872 8760 14884
rect 8588 14844 8760 14872
rect 8021 14835 8079 14841
rect 8754 14832 8760 14844
rect 8812 14832 8818 14884
rect 8864 14872 8892 14980
rect 9950 14968 9956 15020
rect 10008 15008 10014 15020
rect 10597 15011 10655 15017
rect 10597 15008 10609 15011
rect 10008 14980 10609 15008
rect 10008 14968 10014 14980
rect 10597 14977 10609 14980
rect 10643 15008 10655 15011
rect 11146 15008 11152 15020
rect 10643 14980 11152 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 11885 15011 11943 15017
rect 11885 14977 11897 15011
rect 11931 15008 11943 15011
rect 13262 15008 13268 15020
rect 11931 14980 13268 15008
rect 11931 14977 11943 14980
rect 11885 14971 11943 14977
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13906 14968 13912 15020
rect 13964 14968 13970 15020
rect 15212 15008 15240 15048
rect 16758 15036 16764 15048
rect 16816 15036 16822 15088
rect 14108 14980 15240 15008
rect 10134 14900 10140 14952
rect 10192 14940 10198 14952
rect 10321 14943 10379 14949
rect 10321 14940 10333 14943
rect 10192 14912 10333 14940
rect 10192 14900 10198 14912
rect 10321 14909 10333 14912
rect 10367 14909 10379 14943
rect 10962 14940 10968 14952
rect 10321 14903 10379 14909
rect 10704 14912 10968 14940
rect 9677 14875 9735 14881
rect 9677 14872 9689 14875
rect 8864 14844 9689 14872
rect 9677 14841 9689 14844
rect 9723 14872 9735 14875
rect 10704 14872 10732 14912
rect 10962 14900 10968 14912
rect 11020 14900 11026 14952
rect 11609 14943 11667 14949
rect 11609 14909 11621 14943
rect 11655 14940 11667 14943
rect 11655 14912 12204 14940
rect 11655 14909 11667 14912
rect 11609 14903 11667 14909
rect 12176 14884 12204 14912
rect 12066 14872 12072 14884
rect 9723 14844 10732 14872
rect 10796 14844 12072 14872
rect 9723 14841 9735 14844
rect 9677 14835 9735 14841
rect 7374 14804 7380 14816
rect 7300 14776 7380 14804
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 9030 14764 9036 14816
rect 9088 14764 9094 14816
rect 9766 14764 9772 14816
rect 9824 14764 9830 14816
rect 10502 14764 10508 14816
rect 10560 14804 10566 14816
rect 10796 14813 10824 14844
rect 12066 14832 12072 14844
rect 12124 14832 12130 14884
rect 12158 14832 12164 14884
rect 12216 14832 12222 14884
rect 13170 14832 13176 14884
rect 13228 14832 13234 14884
rect 13630 14832 13636 14884
rect 13688 14832 13694 14884
rect 14108 14872 14136 14980
rect 14182 14900 14188 14952
rect 14240 14900 14246 14952
rect 14734 14900 14740 14952
rect 14792 14900 14798 14952
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 15212 14940 15240 14980
rect 15289 15011 15347 15017
rect 15289 14977 15301 15011
rect 15335 15008 15347 15011
rect 15335 14980 15976 15008
rect 15335 14977 15347 14980
rect 15289 14971 15347 14977
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 14875 14912 15148 14940
rect 15212 14912 15393 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 13832 14844 14136 14872
rect 14200 14872 14228 14900
rect 14921 14875 14979 14881
rect 14921 14872 14933 14875
rect 14200 14844 14933 14872
rect 13832 14816 13860 14844
rect 14921 14841 14933 14844
rect 14967 14841 14979 14875
rect 15120 14872 15148 14912
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 15838 14900 15844 14952
rect 15896 14900 15902 14952
rect 15948 14940 15976 14980
rect 16482 14968 16488 15020
rect 16540 15008 16546 15020
rect 16868 15017 16896 15116
rect 17862 15104 17868 15116
rect 17920 15104 17926 15156
rect 17954 15104 17960 15156
rect 18012 15144 18018 15156
rect 18414 15144 18420 15156
rect 18012 15116 18420 15144
rect 18012 15104 18018 15116
rect 18414 15104 18420 15116
rect 18472 15104 18478 15156
rect 19426 15144 19432 15156
rect 18524 15116 19432 15144
rect 17497 15079 17555 15085
rect 17497 15045 17509 15079
rect 17543 15076 17555 15079
rect 18138 15076 18144 15088
rect 17543 15048 18144 15076
rect 17543 15045 17555 15048
rect 17497 15039 17555 15045
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 16853 15011 16911 15017
rect 16853 15008 16865 15011
rect 16540 14980 16865 15008
rect 16540 14968 16546 14980
rect 16853 14977 16865 14980
rect 16899 14977 16911 15011
rect 16853 14971 16911 14977
rect 17126 14968 17132 15020
rect 17184 15008 17190 15020
rect 18524 15017 18552 15116
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 19613 15147 19671 15153
rect 19613 15113 19625 15147
rect 19659 15144 19671 15147
rect 19659 15116 19932 15144
rect 19659 15113 19671 15116
rect 19613 15107 19671 15113
rect 19904 15088 19932 15116
rect 20438 15104 20444 15156
rect 20496 15144 20502 15156
rect 20496 15116 21956 15144
rect 20496 15104 20502 15116
rect 18601 15079 18659 15085
rect 18601 15045 18613 15079
rect 18647 15045 18659 15079
rect 18601 15039 18659 15045
rect 17865 15011 17923 15017
rect 17865 15008 17877 15011
rect 17184 14980 17877 15008
rect 17184 14968 17190 14980
rect 17865 14977 17877 14980
rect 17911 14977 17923 15011
rect 17865 14971 17923 14977
rect 18509 15011 18567 15017
rect 18509 14977 18521 15011
rect 18555 14977 18567 15011
rect 18616 15008 18644 15039
rect 18690 15036 18696 15088
rect 18748 15076 18754 15088
rect 19797 15079 19855 15085
rect 19797 15076 19809 15079
rect 18748 15048 19809 15076
rect 18748 15036 18754 15048
rect 19797 15045 19809 15048
rect 19843 15045 19855 15079
rect 19797 15039 19855 15045
rect 19886 15036 19892 15088
rect 19944 15076 19950 15088
rect 20165 15079 20223 15085
rect 20165 15076 20177 15079
rect 19944 15048 20177 15076
rect 19944 15036 19950 15048
rect 20165 15045 20177 15048
rect 20211 15045 20223 15079
rect 21634 15076 21640 15088
rect 20165 15039 20223 15045
rect 20272 15048 21640 15076
rect 20073 15011 20131 15017
rect 18616 14980 19472 15008
rect 18509 14971 18567 14977
rect 16666 14940 16672 14952
rect 15948 14912 16672 14940
rect 16666 14900 16672 14912
rect 16724 14940 16730 14952
rect 16942 14940 16948 14952
rect 16724 14912 16948 14940
rect 16724 14900 16730 14912
rect 16942 14900 16948 14912
rect 17000 14900 17006 14952
rect 17589 14943 17647 14949
rect 17589 14909 17601 14943
rect 17635 14940 17647 14943
rect 17678 14940 17684 14952
rect 17635 14912 17684 14940
rect 17635 14909 17647 14912
rect 17589 14903 17647 14909
rect 17678 14900 17684 14912
rect 17736 14900 17742 14952
rect 17773 14943 17831 14949
rect 17773 14909 17785 14943
rect 17819 14940 17831 14943
rect 17819 14912 17899 14940
rect 17819 14909 17831 14912
rect 17773 14903 17831 14909
rect 15120 14844 15516 14872
rect 14921 14835 14979 14841
rect 15488 14816 15516 14844
rect 16206 14832 16212 14884
rect 16264 14872 16270 14884
rect 16577 14875 16635 14881
rect 16577 14872 16589 14875
rect 16264 14844 16589 14872
rect 16264 14832 16270 14844
rect 16577 14841 16589 14844
rect 16623 14841 16635 14875
rect 16577 14835 16635 14841
rect 10781 14807 10839 14813
rect 10781 14804 10793 14807
rect 10560 14776 10793 14804
rect 10560 14764 10566 14776
rect 10781 14773 10793 14776
rect 10827 14773 10839 14807
rect 10781 14767 10839 14773
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11517 14807 11575 14813
rect 11517 14804 11529 14807
rect 11480 14776 11529 14804
rect 11480 14764 11486 14776
rect 11517 14773 11529 14776
rect 11563 14773 11575 14807
rect 11517 14767 11575 14773
rect 13814 14764 13820 14816
rect 13872 14764 13878 14816
rect 13906 14764 13912 14816
rect 13964 14804 13970 14816
rect 14185 14807 14243 14813
rect 14185 14804 14197 14807
rect 13964 14776 14197 14804
rect 13964 14764 13970 14776
rect 14185 14773 14197 14776
rect 14231 14773 14243 14807
rect 14185 14767 14243 14773
rect 14458 14764 14464 14816
rect 14516 14764 14522 14816
rect 15470 14764 15476 14816
rect 15528 14764 15534 14816
rect 15562 14764 15568 14816
rect 15620 14764 15626 14816
rect 16114 14764 16120 14816
rect 16172 14804 16178 14816
rect 17310 14804 17316 14816
rect 16172 14776 17316 14804
rect 16172 14764 16178 14776
rect 17310 14764 17316 14776
rect 17368 14804 17374 14816
rect 17681 14807 17739 14813
rect 17681 14804 17693 14807
rect 17368 14776 17693 14804
rect 17368 14764 17374 14776
rect 17681 14773 17693 14776
rect 17727 14773 17739 14807
rect 17871 14804 17899 14912
rect 17954 14900 17960 14952
rect 18012 14940 18018 14952
rect 18601 14943 18659 14949
rect 18601 14940 18613 14943
rect 18012 14912 18613 14940
rect 18012 14900 18018 14912
rect 18601 14909 18613 14912
rect 18647 14909 18659 14943
rect 18601 14903 18659 14909
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 19444 14949 19472 14980
rect 20073 14977 20085 15011
rect 20119 15008 20131 15011
rect 20272 15008 20300 15048
rect 21634 15036 21640 15048
rect 21692 15036 21698 15088
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20119 14980 20300 15008
rect 20364 14980 21097 15008
rect 20119 14977 20131 14980
rect 20073 14971 20131 14977
rect 19429 14943 19487 14949
rect 19429 14909 19441 14943
rect 19475 14909 19487 14943
rect 19429 14903 19487 14909
rect 19978 14900 19984 14952
rect 20036 14900 20042 14952
rect 18874 14832 18880 14884
rect 18932 14832 18938 14884
rect 20088 14872 20116 14971
rect 18984 14844 20116 14872
rect 18984 14804 19012 14844
rect 17871 14776 19012 14804
rect 17681 14767 17739 14773
rect 19242 14764 19248 14816
rect 19300 14804 19306 14816
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 19300 14776 19349 14804
rect 19300 14764 19306 14776
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 19337 14767 19395 14773
rect 19886 14764 19892 14816
rect 19944 14804 19950 14816
rect 20364 14804 20392 14980
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 21177 15011 21235 15017
rect 21177 14977 21189 15011
rect 21223 15008 21235 15011
rect 21818 15008 21824 15020
rect 21223 14980 21824 15008
rect 21223 14977 21235 14980
rect 21177 14971 21235 14977
rect 21818 14968 21824 14980
rect 21876 14968 21882 15020
rect 21928 15017 21956 15116
rect 23474 15104 23480 15156
rect 23532 15144 23538 15156
rect 23799 15147 23857 15153
rect 23799 15144 23811 15147
rect 23532 15116 23811 15144
rect 23532 15104 23538 15116
rect 23799 15113 23811 15116
rect 23845 15113 23857 15147
rect 27522 15144 27528 15156
rect 23799 15107 23857 15113
rect 27080 15116 27528 15144
rect 23201 15079 23259 15085
rect 23201 15045 23213 15079
rect 23247 15076 23259 15079
rect 24394 15076 24400 15088
rect 23247 15048 24400 15076
rect 23247 15045 23259 15048
rect 23201 15039 23259 15045
rect 24394 15036 24400 15048
rect 24452 15036 24458 15088
rect 27080 15017 27108 15116
rect 27522 15104 27528 15116
rect 27580 15104 27586 15156
rect 31294 15104 31300 15156
rect 31352 15104 31358 15156
rect 33594 15104 33600 15156
rect 33652 15104 33658 15156
rect 21913 15011 21971 15017
rect 21913 14977 21925 15011
rect 21959 14977 21971 15011
rect 21913 14971 21971 14977
rect 25593 15011 25651 15017
rect 25593 14977 25605 15011
rect 25639 15008 25651 15011
rect 27065 15011 27123 15017
rect 27065 15008 27077 15011
rect 25639 14980 27077 15008
rect 25639 14977 25651 14980
rect 25593 14971 25651 14977
rect 27065 14977 27077 14980
rect 27111 14977 27123 15011
rect 27065 14971 27123 14977
rect 28718 14968 28724 15020
rect 28776 14968 28782 15020
rect 31846 14968 31852 15020
rect 31904 14968 31910 15020
rect 20898 14900 20904 14952
rect 20956 14900 20962 14952
rect 22281 14943 22339 14949
rect 22281 14940 22293 14943
rect 21192 14912 22293 14940
rect 20530 14832 20536 14884
rect 20588 14832 20594 14884
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 21192 14872 21220 14912
rect 22281 14909 22293 14912
rect 22327 14909 22339 14943
rect 22281 14903 22339 14909
rect 21796 14875 21854 14881
rect 20772 14844 21220 14872
rect 21284 14844 21680 14872
rect 20772 14832 20778 14844
rect 19944 14776 20392 14804
rect 19944 14764 19950 14776
rect 20622 14764 20628 14816
rect 20680 14804 20686 14816
rect 21284 14804 21312 14844
rect 20680 14776 21312 14804
rect 20680 14764 20686 14776
rect 21542 14764 21548 14816
rect 21600 14764 21606 14816
rect 21652 14813 21680 14844
rect 21796 14841 21808 14875
rect 21842 14872 21854 14875
rect 22094 14872 22100 14884
rect 21842 14844 22100 14872
rect 21842 14841 21854 14844
rect 21796 14835 21854 14841
rect 22094 14832 22100 14844
rect 22152 14832 22158 14884
rect 22296 14872 22324 14903
rect 22462 14900 22468 14952
rect 22520 14900 22526 14952
rect 23109 14943 23167 14949
rect 23109 14909 23121 14943
rect 23155 14909 23167 14943
rect 23109 14903 23167 14909
rect 23293 14943 23351 14949
rect 23293 14909 23305 14943
rect 23339 14940 23351 14943
rect 25225 14943 25283 14949
rect 23339 14912 23428 14940
rect 23339 14909 23351 14912
rect 23293 14903 23351 14909
rect 23017 14875 23075 14881
rect 23017 14872 23029 14875
rect 22296 14844 23029 14872
rect 23017 14841 23029 14844
rect 23063 14872 23075 14875
rect 23124 14872 23152 14903
rect 23063 14844 23152 14872
rect 23063 14841 23075 14844
rect 23017 14835 23075 14841
rect 23400 14816 23428 14912
rect 25225 14909 25237 14943
rect 25271 14940 25283 14943
rect 26053 14943 26111 14949
rect 26053 14940 26065 14943
rect 25271 14912 26065 14940
rect 25271 14909 25283 14912
rect 25225 14903 25283 14909
rect 26053 14909 26065 14912
rect 26099 14909 26111 14943
rect 26053 14903 26111 14909
rect 26694 14900 26700 14952
rect 26752 14900 26758 14952
rect 28736 14940 28764 14968
rect 29089 14943 29147 14949
rect 29089 14940 29101 14943
rect 28736 14912 29101 14940
rect 29089 14909 29101 14912
rect 29135 14909 29147 14943
rect 29089 14903 29147 14909
rect 29822 14900 29828 14952
rect 29880 14900 29886 14952
rect 30006 14900 30012 14952
rect 30064 14900 30070 14952
rect 31389 14943 31447 14949
rect 31389 14909 31401 14943
rect 31435 14909 31447 14943
rect 31389 14903 31447 14909
rect 31665 14943 31723 14949
rect 31665 14909 31677 14943
rect 31711 14940 31723 14943
rect 33870 14940 33876 14952
rect 31711 14912 31745 14940
rect 33258 14912 33876 14940
rect 31711 14909 31723 14912
rect 31665 14903 31723 14909
rect 24670 14832 24676 14884
rect 24728 14832 24734 14884
rect 27338 14832 27344 14884
rect 27396 14832 27402 14884
rect 28074 14832 28080 14884
rect 28132 14832 28138 14884
rect 28626 14832 28632 14884
rect 28684 14872 28690 14884
rect 31404 14872 31432 14903
rect 31680 14872 31708 14903
rect 33870 14900 33876 14912
rect 33928 14900 33934 14952
rect 32030 14872 32036 14884
rect 28684 14844 32036 14872
rect 28684 14832 28690 14844
rect 32030 14832 32036 14844
rect 32088 14832 32094 14884
rect 32122 14832 32128 14884
rect 32180 14832 32186 14884
rect 21637 14807 21695 14813
rect 21637 14773 21649 14807
rect 21683 14773 21695 14807
rect 21637 14767 21695 14773
rect 22002 14764 22008 14816
rect 22060 14804 22066 14816
rect 23382 14804 23388 14816
rect 22060 14776 23388 14804
rect 22060 14764 22066 14776
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 29273 14807 29331 14813
rect 29273 14773 29285 14807
rect 29319 14804 29331 14807
rect 29454 14804 29460 14816
rect 29319 14776 29460 14804
rect 29319 14773 29331 14776
rect 29273 14767 29331 14773
rect 29454 14764 29460 14776
rect 29512 14764 29518 14816
rect 30650 14764 30656 14816
rect 30708 14764 30714 14816
rect 31202 14764 31208 14816
rect 31260 14804 31266 14816
rect 31573 14807 31631 14813
rect 31573 14804 31585 14807
rect 31260 14776 31585 14804
rect 31260 14764 31266 14776
rect 31573 14773 31585 14776
rect 31619 14773 31631 14807
rect 31573 14767 31631 14773
rect 2760 14714 34316 14736
rect 2760 14662 7210 14714
rect 7262 14662 7274 14714
rect 7326 14662 7338 14714
rect 7390 14662 7402 14714
rect 7454 14662 7466 14714
rect 7518 14662 15099 14714
rect 15151 14662 15163 14714
rect 15215 14662 15227 14714
rect 15279 14662 15291 14714
rect 15343 14662 15355 14714
rect 15407 14662 22988 14714
rect 23040 14662 23052 14714
rect 23104 14662 23116 14714
rect 23168 14662 23180 14714
rect 23232 14662 23244 14714
rect 23296 14662 30877 14714
rect 30929 14662 30941 14714
rect 30993 14662 31005 14714
rect 31057 14662 31069 14714
rect 31121 14662 31133 14714
rect 31185 14662 34316 14714
rect 2760 14640 34316 14662
rect 2700 14572 2774 14600
rect 2746 14532 2774 14572
rect 4154 14560 4160 14612
rect 4212 14600 4218 14612
rect 4893 14603 4951 14609
rect 4893 14600 4905 14603
rect 4212 14572 4905 14600
rect 4212 14560 4218 14572
rect 4893 14569 4905 14572
rect 4939 14600 4951 14603
rect 6641 14603 6699 14609
rect 4939 14572 5120 14600
rect 4939 14569 4951 14572
rect 4893 14563 4951 14569
rect 3329 14535 3387 14541
rect 3329 14532 3341 14535
rect 2746 14504 3341 14532
rect 3329 14501 3341 14504
rect 3375 14501 3387 14535
rect 4982 14532 4988 14544
rect 4554 14504 4988 14532
rect 3329 14495 3387 14501
rect 4982 14492 4988 14504
rect 5040 14492 5046 14544
rect 5092 14532 5120 14572
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 7098 14600 7104 14612
rect 6687 14572 7104 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7742 14560 7748 14612
rect 7800 14560 7806 14612
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 10134 14600 10140 14612
rect 8904 14572 10140 14600
rect 8904 14560 8910 14572
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 13630 14560 13636 14612
rect 13688 14600 13694 14612
rect 13909 14603 13967 14609
rect 13909 14600 13921 14603
rect 13688 14572 13921 14600
rect 13688 14560 13694 14572
rect 13909 14569 13921 14572
rect 13955 14569 13967 14603
rect 13909 14563 13967 14569
rect 14458 14560 14464 14612
rect 14516 14560 14522 14612
rect 15194 14560 15200 14612
rect 15252 14560 15258 14612
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15838 14600 15844 14612
rect 15611 14572 15844 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15838 14560 15844 14572
rect 15896 14560 15902 14612
rect 16390 14560 16396 14612
rect 16448 14600 16454 14612
rect 17126 14600 17132 14612
rect 16448 14572 17132 14600
rect 16448 14560 16454 14572
rect 17126 14560 17132 14572
rect 17184 14560 17190 14612
rect 17310 14560 17316 14612
rect 17368 14560 17374 14612
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 17460 14572 17908 14600
rect 17460 14560 17466 14572
rect 5905 14535 5963 14541
rect 5905 14532 5917 14535
rect 5092 14504 5917 14532
rect 5905 14501 5917 14504
rect 5951 14501 5963 14535
rect 5905 14495 5963 14501
rect 5997 14535 6055 14541
rect 5997 14501 6009 14535
rect 6043 14532 6055 14535
rect 10042 14532 10048 14544
rect 6043 14504 6132 14532
rect 9798 14504 10048 14532
rect 6043 14501 6055 14504
rect 5997 14495 6055 14501
rect 3050 14424 3056 14476
rect 3108 14424 3114 14476
rect 5810 14424 5816 14476
rect 5868 14424 5874 14476
rect 5442 14356 5448 14408
rect 5500 14356 5506 14408
rect 4430 14288 4436 14340
rect 4488 14328 4494 14340
rect 4801 14331 4859 14337
rect 4801 14328 4813 14331
rect 4488 14300 4813 14328
rect 4488 14288 4494 14300
rect 4801 14297 4813 14300
rect 4847 14297 4859 14331
rect 6104 14328 6132 14504
rect 10042 14492 10048 14504
rect 10100 14492 10106 14544
rect 6181 14467 6239 14473
rect 6181 14433 6193 14467
rect 6227 14464 6239 14467
rect 6822 14464 6828 14476
rect 6227 14436 6828 14464
rect 6227 14433 6239 14436
rect 6181 14427 6239 14433
rect 6822 14424 6828 14436
rect 6880 14424 6886 14476
rect 7466 14424 7472 14476
rect 7524 14464 7530 14476
rect 8018 14464 8024 14476
rect 7524 14436 8024 14464
rect 7524 14424 7530 14436
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14433 8263 14467
rect 8205 14427 8263 14433
rect 4801 14291 4859 14297
rect 5920 14300 6132 14328
rect 6273 14331 6331 14337
rect 5920 14272 5948 14300
rect 6273 14297 6285 14331
rect 6319 14328 6331 14331
rect 6362 14328 6368 14340
rect 6319 14300 6368 14328
rect 6319 14297 6331 14300
rect 6273 14291 6331 14297
rect 6362 14288 6368 14300
rect 6420 14288 6426 14340
rect 6454 14288 6460 14340
rect 6512 14328 6518 14340
rect 6825 14331 6883 14337
rect 6825 14328 6837 14331
rect 6512 14300 6837 14328
rect 6512 14288 6518 14300
rect 6825 14297 6837 14300
rect 6871 14297 6883 14331
rect 8220 14328 8248 14427
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8573 14399 8631 14405
rect 8343 14368 8432 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8220 14300 8340 14328
rect 6825 14291 6883 14297
rect 8312 14272 8340 14300
rect 5626 14220 5632 14272
rect 5684 14220 5690 14272
rect 5902 14220 5908 14272
rect 5960 14220 5966 14272
rect 6641 14263 6699 14269
rect 6641 14229 6653 14263
rect 6687 14260 6699 14263
rect 7466 14260 7472 14272
rect 6687 14232 7472 14260
rect 6687 14229 6699 14232
rect 6641 14223 6699 14229
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 8113 14263 8171 14269
rect 8113 14229 8125 14263
rect 8159 14260 8171 14263
rect 8202 14260 8208 14272
rect 8159 14232 8208 14260
rect 8159 14229 8171 14232
rect 8113 14223 8171 14229
rect 8202 14220 8208 14232
rect 8260 14220 8266 14272
rect 8294 14220 8300 14272
rect 8352 14220 8358 14272
rect 8404 14260 8432 14368
rect 8573 14365 8585 14399
rect 8619 14396 8631 14399
rect 9122 14396 9128 14408
rect 8619 14368 9128 14396
rect 8619 14365 8631 14368
rect 8573 14359 8631 14365
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 10045 14399 10103 14405
rect 10045 14365 10057 14399
rect 10091 14396 10103 14399
rect 10152 14396 10180 14560
rect 11422 14492 11428 14544
rect 11480 14492 11486 14544
rect 13262 14424 13268 14476
rect 13320 14424 13326 14476
rect 13817 14467 13875 14473
rect 13817 14433 13829 14467
rect 13863 14464 13875 14467
rect 14185 14467 14243 14473
rect 14185 14464 14197 14467
rect 13863 14436 14197 14464
rect 13863 14433 13875 14436
rect 13817 14427 13875 14433
rect 14185 14433 14197 14436
rect 14231 14433 14243 14467
rect 14185 14427 14243 14433
rect 10091 14368 10180 14396
rect 10091 14365 10103 14368
rect 10045 14359 10103 14365
rect 10226 14356 10232 14408
rect 10284 14396 10290 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 10284 14368 10425 14396
rect 10284 14356 10290 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 10686 14356 10692 14408
rect 10744 14356 10750 14408
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12207 14368 12265 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 13906 14356 13912 14408
rect 13964 14356 13970 14408
rect 14093 14399 14151 14405
rect 14093 14365 14105 14399
rect 14139 14396 14151 14399
rect 14476 14396 14504 14560
rect 15212 14532 15240 14560
rect 16114 14532 16120 14544
rect 15212 14504 16120 14532
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 17328 14532 17356 14560
rect 17880 14532 17908 14572
rect 17954 14560 17960 14612
rect 18012 14600 18018 14612
rect 19886 14600 19892 14612
rect 18012 14572 19892 14600
rect 18012 14560 18018 14572
rect 19886 14560 19892 14572
rect 19944 14560 19950 14612
rect 20346 14560 20352 14612
rect 20404 14600 20410 14612
rect 22186 14600 22192 14612
rect 20404 14572 22192 14600
rect 20404 14560 20410 14572
rect 22186 14560 22192 14572
rect 22244 14560 22250 14612
rect 22462 14560 22468 14612
rect 22520 14600 22526 14612
rect 22649 14603 22707 14609
rect 22649 14600 22661 14603
rect 22520 14572 22661 14600
rect 22520 14560 22526 14572
rect 22649 14569 22661 14572
rect 22695 14569 22707 14603
rect 22649 14563 22707 14569
rect 24026 14560 24032 14612
rect 24084 14560 24090 14612
rect 24670 14560 24676 14612
rect 24728 14600 24734 14612
rect 24765 14603 24823 14609
rect 24765 14600 24777 14603
rect 24728 14572 24777 14600
rect 24728 14560 24734 14572
rect 24765 14569 24777 14572
rect 24811 14569 24823 14603
rect 24765 14563 24823 14569
rect 25593 14603 25651 14609
rect 25593 14569 25605 14603
rect 25639 14600 25651 14603
rect 26418 14600 26424 14612
rect 25639 14572 26424 14600
rect 25639 14569 25651 14572
rect 25593 14563 25651 14569
rect 26418 14560 26424 14572
rect 26476 14560 26482 14612
rect 26694 14560 26700 14612
rect 26752 14560 26758 14612
rect 27338 14560 27344 14612
rect 27396 14600 27402 14612
rect 27709 14603 27767 14609
rect 27709 14600 27721 14603
rect 27396 14572 27721 14600
rect 27396 14560 27402 14572
rect 27709 14569 27721 14572
rect 27755 14569 27767 14603
rect 27709 14563 27767 14569
rect 29733 14603 29791 14609
rect 29733 14569 29745 14603
rect 29779 14569 29791 14603
rect 29733 14563 29791 14569
rect 18690 14532 18696 14544
rect 17328 14504 17632 14532
rect 17880 14504 18696 14532
rect 14918 14424 14924 14476
rect 14976 14464 14982 14476
rect 15013 14467 15071 14473
rect 15013 14464 15025 14467
rect 14976 14436 15025 14464
rect 14976 14424 14982 14436
rect 15013 14433 15025 14436
rect 15059 14433 15071 14467
rect 15013 14427 15071 14433
rect 15930 14424 15936 14476
rect 15988 14464 15994 14476
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 15988 14436 16313 14464
rect 15988 14424 15994 14436
rect 16301 14433 16313 14436
rect 16347 14464 16359 14467
rect 16393 14467 16451 14473
rect 16393 14464 16405 14467
rect 16347 14436 16405 14464
rect 16347 14433 16359 14436
rect 16301 14427 16359 14433
rect 16393 14433 16405 14436
rect 16439 14464 16451 14467
rect 16482 14464 16488 14476
rect 16439 14436 16488 14464
rect 16439 14433 16451 14436
rect 16393 14427 16451 14433
rect 16482 14424 16488 14436
rect 16540 14424 16546 14476
rect 17494 14424 17500 14476
rect 17552 14424 17558 14476
rect 17604 14473 17632 14504
rect 18690 14492 18696 14504
rect 18748 14492 18754 14544
rect 18782 14492 18788 14544
rect 18840 14532 18846 14544
rect 18840 14504 18906 14532
rect 18840 14492 18846 14504
rect 20070 14492 20076 14544
rect 20128 14532 20134 14544
rect 21174 14532 21180 14544
rect 20128 14504 20392 14532
rect 20128 14492 20134 14504
rect 17589 14467 17647 14473
rect 17589 14433 17601 14467
rect 17635 14433 17647 14467
rect 17589 14427 17647 14433
rect 17770 14424 17776 14476
rect 17828 14424 17834 14476
rect 17862 14424 17868 14476
rect 17920 14424 17926 14476
rect 20364 14464 20392 14504
rect 20824 14504 21180 14532
rect 20441 14467 20499 14473
rect 20441 14464 20453 14467
rect 20364 14436 20453 14464
rect 20441 14433 20453 14436
rect 20487 14433 20499 14467
rect 20441 14427 20499 14433
rect 20530 14424 20536 14476
rect 20588 14424 20594 14476
rect 20824 14473 20852 14504
rect 21174 14492 21180 14504
rect 21232 14492 21238 14544
rect 22833 14535 22891 14541
rect 22833 14532 22845 14535
rect 22402 14504 22845 14532
rect 22833 14501 22845 14504
rect 22879 14501 22891 14535
rect 22833 14495 22891 14501
rect 26050 14492 26056 14544
rect 26108 14532 26114 14544
rect 26191 14535 26249 14541
rect 26191 14532 26203 14535
rect 26108 14504 26203 14532
rect 26108 14492 26114 14504
rect 26191 14501 26203 14504
rect 26237 14501 26249 14535
rect 27982 14532 27988 14544
rect 26191 14495 26249 14501
rect 26620 14504 27988 14532
rect 20809 14467 20867 14473
rect 20809 14433 20821 14467
rect 20855 14433 20867 14467
rect 20809 14427 20867 14433
rect 22462 14424 22468 14476
rect 22520 14424 22526 14476
rect 22646 14424 22652 14476
rect 22704 14424 22710 14476
rect 22925 14467 22983 14473
rect 22925 14433 22937 14467
rect 22971 14464 22983 14467
rect 23750 14464 23756 14476
rect 22971 14436 23756 14464
rect 22971 14433 22983 14436
rect 22925 14427 22983 14433
rect 23750 14424 23756 14436
rect 23808 14464 23814 14476
rect 24857 14467 24915 14473
rect 24857 14464 24869 14467
rect 23808 14436 24869 14464
rect 23808 14424 23814 14436
rect 24857 14433 24869 14436
rect 24903 14464 24915 14467
rect 24946 14464 24952 14476
rect 24903 14436 24952 14464
rect 24903 14433 24915 14436
rect 24857 14427 24915 14433
rect 24946 14424 24952 14436
rect 25004 14424 25010 14476
rect 25774 14424 25780 14476
rect 25832 14424 25838 14476
rect 25958 14424 25964 14476
rect 26016 14424 26022 14476
rect 26329 14467 26387 14473
rect 26329 14433 26341 14467
rect 26375 14433 26387 14467
rect 26329 14427 26387 14433
rect 14139 14368 14504 14396
rect 14553 14399 14611 14405
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 10244 14328 10272 14356
rect 9600 14300 10272 14328
rect 13924 14328 13952 14356
rect 14568 14328 14596 14359
rect 14734 14356 14740 14408
rect 14792 14396 14798 14408
rect 16114 14396 16120 14408
rect 14792 14368 16120 14396
rect 14792 14356 14798 14368
rect 16114 14356 16120 14368
rect 16172 14396 16178 14408
rect 16669 14399 16727 14405
rect 16669 14396 16681 14399
rect 16172 14368 16681 14396
rect 16172 14356 16178 14368
rect 16669 14365 16681 14368
rect 16715 14396 16727 14399
rect 17313 14399 17371 14405
rect 16715 14368 17264 14396
rect 16715 14365 16727 14368
rect 16669 14359 16727 14365
rect 17236 14340 17264 14368
rect 17313 14365 17325 14399
rect 17359 14396 17371 14399
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 17359 14368 20085 14396
rect 17359 14365 17371 14368
rect 17313 14359 17371 14365
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 20073 14359 20131 14365
rect 20349 14399 20407 14405
rect 20349 14365 20361 14399
rect 20395 14365 20407 14399
rect 20349 14359 20407 14365
rect 20901 14399 20959 14405
rect 20901 14365 20913 14399
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 13924 14300 14596 14328
rect 14752 14300 17080 14328
rect 9600 14260 9628 14300
rect 8404 14232 9628 14260
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 12860 14232 12909 14260
rect 12860 14220 12866 14232
rect 12897 14229 12909 14232
rect 12943 14229 12955 14263
rect 12897 14223 12955 14229
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 14752 14260 14780 14300
rect 14148 14232 14780 14260
rect 14829 14263 14887 14269
rect 14148 14220 14154 14232
rect 14829 14229 14841 14263
rect 14875 14260 14887 14263
rect 14918 14260 14924 14272
rect 14875 14232 14924 14260
rect 14875 14229 14887 14232
rect 14829 14223 14887 14229
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 15654 14220 15660 14272
rect 15712 14220 15718 14272
rect 17052 14260 17080 14300
rect 17218 14288 17224 14340
rect 17276 14288 17282 14340
rect 18322 14328 18328 14340
rect 17972 14300 18328 14328
rect 17972 14260 18000 14300
rect 18322 14288 18328 14300
rect 18380 14288 18386 14340
rect 18874 14328 18880 14340
rect 18616 14300 18880 14328
rect 17052 14232 18000 14260
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 18616 14269 18644 14300
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 20364 14328 20392 14359
rect 20916 14328 20944 14359
rect 21174 14356 21180 14408
rect 21232 14356 21238 14408
rect 21266 14356 21272 14408
rect 21324 14396 21330 14408
rect 22480 14396 22508 14424
rect 21324 14368 22508 14396
rect 22664 14396 22692 14424
rect 23198 14396 23204 14408
rect 22664 14368 23204 14396
rect 21324 14356 21330 14368
rect 23198 14356 23204 14368
rect 23256 14356 23262 14408
rect 23382 14356 23388 14408
rect 23440 14396 23446 14408
rect 26053 14399 26111 14405
rect 26053 14396 26065 14399
rect 23440 14368 26065 14396
rect 23440 14356 23446 14368
rect 26053 14365 26065 14368
rect 26099 14365 26111 14399
rect 26344 14396 26372 14427
rect 26418 14424 26424 14476
rect 26476 14424 26482 14476
rect 26513 14467 26571 14473
rect 26513 14433 26525 14467
rect 26559 14464 26571 14467
rect 26620 14464 26648 14504
rect 27982 14492 27988 14504
rect 28040 14532 28046 14544
rect 28445 14535 28503 14541
rect 28445 14532 28457 14535
rect 28040 14504 28457 14532
rect 28040 14492 28046 14504
rect 28445 14501 28457 14504
rect 28491 14501 28503 14535
rect 28445 14495 28503 14501
rect 28994 14492 29000 14544
rect 29052 14532 29058 14544
rect 29365 14535 29423 14541
rect 29365 14532 29377 14535
rect 29052 14504 29377 14532
rect 29052 14492 29058 14504
rect 29365 14501 29377 14504
rect 29411 14501 29423 14535
rect 29748 14532 29776 14563
rect 29822 14560 29828 14612
rect 29880 14560 29886 14612
rect 30006 14560 30012 14612
rect 30064 14560 30070 14612
rect 30650 14560 30656 14612
rect 30708 14600 30714 14612
rect 30708 14572 31340 14600
rect 30708 14560 30714 14572
rect 30024 14532 30052 14560
rect 31202 14532 31208 14544
rect 29748 14504 30052 14532
rect 30866 14504 31208 14532
rect 29365 14495 29423 14501
rect 31202 14492 31208 14504
rect 31260 14492 31266 14544
rect 31312 14541 31340 14572
rect 31297 14535 31355 14541
rect 31297 14501 31309 14535
rect 31343 14501 31355 14535
rect 31297 14495 31355 14501
rect 26559 14436 26648 14464
rect 26559 14433 26571 14436
rect 26513 14427 26571 14433
rect 26694 14424 26700 14476
rect 26752 14464 26758 14476
rect 27801 14467 27859 14473
rect 27801 14464 27813 14467
rect 26752 14436 27813 14464
rect 26752 14424 26758 14436
rect 27801 14433 27813 14436
rect 27847 14433 27859 14467
rect 27801 14427 27859 14433
rect 28626 14424 28632 14476
rect 28684 14464 28690 14476
rect 29089 14467 29147 14473
rect 29089 14464 29101 14467
rect 28684 14436 29101 14464
rect 28684 14424 28690 14436
rect 29089 14433 29101 14436
rect 29135 14433 29147 14467
rect 29089 14427 29147 14433
rect 29178 14424 29184 14476
rect 29236 14424 29242 14476
rect 29454 14424 29460 14476
rect 29512 14424 29518 14476
rect 29549 14467 29607 14473
rect 29549 14433 29561 14467
rect 29595 14464 29607 14467
rect 29822 14464 29828 14476
rect 29595 14436 29828 14464
rect 29595 14433 29607 14436
rect 29549 14427 29607 14433
rect 29822 14424 29828 14436
rect 29880 14424 29886 14476
rect 31573 14467 31631 14473
rect 31573 14433 31585 14467
rect 31619 14464 31631 14467
rect 31846 14464 31852 14476
rect 31619 14436 31852 14464
rect 31619 14433 31631 14436
rect 31573 14427 31631 14433
rect 31846 14424 31852 14436
rect 31904 14464 31910 14476
rect 32306 14464 32312 14476
rect 31904 14436 32312 14464
rect 31904 14424 31910 14436
rect 32306 14424 32312 14436
rect 32364 14424 32370 14476
rect 32769 14467 32827 14473
rect 32769 14433 32781 14467
rect 32815 14433 32827 14467
rect 32769 14427 32827 14433
rect 26344 14368 26924 14396
rect 26053 14359 26111 14365
rect 26896 14340 26924 14368
rect 27062 14356 27068 14408
rect 27120 14356 27126 14408
rect 29472 14396 29500 14424
rect 32784 14396 32812 14427
rect 29472 14368 32812 14396
rect 32858 14356 32864 14408
rect 32916 14356 32922 14408
rect 33045 14399 33103 14405
rect 33045 14365 33057 14399
rect 33091 14396 33103 14399
rect 33686 14396 33692 14408
rect 33091 14368 33692 14396
rect 33091 14365 33103 14368
rect 33045 14359 33103 14365
rect 20364 14300 20944 14328
rect 18601 14263 18659 14269
rect 18601 14260 18613 14263
rect 18104 14232 18613 14260
rect 18104 14220 18110 14232
rect 18601 14229 18613 14232
rect 18647 14229 18659 14263
rect 18601 14223 18659 14229
rect 18690 14220 18696 14272
rect 18748 14260 18754 14272
rect 20530 14260 20536 14272
rect 18748 14232 20536 14260
rect 18748 14220 18754 14232
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 20916 14260 20944 14300
rect 22278 14288 22284 14340
rect 22336 14328 22342 14340
rect 24486 14328 24492 14340
rect 22336 14300 24492 14328
rect 22336 14288 22342 14300
rect 24486 14288 24492 14300
rect 24544 14288 24550 14340
rect 26878 14288 26884 14340
rect 26936 14328 26942 14340
rect 28810 14328 28816 14340
rect 26936 14300 28816 14328
rect 26936 14288 26942 14300
rect 28810 14288 28816 14300
rect 28868 14328 28874 14340
rect 30006 14328 30012 14340
rect 28868 14300 30012 14328
rect 28868 14288 28874 14300
rect 30006 14288 30012 14300
rect 30064 14288 30070 14340
rect 33520 14272 33548 14368
rect 33686 14356 33692 14368
rect 33744 14356 33750 14408
rect 22186 14260 22192 14272
rect 20916 14232 22192 14260
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 22922 14220 22928 14272
rect 22980 14260 22986 14272
rect 23201 14263 23259 14269
rect 23201 14260 23213 14263
rect 22980 14232 23213 14260
rect 22980 14220 22986 14232
rect 23201 14229 23213 14232
rect 23247 14229 23259 14263
rect 23201 14223 23259 14229
rect 23382 14220 23388 14272
rect 23440 14260 23446 14272
rect 23661 14263 23719 14269
rect 23661 14260 23673 14263
rect 23440 14232 23673 14260
rect 23440 14220 23446 14232
rect 23661 14229 23673 14232
rect 23707 14229 23719 14263
rect 23661 14223 23719 14229
rect 26418 14220 26424 14272
rect 26476 14260 26482 14272
rect 26786 14260 26792 14272
rect 26476 14232 26792 14260
rect 26476 14220 26482 14232
rect 26786 14220 26792 14232
rect 26844 14260 26850 14272
rect 28902 14260 28908 14272
rect 26844 14232 28908 14260
rect 26844 14220 26850 14232
rect 28902 14220 28908 14232
rect 28960 14220 28966 14272
rect 28994 14220 29000 14272
rect 29052 14220 29058 14272
rect 32398 14220 32404 14272
rect 32456 14220 32462 14272
rect 33502 14220 33508 14272
rect 33560 14220 33566 14272
rect 2760 14170 34316 14192
rect 2760 14118 6550 14170
rect 6602 14118 6614 14170
rect 6666 14118 6678 14170
rect 6730 14118 6742 14170
rect 6794 14118 6806 14170
rect 6858 14118 14439 14170
rect 14491 14118 14503 14170
rect 14555 14118 14567 14170
rect 14619 14118 14631 14170
rect 14683 14118 14695 14170
rect 14747 14118 22328 14170
rect 22380 14118 22392 14170
rect 22444 14118 22456 14170
rect 22508 14118 22520 14170
rect 22572 14118 22584 14170
rect 22636 14118 30217 14170
rect 30269 14118 30281 14170
rect 30333 14118 30345 14170
rect 30397 14118 30409 14170
rect 30461 14118 30473 14170
rect 30525 14118 34316 14170
rect 2760 14096 34316 14118
rect 4522 14016 4528 14068
rect 4580 14056 4586 14068
rect 4706 14056 4712 14068
rect 4580 14028 4712 14056
rect 4580 14016 4586 14028
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 4982 14016 4988 14068
rect 5040 14016 5046 14068
rect 5626 14016 5632 14068
rect 5684 14016 5690 14068
rect 5810 14016 5816 14068
rect 5868 14056 5874 14068
rect 6178 14056 6184 14068
rect 5868 14028 6184 14056
rect 5868 14016 5874 14028
rect 6178 14016 6184 14028
rect 6236 14056 6242 14068
rect 6825 14059 6883 14065
rect 6825 14056 6837 14059
rect 6236 14028 6837 14056
rect 6236 14016 6242 14028
rect 6825 14025 6837 14028
rect 6871 14056 6883 14059
rect 6871 14028 8248 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 1302 13880 1308 13932
rect 1360 13920 1366 13932
rect 3237 13923 3295 13929
rect 3237 13920 3249 13923
rect 1360 13892 3249 13920
rect 1360 13880 1366 13892
rect 3237 13889 3249 13892
rect 3283 13889 3295 13923
rect 5644 13920 5672 14016
rect 6914 13948 6920 14000
rect 6972 13948 6978 14000
rect 8220 13988 8248 14028
rect 8662 14016 8668 14068
rect 8720 14016 8726 14068
rect 9122 14016 9128 14068
rect 9180 14016 9186 14068
rect 9766 14016 9772 14068
rect 9824 14016 9830 14068
rect 10042 14016 10048 14068
rect 10100 14016 10106 14068
rect 10686 14016 10692 14068
rect 10744 14056 10750 14068
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 10744 14028 11069 14056
rect 10744 14016 10750 14028
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 11057 14019 11115 14025
rect 12526 14016 12532 14068
rect 12584 14056 12590 14068
rect 13633 14059 13691 14065
rect 12584 14028 13124 14056
rect 12584 14016 12590 14028
rect 8938 13988 8944 14000
rect 8220 13960 8944 13988
rect 8938 13948 8944 13960
rect 8996 13948 9002 14000
rect 9784 13988 9812 14016
rect 12802 13988 12808 14000
rect 9600 13960 9812 13988
rect 11532 13960 12808 13988
rect 5813 13923 5871 13929
rect 5813 13920 5825 13923
rect 5644 13892 5825 13920
rect 3237 13883 3295 13889
rect 5813 13889 5825 13892
rect 5859 13889 5871 13923
rect 6932 13920 6960 13948
rect 9600 13929 9628 13960
rect 11532 13929 11560 13960
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 12894 13948 12900 14000
rect 12952 13948 12958 14000
rect 13096 13988 13124 14028
rect 13633 14025 13645 14059
rect 13679 14056 13691 14059
rect 13814 14056 13820 14068
rect 13679 14028 13820 14056
rect 13679 14025 13691 14028
rect 13633 14019 13691 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14332 14028 14749 14056
rect 14332 14016 14338 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 15562 14056 15568 14068
rect 14737 14019 14795 14025
rect 15028 14028 15568 14056
rect 13722 13988 13728 14000
rect 13096 13960 13728 13988
rect 13722 13948 13728 13960
rect 13780 13988 13786 14000
rect 14185 13991 14243 13997
rect 14185 13988 14197 13991
rect 13780 13960 14197 13988
rect 13780 13948 13786 13960
rect 14185 13957 14197 13960
rect 14231 13957 14243 13991
rect 14185 13951 14243 13957
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 6932 13892 7205 13920
rect 5813 13883 5871 13889
rect 7193 13889 7205 13892
rect 7239 13889 7251 13923
rect 7193 13883 7251 13889
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 9723 13892 10793 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13821 4491 13855
rect 4433 13815 4491 13821
rect 5077 13855 5135 13861
rect 5077 13821 5089 13855
rect 5123 13852 5135 13855
rect 5166 13852 5172 13864
rect 5123 13824 5172 13852
rect 5123 13821 5135 13824
rect 5077 13815 5135 13821
rect 4448 13784 4476 13815
rect 5166 13812 5172 13824
rect 5224 13852 5230 13864
rect 5629 13855 5687 13861
rect 5629 13852 5641 13855
rect 5224 13824 5641 13852
rect 5224 13812 5230 13824
rect 5629 13821 5641 13824
rect 5675 13821 5687 13855
rect 5629 13815 5687 13821
rect 6362 13812 6368 13864
rect 6420 13852 6426 13864
rect 6917 13855 6975 13861
rect 6917 13852 6929 13855
rect 6420 13824 6929 13852
rect 6420 13812 6426 13824
rect 6917 13821 6929 13824
rect 6963 13821 6975 13855
rect 6917 13815 6975 13821
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 8260 13824 8326 13852
rect 8260 13812 8266 13824
rect 8662 13812 8668 13864
rect 8720 13852 8726 13864
rect 9692 13852 9720 13883
rect 11698 13880 11704 13932
rect 11756 13920 11762 13932
rect 12618 13920 12624 13932
rect 11756 13892 12624 13920
rect 11756 13880 11762 13892
rect 12618 13880 12624 13892
rect 12676 13880 12682 13932
rect 12820 13920 12848 13948
rect 13170 13920 13176 13932
rect 12820 13892 13176 13920
rect 13170 13880 13176 13892
rect 13228 13920 13234 13932
rect 13449 13923 13507 13929
rect 13449 13920 13461 13923
rect 13228 13892 13461 13920
rect 13228 13880 13234 13892
rect 13449 13889 13461 13892
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 14090 13880 14096 13932
rect 14148 13920 14154 13932
rect 15028 13920 15056 14028
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 16114 14056 16120 14068
rect 15672 14028 16120 14056
rect 15672 13988 15700 14028
rect 16114 14016 16120 14028
rect 16172 14016 16178 14068
rect 16853 14059 16911 14065
rect 16408 14028 16804 14056
rect 15396 13960 15700 13988
rect 15749 13991 15807 13997
rect 15396 13929 15424 13960
rect 15749 13957 15761 13991
rect 15795 13988 15807 13991
rect 16022 13988 16028 14000
rect 15795 13960 16028 13988
rect 15795 13957 15807 13960
rect 15749 13951 15807 13957
rect 16022 13948 16028 13960
rect 16080 13948 16086 14000
rect 16298 13948 16304 14000
rect 16356 13948 16362 14000
rect 14148 13892 14412 13920
rect 14148 13880 14154 13892
rect 8720 13824 9720 13852
rect 8720 13812 8726 13824
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 10137 13855 10195 13861
rect 10137 13852 10149 13855
rect 10100 13824 10149 13852
rect 10100 13812 10106 13824
rect 10137 13821 10149 13824
rect 10183 13852 10195 13855
rect 10183 13824 10272 13852
rect 10183 13821 10195 13824
rect 10137 13815 10195 13821
rect 4448 13756 6592 13784
rect 5534 13676 5540 13728
rect 5592 13676 5598 13728
rect 6454 13676 6460 13728
rect 6512 13676 6518 13728
rect 6564 13716 6592 13756
rect 8846 13744 8852 13796
rect 8904 13744 8910 13796
rect 9493 13787 9551 13793
rect 9493 13753 9505 13787
rect 9539 13784 9551 13787
rect 9950 13784 9956 13796
rect 9539 13756 9956 13784
rect 9539 13753 9551 13756
rect 9493 13747 9551 13753
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 10244 13784 10272 13824
rect 10318 13812 10324 13864
rect 10376 13852 10382 13864
rect 11885 13855 11943 13861
rect 11885 13852 11897 13855
rect 10376 13824 11897 13852
rect 10376 13812 10382 13824
rect 11885 13821 11897 13824
rect 11931 13821 11943 13855
rect 11885 13815 11943 13821
rect 12342 13812 12348 13864
rect 12400 13812 12406 13864
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13852 12587 13855
rect 13262 13852 13268 13864
rect 12575 13824 13268 13852
rect 12575 13821 12587 13824
rect 12529 13815 12587 13821
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 14274 13812 14280 13864
rect 14332 13812 14338 13864
rect 14384 13861 14412 13892
rect 14936 13892 15056 13920
rect 15381 13923 15439 13929
rect 14369 13855 14427 13861
rect 14369 13821 14381 13855
rect 14415 13821 14427 13855
rect 14369 13815 14427 13821
rect 14458 13812 14464 13864
rect 14516 13812 14522 13864
rect 14936 13861 14964 13892
rect 15381 13889 15393 13923
rect 15427 13889 15439 13923
rect 15381 13883 15439 13889
rect 15562 13880 15568 13932
rect 15620 13920 15626 13932
rect 16114 13920 16120 13932
rect 15620 13892 15976 13920
rect 15620 13880 15626 13892
rect 14645 13855 14703 13861
rect 14645 13852 14657 13855
rect 14568 13824 14657 13852
rect 10410 13784 10416 13796
rect 10244 13756 10416 13784
rect 10410 13744 10416 13756
rect 10468 13744 10474 13796
rect 11425 13787 11483 13793
rect 11425 13753 11437 13787
rect 11471 13784 11483 13787
rect 12360 13784 12388 13812
rect 11471 13756 12388 13784
rect 12897 13787 12955 13793
rect 11471 13753 11483 13756
rect 11425 13747 11483 13753
rect 12897 13753 12909 13787
rect 12943 13784 12955 13787
rect 13078 13784 13084 13796
rect 12943 13756 13084 13784
rect 12943 13753 12955 13756
rect 12897 13747 12955 13753
rect 13078 13744 13084 13756
rect 13136 13744 13142 13796
rect 14292 13784 14320 13812
rect 14568 13784 14596 13824
rect 14645 13821 14657 13824
rect 14691 13821 14703 13855
rect 14645 13815 14703 13821
rect 14921 13855 14979 13861
rect 14921 13821 14933 13855
rect 14967 13821 14979 13855
rect 14921 13815 14979 13821
rect 15243 13855 15301 13861
rect 15243 13821 15255 13855
rect 15289 13852 15301 13855
rect 15470 13852 15476 13864
rect 15289 13824 15476 13852
rect 15289 13821 15301 13824
rect 15243 13815 15301 13821
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15746 13812 15752 13864
rect 15804 13812 15810 13864
rect 15948 13861 15976 13892
rect 16040 13892 16120 13920
rect 16040 13861 16068 13892
rect 16114 13880 16120 13892
rect 16172 13920 16178 13932
rect 16316 13920 16344 13948
rect 16408 13929 16436 14028
rect 16776 13988 16804 14028
rect 16853 14025 16865 14059
rect 16899 14056 16911 14059
rect 17034 14056 17040 14068
rect 16899 14028 17040 14056
rect 16899 14025 16911 14028
rect 16853 14019 16911 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 17129 14059 17187 14065
rect 17129 14025 17141 14059
rect 17175 14056 17187 14059
rect 17218 14056 17224 14068
rect 17175 14028 17224 14056
rect 17175 14025 17187 14028
rect 17129 14019 17187 14025
rect 17218 14016 17224 14028
rect 17276 14016 17282 14068
rect 18414 14016 18420 14068
rect 18472 14016 18478 14068
rect 18782 14016 18788 14068
rect 18840 14016 18846 14068
rect 19058 14016 19064 14068
rect 19116 14056 19122 14068
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19116 14028 19901 14056
rect 19116 14016 19122 14028
rect 19889 14025 19901 14028
rect 19935 14056 19947 14059
rect 20162 14056 20168 14068
rect 19935 14028 20168 14056
rect 19935 14025 19947 14028
rect 19889 14019 19947 14025
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20530 14056 20536 14068
rect 20404 14028 20536 14056
rect 20404 14016 20410 14028
rect 20530 14016 20536 14028
rect 20588 14016 20594 14068
rect 21542 14056 21548 14068
rect 20640 14028 21548 14056
rect 16776 13960 17080 13988
rect 16172 13892 16344 13920
rect 16393 13923 16451 13929
rect 16172 13880 16178 13892
rect 16393 13889 16405 13923
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 16758 13886 16764 13932
rect 16687 13880 16764 13886
rect 16816 13880 16822 13932
rect 16942 13880 16948 13932
rect 17000 13880 17006 13932
rect 16687 13861 16804 13880
rect 15933 13855 15991 13861
rect 15933 13821 15945 13855
rect 15979 13821 15991 13855
rect 15933 13815 15991 13821
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13821 16083 13855
rect 16484 13855 16542 13861
rect 16484 13852 16496 13855
rect 16025 13815 16083 13821
rect 16132 13824 16496 13852
rect 13188 13756 14044 13784
rect 14292 13756 14596 13784
rect 8864 13716 8892 13744
rect 6564 13688 8892 13716
rect 9858 13676 9864 13728
rect 9916 13716 9922 13728
rect 13188 13716 13216 13756
rect 9916 13688 13216 13716
rect 9916 13676 9922 13688
rect 13354 13676 13360 13728
rect 13412 13676 13418 13728
rect 14016 13725 14044 13756
rect 15010 13744 15016 13796
rect 15068 13744 15074 13796
rect 15105 13787 15163 13793
rect 15105 13753 15117 13787
rect 15151 13784 15163 13787
rect 15838 13784 15844 13796
rect 15151 13756 15844 13784
rect 15151 13753 15163 13756
rect 15105 13747 15163 13753
rect 15838 13744 15844 13756
rect 15896 13784 15902 13796
rect 16132 13784 16160 13824
rect 16484 13821 16496 13824
rect 16530 13821 16542 13855
rect 16484 13815 16542 13821
rect 16577 13855 16635 13861
rect 16577 13821 16589 13855
rect 16623 13821 16635 13855
rect 16577 13815 16635 13821
rect 16669 13858 16804 13861
rect 16669 13855 16727 13858
rect 16669 13821 16681 13855
rect 16715 13821 16727 13855
rect 16960 13852 16988 13880
rect 16669 13815 16727 13821
rect 16868 13824 16988 13852
rect 16868 13818 16896 13824
rect 15896 13756 16160 13784
rect 16592 13784 16620 13815
rect 16776 13790 16896 13818
rect 16776 13784 16804 13790
rect 16592 13756 16804 13784
rect 15896 13744 15902 13756
rect 14001 13719 14059 13725
rect 14001 13685 14013 13719
rect 14047 13716 14059 13719
rect 14458 13716 14464 13728
rect 14047 13688 14464 13716
rect 14047 13685 14059 13688
rect 14001 13679 14059 13685
rect 14458 13676 14464 13688
rect 14516 13676 14522 13728
rect 14553 13719 14611 13725
rect 14553 13685 14565 13719
rect 14599 13716 14611 13719
rect 16482 13716 16488 13728
rect 14599 13688 16488 13716
rect 14599 13685 14611 13688
rect 14553 13679 14611 13685
rect 16482 13676 16488 13688
rect 16540 13676 16546 13728
rect 16850 13676 16856 13728
rect 16908 13716 16914 13728
rect 16945 13719 17003 13725
rect 16945 13716 16957 13719
rect 16908 13688 16957 13716
rect 16908 13676 16914 13688
rect 16945 13685 16957 13688
rect 16991 13716 17003 13719
rect 17052 13716 17080 13960
rect 17402 13948 17408 14000
rect 17460 13988 17466 14000
rect 17497 13991 17555 13997
rect 17497 13988 17509 13991
rect 17460 13960 17509 13988
rect 17460 13948 17466 13960
rect 17497 13957 17509 13960
rect 17543 13957 17555 13991
rect 18432 13988 18460 14016
rect 19242 13988 19248 14000
rect 18432 13960 19248 13988
rect 17497 13951 17555 13957
rect 19242 13948 19248 13960
rect 19300 13948 19306 14000
rect 19260 13920 19288 13948
rect 20640 13920 20668 14028
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 22281 14059 22339 14065
rect 22281 14025 22293 14059
rect 22327 14056 22339 14059
rect 22327 14028 24440 14056
rect 22327 14025 22339 14028
rect 22281 14019 22339 14025
rect 22094 13948 22100 14000
rect 22152 13988 22158 14000
rect 22370 13988 22376 14000
rect 22152 13960 22376 13988
rect 22152 13948 22158 13960
rect 22370 13948 22376 13960
rect 22428 13948 22434 14000
rect 19260 13892 20668 13920
rect 21191 13892 22048 13920
rect 17586 13812 17592 13864
rect 17644 13852 17650 13864
rect 17773 13855 17831 13861
rect 17773 13852 17785 13855
rect 17644 13824 17785 13852
rect 17644 13812 17650 13824
rect 17773 13821 17785 13824
rect 17819 13821 17831 13855
rect 17773 13815 17831 13821
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18693 13855 18751 13861
rect 18003 13824 18368 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18046 13744 18052 13796
rect 18104 13784 18110 13796
rect 18233 13787 18291 13793
rect 18233 13784 18245 13787
rect 18104 13756 18245 13784
rect 18104 13744 18110 13756
rect 18233 13753 18245 13756
rect 18279 13753 18291 13787
rect 18340 13784 18368 13824
rect 18693 13821 18705 13855
rect 18739 13852 18751 13855
rect 19334 13852 19340 13864
rect 18739 13824 19340 13852
rect 18739 13821 18751 13824
rect 18693 13815 18751 13821
rect 19334 13812 19340 13824
rect 19392 13852 19398 13864
rect 20346 13852 20352 13864
rect 19392 13824 20352 13852
rect 19392 13812 19398 13824
rect 20346 13812 20352 13824
rect 20404 13812 20410 13864
rect 21191 13861 21219 13892
rect 22020 13864 22048 13892
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22922 13920 22928 13932
rect 22336 13892 22928 13920
rect 22336 13880 22342 13892
rect 22922 13880 22928 13892
rect 22980 13880 22986 13932
rect 23084 13923 23142 13929
rect 23084 13889 23096 13923
rect 23130 13920 23142 13923
rect 23382 13920 23388 13932
rect 23130 13892 23388 13920
rect 23130 13889 23142 13892
rect 23084 13883 23142 13889
rect 23382 13880 23388 13892
rect 23440 13880 23446 13932
rect 23474 13880 23480 13932
rect 23532 13880 23538 13932
rect 24210 13920 24216 13932
rect 23952 13892 24216 13920
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13852 20775 13855
rect 20901 13855 20959 13861
rect 20901 13852 20913 13855
rect 20763 13824 20913 13852
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 20901 13821 20913 13824
rect 20947 13821 20959 13855
rect 20901 13815 20959 13821
rect 21176 13855 21234 13861
rect 21176 13821 21188 13855
rect 21222 13821 21234 13855
rect 21176 13815 21234 13821
rect 21266 13812 21272 13864
rect 21324 13812 21330 13864
rect 21545 13855 21603 13861
rect 21545 13821 21557 13855
rect 21591 13821 21603 13855
rect 21545 13815 21603 13821
rect 18506 13784 18512 13796
rect 18340 13756 18512 13784
rect 18233 13747 18291 13753
rect 18506 13744 18512 13756
rect 18564 13784 18570 13796
rect 19058 13784 19064 13796
rect 18564 13756 19064 13784
rect 18564 13744 18570 13756
rect 19058 13744 19064 13756
rect 19116 13744 19122 13796
rect 20806 13744 20812 13796
rect 20864 13784 20870 13796
rect 21560 13784 21588 13815
rect 21634 13812 21640 13864
rect 21692 13812 21698 13864
rect 21821 13855 21879 13861
rect 21821 13852 21833 13855
rect 21744 13824 21833 13852
rect 20864 13756 21588 13784
rect 20864 13744 20870 13756
rect 16991 13688 17080 13716
rect 16991 13685 17003 13688
rect 16945 13679 17003 13685
rect 17126 13676 17132 13728
rect 17184 13716 17190 13728
rect 18141 13719 18199 13725
rect 18141 13716 18153 13719
rect 17184 13688 18153 13716
rect 17184 13676 17190 13688
rect 18141 13685 18153 13688
rect 18187 13716 18199 13719
rect 19150 13716 19156 13728
rect 18187 13688 19156 13716
rect 18187 13685 18199 13688
rect 18141 13679 18199 13685
rect 19150 13676 19156 13688
rect 19208 13676 19214 13728
rect 20070 13676 20076 13728
rect 20128 13676 20134 13728
rect 20438 13676 20444 13728
rect 20496 13716 20502 13728
rect 21744 13716 21772 13824
rect 21821 13821 21833 13824
rect 21867 13821 21879 13855
rect 21821 13815 21879 13821
rect 21913 13855 21971 13861
rect 21913 13821 21925 13855
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 20496 13688 21772 13716
rect 21928 13716 21956 13815
rect 22002 13812 22008 13864
rect 22060 13812 22066 13864
rect 22097 13855 22155 13861
rect 22097 13821 22109 13855
rect 22143 13852 22155 13855
rect 22143 13824 22416 13852
rect 22143 13821 22155 13824
rect 22097 13815 22155 13821
rect 22002 13716 22008 13728
rect 21928 13688 22008 13716
rect 20496 13676 20502 13688
rect 22002 13676 22008 13688
rect 22060 13676 22066 13728
rect 22388 13716 22416 13824
rect 23198 13812 23204 13864
rect 23256 13812 23262 13864
rect 23952 13861 23980 13892
rect 24210 13880 24216 13892
rect 24268 13880 24274 13932
rect 23937 13855 23995 13861
rect 23937 13821 23949 13855
rect 23983 13821 23995 13855
rect 23937 13815 23995 13821
rect 24118 13812 24124 13864
rect 24176 13812 24182 13864
rect 24412 13861 24440 14028
rect 24486 14016 24492 14068
rect 24544 14016 24550 14068
rect 25774 14016 25780 14068
rect 25832 14056 25838 14068
rect 25869 14059 25927 14065
rect 25869 14056 25881 14059
rect 25832 14028 25881 14056
rect 25832 14016 25838 14028
rect 25869 14025 25881 14028
rect 25915 14025 25927 14059
rect 25869 14019 25927 14025
rect 25958 14016 25964 14068
rect 26016 14056 26022 14068
rect 26053 14059 26111 14065
rect 26053 14056 26065 14059
rect 26016 14028 26065 14056
rect 26016 14016 26022 14028
rect 26053 14025 26065 14028
rect 26099 14025 26111 14059
rect 26053 14019 26111 14025
rect 26878 14016 26884 14068
rect 26936 14016 26942 14068
rect 27062 14016 27068 14068
rect 27120 14016 27126 14068
rect 27614 14056 27620 14068
rect 27264 14028 27620 14056
rect 24504 13920 24532 14016
rect 25682 13948 25688 14000
rect 25740 13948 25746 14000
rect 26602 13988 26608 14000
rect 26252 13960 26608 13988
rect 24581 13923 24639 13929
rect 24581 13920 24593 13923
rect 24504 13892 24593 13920
rect 24581 13889 24593 13892
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13920 25467 13923
rect 26252 13920 26280 13960
rect 26602 13948 26608 13960
rect 26660 13948 26666 14000
rect 26896 13929 26924 14016
rect 26881 13923 26939 13929
rect 26881 13920 26893 13923
rect 25455 13892 26280 13920
rect 26344 13892 26893 13920
rect 25455 13889 25467 13892
rect 25409 13883 25467 13889
rect 26344 13861 26372 13892
rect 26881 13889 26893 13892
rect 26927 13889 26939 13923
rect 26881 13883 26939 13889
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13920 27215 13923
rect 27264 13920 27292 14028
rect 27614 14016 27620 14028
rect 27672 14016 27678 14068
rect 28902 14016 28908 14068
rect 28960 14056 28966 14068
rect 29086 14056 29092 14068
rect 28960 14028 29092 14056
rect 28960 14016 28966 14028
rect 29086 14016 29092 14028
rect 29144 14056 29150 14068
rect 29144 14028 31432 14056
rect 29144 14016 29150 14028
rect 29564 13960 30788 13988
rect 27203 13892 27292 13920
rect 27203 13889 27215 13892
rect 27157 13883 27215 13889
rect 27522 13880 27528 13932
rect 27580 13920 27586 13932
rect 27580 13892 29408 13920
rect 27580 13880 27586 13892
rect 24397 13855 24455 13861
rect 24397 13821 24409 13855
rect 24443 13821 24455 13855
rect 24397 13815 24455 13821
rect 26237 13855 26295 13861
rect 26237 13821 26249 13855
rect 26283 13821 26295 13855
rect 26237 13815 26295 13821
rect 26329 13855 26387 13861
rect 26329 13821 26341 13855
rect 26375 13821 26387 13855
rect 26329 13815 26387 13821
rect 24026 13716 24032 13728
rect 22388 13688 24032 13716
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 24210 13676 24216 13728
rect 24268 13676 24274 13728
rect 26252 13716 26280 13815
rect 26418 13812 26424 13864
rect 26476 13812 26482 13864
rect 26602 13812 26608 13864
rect 26660 13812 26666 13864
rect 26694 13812 26700 13864
rect 26752 13812 26758 13864
rect 26786 13812 26792 13864
rect 26844 13812 26850 13864
rect 27062 13812 27068 13864
rect 27120 13812 27126 13864
rect 28994 13812 29000 13864
rect 29052 13812 29058 13864
rect 29086 13812 29092 13864
rect 29144 13812 29150 13864
rect 29380 13861 29408 13892
rect 29564 13861 29592 13960
rect 30006 13880 30012 13932
rect 30064 13920 30070 13932
rect 30064 13892 30696 13920
rect 30064 13880 30070 13892
rect 29365 13855 29423 13861
rect 29365 13821 29377 13855
rect 29411 13821 29423 13855
rect 29365 13815 29423 13821
rect 29549 13855 29607 13861
rect 29549 13821 29561 13855
rect 29595 13852 29607 13855
rect 29730 13852 29736 13864
rect 29595 13824 29736 13852
rect 29595 13821 29607 13824
rect 29549 13815 29607 13821
rect 29730 13812 29736 13824
rect 29788 13812 29794 13864
rect 29822 13812 29828 13864
rect 29880 13812 29886 13864
rect 29914 13812 29920 13864
rect 29972 13852 29978 13864
rect 30122 13852 30328 13862
rect 30668 13861 30696 13892
rect 30760 13861 30788 13960
rect 30377 13855 30435 13861
rect 30377 13852 30389 13855
rect 29972 13834 30389 13852
rect 29972 13824 30150 13834
rect 30300 13824 30389 13834
rect 29972 13812 29978 13824
rect 30377 13821 30389 13824
rect 30423 13821 30435 13855
rect 30377 13815 30435 13821
rect 30653 13855 30711 13861
rect 30653 13821 30665 13855
rect 30699 13821 30711 13855
rect 30653 13815 30711 13821
rect 30745 13855 30803 13861
rect 30745 13821 30757 13855
rect 30791 13821 30803 13855
rect 30745 13815 30803 13821
rect 31202 13812 31208 13864
rect 31260 13812 31266 13864
rect 31404 13861 31432 14028
rect 32122 14016 32128 14068
rect 32180 14056 32186 14068
rect 32309 14059 32367 14065
rect 32309 14056 32321 14059
rect 32180 14028 32321 14056
rect 32180 14016 32186 14028
rect 32309 14025 32321 14028
rect 32355 14025 32367 14059
rect 32309 14019 32367 14025
rect 32398 14016 32404 14068
rect 32456 14016 32462 14068
rect 32858 14016 32864 14068
rect 32916 14056 32922 14068
rect 33229 14059 33287 14065
rect 33229 14056 33241 14059
rect 32916 14028 33241 14056
rect 32916 14016 32922 14028
rect 33229 14025 33241 14028
rect 33275 14025 33287 14059
rect 33229 14019 33287 14025
rect 32416 13920 32444 14016
rect 32861 13923 32919 13929
rect 32861 13920 32873 13923
rect 32416 13892 32873 13920
rect 32861 13889 32873 13892
rect 32907 13889 32919 13923
rect 32861 13883 32919 13889
rect 33594 13880 33600 13932
rect 33652 13920 33658 13932
rect 33781 13923 33839 13929
rect 33781 13920 33793 13923
rect 33652 13892 33793 13920
rect 33652 13880 33658 13892
rect 33781 13889 33793 13892
rect 33827 13889 33839 13923
rect 33781 13883 33839 13889
rect 31389 13855 31447 13861
rect 31389 13821 31401 13855
rect 31435 13821 31447 13855
rect 31389 13815 31447 13821
rect 31478 13812 31484 13864
rect 31536 13812 31542 13864
rect 27430 13744 27436 13796
rect 27488 13744 27494 13796
rect 29012 13784 29040 13812
rect 28658 13756 29040 13784
rect 30190 13744 30196 13796
rect 30248 13744 30254 13796
rect 30558 13744 30564 13796
rect 30616 13744 30622 13796
rect 27706 13716 27712 13728
rect 26252 13688 27712 13716
rect 27706 13676 27712 13688
rect 27764 13676 27770 13728
rect 28902 13676 28908 13728
rect 28960 13676 28966 13728
rect 29086 13676 29092 13728
rect 29144 13716 29150 13728
rect 29181 13719 29239 13725
rect 29181 13716 29193 13719
rect 29144 13688 29193 13716
rect 29144 13676 29150 13688
rect 29181 13685 29193 13688
rect 29227 13716 29239 13719
rect 30466 13716 30472 13728
rect 29227 13688 30472 13716
rect 29227 13685 29239 13688
rect 29181 13679 29239 13685
rect 30466 13676 30472 13688
rect 30524 13676 30530 13728
rect 30929 13719 30987 13725
rect 30929 13685 30941 13719
rect 30975 13716 30987 13719
rect 31294 13716 31300 13728
rect 30975 13688 31300 13716
rect 30975 13685 30987 13688
rect 30929 13679 30987 13685
rect 31294 13676 31300 13688
rect 31352 13676 31358 13728
rect 2760 13626 34316 13648
rect 2760 13574 7210 13626
rect 7262 13574 7274 13626
rect 7326 13574 7338 13626
rect 7390 13574 7402 13626
rect 7454 13574 7466 13626
rect 7518 13574 15099 13626
rect 15151 13574 15163 13626
rect 15215 13574 15227 13626
rect 15279 13574 15291 13626
rect 15343 13574 15355 13626
rect 15407 13574 22988 13626
rect 23040 13574 23052 13626
rect 23104 13574 23116 13626
rect 23168 13574 23180 13626
rect 23232 13574 23244 13626
rect 23296 13574 30877 13626
rect 30929 13574 30941 13626
rect 30993 13574 31005 13626
rect 31057 13574 31069 13626
rect 31121 13574 31133 13626
rect 31185 13574 34316 13626
rect 2760 13552 34316 13574
rect 4617 13515 4675 13521
rect 4617 13481 4629 13515
rect 4663 13512 4675 13515
rect 5442 13512 5448 13524
rect 4663 13484 5448 13512
rect 4663 13481 4675 13484
rect 4617 13475 4675 13481
rect 5442 13472 5448 13484
rect 5500 13472 5506 13524
rect 6270 13472 6276 13524
rect 6328 13512 6334 13524
rect 6641 13515 6699 13521
rect 6641 13512 6653 13515
rect 6328 13484 6653 13512
rect 6328 13472 6334 13484
rect 6641 13481 6653 13484
rect 6687 13481 6699 13515
rect 6641 13475 6699 13481
rect 7837 13515 7895 13521
rect 7837 13481 7849 13515
rect 7883 13512 7895 13515
rect 7926 13512 7932 13524
rect 7883 13484 7932 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 9122 13472 9128 13524
rect 9180 13512 9186 13524
rect 9309 13515 9367 13521
rect 9309 13512 9321 13515
rect 9180 13484 9321 13512
rect 9180 13472 9186 13484
rect 9309 13481 9321 13484
rect 9355 13512 9367 13515
rect 9585 13515 9643 13521
rect 9585 13512 9597 13515
rect 9355 13484 9597 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 9585 13481 9597 13484
rect 9631 13512 9643 13515
rect 9858 13512 9864 13524
rect 9631 13484 9864 13512
rect 9631 13481 9643 13484
rect 9585 13475 9643 13481
rect 9858 13472 9864 13484
rect 9916 13472 9922 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 11241 13515 11299 13521
rect 10468 13484 11192 13512
rect 10468 13472 10474 13484
rect 5534 13404 5540 13456
rect 5592 13404 5598 13456
rect 6089 13447 6147 13453
rect 6089 13413 6101 13447
rect 6135 13444 6147 13447
rect 6454 13444 6460 13456
rect 6135 13416 6460 13444
rect 6135 13413 6147 13416
rect 6089 13407 6147 13413
rect 6454 13404 6460 13416
rect 6512 13404 6518 13456
rect 8478 13404 8484 13456
rect 8536 13444 8542 13456
rect 9953 13447 10011 13453
rect 9953 13444 9965 13447
rect 8536 13416 9965 13444
rect 8536 13404 8542 13416
rect 9953 13413 9965 13416
rect 9999 13413 10011 13447
rect 9953 13407 10011 13413
rect 10505 13447 10563 13453
rect 10505 13413 10517 13447
rect 10551 13444 10563 13447
rect 10594 13444 10600 13456
rect 10551 13416 10600 13444
rect 10551 13413 10563 13416
rect 10505 13407 10563 13413
rect 10594 13404 10600 13416
rect 10652 13404 10658 13456
rect 11164 13444 11192 13484
rect 11241 13481 11253 13515
rect 11287 13512 11299 13515
rect 11609 13515 11667 13521
rect 11609 13512 11621 13515
rect 11287 13484 11621 13512
rect 11287 13481 11299 13484
rect 11241 13475 11299 13481
rect 11609 13481 11621 13484
rect 11655 13512 11667 13515
rect 11698 13512 11704 13524
rect 11655 13484 11704 13512
rect 11655 13481 11667 13484
rect 11609 13475 11667 13481
rect 11698 13472 11704 13484
rect 11756 13472 11762 13524
rect 12894 13472 12900 13524
rect 12952 13512 12958 13524
rect 13449 13515 13507 13521
rect 13449 13512 13461 13515
rect 12952 13484 13461 13512
rect 12952 13472 12958 13484
rect 13449 13481 13461 13484
rect 13495 13481 13507 13515
rect 13449 13475 13507 13481
rect 14458 13472 14464 13524
rect 14516 13512 14522 13524
rect 15562 13512 15568 13524
rect 14516 13484 15568 13512
rect 14516 13472 14522 13484
rect 15562 13472 15568 13484
rect 15620 13472 15626 13524
rect 15746 13472 15752 13524
rect 15804 13472 15810 13524
rect 16853 13515 16911 13521
rect 16040 13484 16804 13512
rect 12986 13444 12992 13456
rect 11164 13416 12992 13444
rect 12986 13404 12992 13416
rect 13044 13404 13050 13456
rect 13078 13404 13084 13456
rect 13136 13444 13142 13456
rect 13658 13447 13716 13453
rect 13658 13444 13670 13447
rect 13136 13416 13670 13444
rect 13136 13404 13142 13416
rect 13658 13413 13670 13416
rect 13704 13444 13716 13447
rect 13814 13444 13820 13456
rect 13704 13416 13820 13444
rect 13704 13413 13716 13416
rect 13658 13407 13716 13413
rect 13814 13404 13820 13416
rect 13872 13404 13878 13456
rect 14550 13404 14556 13456
rect 14608 13444 14614 13456
rect 15764 13444 15792 13472
rect 14608 13416 15792 13444
rect 14608 13404 14614 13416
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4120 13348 4261 13376
rect 4120 13336 4126 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4249 13339 4307 13345
rect 6362 13336 6368 13388
rect 6420 13336 6426 13388
rect 6546 13336 6552 13388
rect 6604 13376 6610 13388
rect 6825 13379 6883 13385
rect 6825 13376 6837 13379
rect 6604 13348 6837 13376
rect 6604 13336 6610 13348
rect 6825 13345 6837 13348
rect 6871 13345 6883 13379
rect 6825 13339 6883 13345
rect 8202 13336 8208 13388
rect 8260 13336 8266 13388
rect 10137 13379 10195 13385
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 10410 13376 10416 13388
rect 10183 13348 10416 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 10410 13336 10416 13348
rect 10468 13376 10474 13388
rect 11606 13376 11612 13388
rect 10468 13348 11612 13376
rect 10468 13336 10474 13348
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 13170 13336 13176 13388
rect 13228 13336 13234 13388
rect 13541 13379 13599 13385
rect 13541 13376 13553 13379
rect 13372 13348 13553 13376
rect 1302 13268 1308 13320
rect 1360 13308 1366 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 1360 13280 3249 13308
rect 1360 13268 1366 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 6380 13308 6408 13336
rect 13372 13320 13400 13348
rect 13541 13345 13553 13348
rect 13587 13345 13599 13379
rect 14734 13376 14740 13388
rect 13541 13339 13599 13345
rect 13832 13348 14740 13376
rect 3237 13271 3295 13277
rect 6288 13280 6408 13308
rect 7469 13311 7527 13317
rect 6288 13184 6316 13280
rect 7469 13277 7481 13311
rect 7515 13308 7527 13311
rect 8018 13308 8024 13320
rect 7515 13280 8024 13308
rect 7515 13277 7527 13280
rect 7469 13271 7527 13277
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13308 8447 13311
rect 11793 13311 11851 13317
rect 8435 13280 8800 13308
rect 8435 13277 8447 13280
rect 8389 13271 8447 13277
rect 6270 13132 6276 13184
rect 6328 13132 6334 13184
rect 6362 13132 6368 13184
rect 6420 13172 6426 13184
rect 8021 13175 8079 13181
rect 8021 13172 8033 13175
rect 6420 13144 8033 13172
rect 6420 13132 6426 13144
rect 8021 13141 8033 13144
rect 8067 13172 8079 13175
rect 8110 13172 8116 13184
rect 8067 13144 8116 13172
rect 8067 13141 8079 13144
rect 8021 13135 8079 13141
rect 8110 13132 8116 13144
rect 8168 13132 8174 13184
rect 8772 13181 8800 13280
rect 11793 13277 11805 13311
rect 11839 13308 11851 13311
rect 12066 13308 12072 13320
rect 11839 13280 12072 13308
rect 11839 13277 11851 13280
rect 11793 13271 11851 13277
rect 12066 13268 12072 13280
rect 12124 13268 12130 13320
rect 13354 13268 13360 13320
rect 13412 13268 13418 13320
rect 13832 13249 13860 13348
rect 14734 13336 14740 13348
rect 14792 13336 14798 13388
rect 15013 13379 15071 13385
rect 15013 13345 15025 13379
rect 15059 13376 15071 13379
rect 15059 13348 15332 13376
rect 15059 13345 15071 13348
rect 15013 13339 15071 13345
rect 14182 13268 14188 13320
rect 14240 13268 14246 13320
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13308 14427 13311
rect 15304 13308 15332 13348
rect 15562 13336 15568 13388
rect 15620 13336 15626 13388
rect 16040 13385 16068 13484
rect 16390 13404 16396 13456
rect 16448 13404 16454 13456
rect 16776 13444 16804 13484
rect 16853 13481 16865 13515
rect 16899 13512 16911 13515
rect 17494 13512 17500 13524
rect 16899 13484 17500 13512
rect 16899 13481 16911 13484
rect 16853 13475 16911 13481
rect 17494 13472 17500 13484
rect 17552 13472 17558 13524
rect 17589 13515 17647 13521
rect 17589 13481 17601 13515
rect 17635 13512 17647 13515
rect 17678 13512 17684 13524
rect 17635 13484 17684 13512
rect 17635 13481 17647 13484
rect 17589 13475 17647 13481
rect 17678 13472 17684 13484
rect 17736 13472 17742 13524
rect 20625 13515 20683 13521
rect 20625 13481 20637 13515
rect 20671 13512 20683 13515
rect 20714 13512 20720 13524
rect 20671 13484 20720 13512
rect 20671 13481 20683 13484
rect 20625 13475 20683 13481
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 20806 13472 20812 13524
rect 20864 13472 20870 13524
rect 21174 13472 21180 13524
rect 21232 13512 21238 13524
rect 21637 13515 21695 13521
rect 21637 13512 21649 13515
rect 21232 13484 21649 13512
rect 21232 13472 21238 13484
rect 21637 13481 21649 13484
rect 21683 13481 21695 13515
rect 23474 13512 23480 13524
rect 21637 13475 21695 13481
rect 22066 13484 23480 13512
rect 18046 13444 18052 13456
rect 16776 13416 18052 13444
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 16025 13379 16083 13385
rect 16025 13345 16037 13379
rect 16071 13345 16083 13379
rect 16025 13339 16083 13345
rect 16301 13379 16359 13385
rect 16301 13345 16313 13379
rect 16347 13376 16359 13379
rect 16408 13376 16436 13404
rect 16347 13348 16436 13376
rect 16347 13345 16359 13348
rect 16301 13339 16359 13345
rect 16482 13336 16488 13388
rect 16540 13336 16546 13388
rect 16758 13336 16764 13388
rect 16816 13376 16822 13388
rect 16945 13379 17003 13385
rect 16945 13376 16957 13379
rect 16816 13348 16957 13376
rect 16816 13336 16822 13348
rect 16945 13345 16957 13348
rect 16991 13345 17003 13379
rect 16945 13339 17003 13345
rect 17221 13379 17279 13385
rect 17221 13345 17233 13379
rect 17267 13376 17279 13379
rect 17402 13376 17408 13388
rect 17267 13348 17408 13376
rect 17267 13345 17279 13348
rect 17221 13339 17279 13345
rect 17402 13336 17408 13348
rect 17460 13336 17466 13388
rect 17770 13336 17776 13388
rect 17828 13336 17834 13388
rect 17957 13379 18015 13385
rect 17957 13345 17969 13379
rect 18003 13345 18015 13379
rect 17957 13339 18015 13345
rect 16577 13311 16635 13317
rect 14415 13280 15056 13308
rect 15304 13280 15516 13308
rect 14415 13277 14427 13280
rect 14369 13271 14427 13277
rect 15028 13252 15056 13280
rect 13817 13243 13875 13249
rect 13817 13209 13829 13243
rect 13863 13209 13875 13243
rect 13817 13203 13875 13209
rect 14642 13200 14648 13252
rect 14700 13240 14706 13252
rect 14829 13243 14887 13249
rect 14829 13240 14841 13243
rect 14700 13212 14841 13240
rect 14700 13200 14706 13212
rect 14829 13209 14841 13212
rect 14875 13209 14887 13243
rect 14829 13203 14887 13209
rect 15010 13200 15016 13252
rect 15068 13200 15074 13252
rect 15488 13184 15516 13280
rect 16577 13277 16589 13311
rect 16623 13308 16635 13311
rect 16850 13308 16856 13320
rect 16623 13280 16856 13308
rect 16623 13277 16635 13280
rect 16577 13271 16635 13277
rect 16850 13268 16856 13280
rect 16908 13308 16914 13320
rect 16908 13280 17080 13308
rect 16908 13268 16914 13280
rect 8757 13175 8815 13181
rect 8757 13141 8769 13175
rect 8803 13172 8815 13175
rect 9030 13172 9036 13184
rect 8803 13144 9036 13172
rect 8803 13141 8815 13144
rect 8757 13135 8815 13141
rect 9030 13132 9036 13144
rect 9088 13132 9094 13184
rect 12345 13175 12403 13181
rect 12345 13141 12357 13175
rect 12391 13172 12403 13175
rect 12434 13172 12440 13184
rect 12391 13144 12440 13172
rect 12391 13141 12403 13144
rect 12345 13135 12403 13141
rect 12434 13132 12440 13144
rect 12492 13172 12498 13184
rect 12894 13172 12900 13184
rect 12492 13144 12900 13172
rect 12492 13132 12498 13144
rect 12894 13132 12900 13144
rect 12952 13132 12958 13184
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 15470 13172 15476 13184
rect 13044 13144 15476 13172
rect 13044 13132 13050 13144
rect 15470 13132 15476 13144
rect 15528 13132 15534 13184
rect 15930 13132 15936 13184
rect 15988 13132 15994 13184
rect 16574 13132 16580 13184
rect 16632 13132 16638 13184
rect 17052 13181 17080 13280
rect 17126 13268 17132 13320
rect 17184 13268 17190 13320
rect 17310 13268 17316 13320
rect 17368 13308 17374 13320
rect 17678 13308 17684 13320
rect 17368 13280 17684 13308
rect 17368 13268 17374 13280
rect 17678 13268 17684 13280
rect 17736 13308 17742 13320
rect 17972 13308 18000 13339
rect 18598 13336 18604 13388
rect 18656 13376 18662 13388
rect 18782 13376 18788 13388
rect 18656 13348 18788 13376
rect 18656 13336 18662 13348
rect 18782 13336 18788 13348
rect 18840 13376 18846 13388
rect 19061 13379 19119 13385
rect 19061 13376 19073 13379
rect 18840 13348 19073 13376
rect 18840 13336 18846 13348
rect 19061 13345 19073 13348
rect 19107 13345 19119 13379
rect 19061 13339 19119 13345
rect 19150 13336 19156 13388
rect 19208 13336 19214 13388
rect 20441 13379 20499 13385
rect 20441 13376 20453 13379
rect 19352 13348 20453 13376
rect 17736 13280 18000 13308
rect 17736 13268 17742 13280
rect 17862 13200 17868 13252
rect 17920 13240 17926 13252
rect 19352 13240 19380 13348
rect 20441 13345 20453 13348
rect 20487 13376 20499 13379
rect 20622 13376 20628 13388
rect 20487 13348 20628 13376
rect 20487 13345 20499 13348
rect 20441 13339 20499 13345
rect 20622 13336 20628 13348
rect 20680 13336 20686 13388
rect 20717 13379 20775 13385
rect 20717 13345 20729 13379
rect 20763 13376 20775 13379
rect 20824 13376 20852 13472
rect 20763 13348 20852 13376
rect 20763 13345 20775 13348
rect 20717 13339 20775 13345
rect 20898 13336 20904 13388
rect 20956 13376 20962 13388
rect 21729 13379 21787 13385
rect 21729 13376 21741 13379
rect 20956 13348 21741 13376
rect 20956 13336 20962 13348
rect 21729 13345 21741 13348
rect 21775 13345 21787 13379
rect 21729 13339 21787 13345
rect 22066 13320 22094 13484
rect 23474 13472 23480 13484
rect 23532 13472 23538 13524
rect 23845 13515 23903 13521
rect 23845 13481 23857 13515
rect 23891 13512 23903 13515
rect 24210 13512 24216 13524
rect 23891 13484 24216 13512
rect 23891 13481 23903 13484
rect 23845 13475 23903 13481
rect 24210 13472 24216 13484
rect 24268 13472 24274 13524
rect 25682 13472 25688 13524
rect 25740 13512 25746 13524
rect 25869 13515 25927 13521
rect 25869 13512 25881 13515
rect 25740 13484 25881 13512
rect 25740 13472 25746 13484
rect 25869 13481 25881 13484
rect 25915 13481 25927 13515
rect 25869 13475 25927 13481
rect 26510 13472 26516 13524
rect 26568 13472 26574 13524
rect 27430 13472 27436 13524
rect 27488 13472 27494 13524
rect 28810 13512 28816 13524
rect 28644 13484 28816 13512
rect 26142 13404 26148 13456
rect 26200 13404 26206 13456
rect 26528 13444 26556 13472
rect 26855 13447 26913 13453
rect 26855 13444 26867 13447
rect 26528 13416 26867 13444
rect 26855 13413 26867 13416
rect 26901 13413 26913 13447
rect 26855 13407 26913 13413
rect 26973 13447 27031 13453
rect 26973 13413 26985 13447
rect 27019 13444 27031 13447
rect 28261 13447 28319 13453
rect 28261 13444 28273 13447
rect 27019 13416 28273 13444
rect 27019 13413 27031 13416
rect 26973 13407 27031 13413
rect 28261 13413 28273 13416
rect 28307 13413 28319 13447
rect 28261 13407 28319 13413
rect 22189 13379 22247 13385
rect 22189 13345 22201 13379
rect 22235 13376 22247 13379
rect 22646 13376 22652 13388
rect 22235 13348 22652 13376
rect 22235 13345 22247 13348
rect 22189 13339 22247 13345
rect 20257 13311 20315 13317
rect 20257 13277 20269 13311
rect 20303 13308 20315 13311
rect 20993 13311 21051 13317
rect 20993 13308 21005 13311
rect 20303 13280 21005 13308
rect 20303 13277 20315 13280
rect 20257 13271 20315 13277
rect 20993 13277 21005 13280
rect 21039 13277 21051 13311
rect 20993 13271 21051 13277
rect 22002 13268 22008 13320
rect 22060 13280 22094 13320
rect 22060 13268 22066 13280
rect 17920 13212 19380 13240
rect 17920 13200 17926 13212
rect 17037 13175 17095 13181
rect 17037 13141 17049 13175
rect 17083 13141 17095 13175
rect 17037 13135 17095 13141
rect 17310 13132 17316 13184
rect 17368 13172 17374 13184
rect 17972 13181 18000 13212
rect 19610 13200 19616 13252
rect 19668 13240 19674 13252
rect 20165 13243 20223 13249
rect 20165 13240 20177 13243
rect 19668 13212 20177 13240
rect 19668 13200 19674 13212
rect 20165 13209 20177 13212
rect 20211 13240 20223 13243
rect 22204 13240 22232 13339
rect 22646 13336 22652 13348
rect 22704 13336 22710 13388
rect 23937 13379 23995 13385
rect 23937 13345 23949 13379
rect 23983 13376 23995 13379
rect 24581 13379 24639 13385
rect 24581 13376 24593 13379
rect 23983 13348 24593 13376
rect 23983 13345 23995 13348
rect 23937 13339 23995 13345
rect 24581 13345 24593 13348
rect 24627 13345 24639 13379
rect 24581 13339 24639 13345
rect 22741 13311 22799 13317
rect 22741 13277 22753 13311
rect 22787 13277 22799 13311
rect 22741 13271 22799 13277
rect 20211 13212 22232 13240
rect 22756 13240 22784 13271
rect 23842 13268 23848 13320
rect 23900 13308 23906 13320
rect 24026 13308 24032 13320
rect 23900 13280 24032 13308
rect 23900 13268 23906 13280
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 24486 13268 24492 13320
rect 24544 13268 24550 13320
rect 24596 13308 24624 13339
rect 24670 13336 24676 13388
rect 24728 13336 24734 13388
rect 26050 13336 26056 13388
rect 26108 13336 26114 13388
rect 26234 13336 26240 13388
rect 26292 13336 26298 13388
rect 26326 13336 26332 13388
rect 26384 13385 26390 13388
rect 26384 13379 26413 13385
rect 26401 13345 26413 13379
rect 26384 13339 26413 13345
rect 26384 13336 26390 13339
rect 27062 13336 27068 13388
rect 27120 13336 27126 13388
rect 27157 13379 27215 13385
rect 27157 13345 27169 13379
rect 27203 13376 27215 13379
rect 27890 13376 27896 13388
rect 27203 13348 27896 13376
rect 27203 13345 27215 13348
rect 27157 13339 27215 13345
rect 27890 13336 27896 13348
rect 27948 13336 27954 13388
rect 28169 13379 28227 13385
rect 28169 13345 28181 13379
rect 28215 13376 28227 13379
rect 28215 13348 28304 13376
rect 28215 13345 28227 13348
rect 28169 13339 28227 13345
rect 25133 13311 25191 13317
rect 25133 13308 25145 13311
rect 24596 13280 25145 13308
rect 25133 13277 25145 13280
rect 25179 13277 25191 13311
rect 25133 13271 25191 13277
rect 25682 13268 25688 13320
rect 25740 13268 25746 13320
rect 26513 13311 26571 13317
rect 26513 13277 26525 13311
rect 26559 13277 26571 13311
rect 26513 13271 26571 13277
rect 23477 13243 23535 13249
rect 23477 13240 23489 13243
rect 22756 13212 23489 13240
rect 20211 13209 20223 13212
rect 20165 13203 20223 13209
rect 23477 13209 23489 13212
rect 23523 13209 23535 13243
rect 26528 13240 26556 13271
rect 26602 13268 26608 13320
rect 26660 13308 26666 13320
rect 26697 13311 26755 13317
rect 26697 13308 26709 13311
rect 26660 13280 26709 13308
rect 26660 13268 26666 13280
rect 26697 13277 26709 13280
rect 26743 13308 26755 13311
rect 27341 13311 27399 13317
rect 26743 13280 27292 13308
rect 26743 13277 26755 13280
rect 26697 13271 26755 13277
rect 26970 13240 26976 13252
rect 23477 13203 23535 13209
rect 24136 13212 26464 13240
rect 26528 13212 26976 13240
rect 24136 13184 24164 13212
rect 17405 13175 17463 13181
rect 17405 13172 17417 13175
rect 17368 13144 17417 13172
rect 17368 13132 17374 13144
rect 17405 13141 17417 13144
rect 17451 13141 17463 13175
rect 17405 13135 17463 13141
rect 17957 13175 18015 13181
rect 17957 13141 17969 13175
rect 18003 13141 18015 13175
rect 17957 13135 18015 13141
rect 19242 13132 19248 13184
rect 19300 13132 19306 13184
rect 19334 13132 19340 13184
rect 19392 13172 19398 13184
rect 21726 13172 21732 13184
rect 19392 13144 21732 13172
rect 19392 13132 19398 13144
rect 21726 13132 21732 13144
rect 21784 13132 21790 13184
rect 22094 13132 22100 13184
rect 22152 13172 22158 13184
rect 22189 13175 22247 13181
rect 22189 13172 22201 13175
rect 22152 13144 22201 13172
rect 22152 13132 22158 13144
rect 22189 13141 22201 13144
rect 22235 13172 22247 13175
rect 22278 13172 22284 13184
rect 22235 13144 22284 13172
rect 22235 13141 22247 13144
rect 22189 13135 22247 13141
rect 22278 13132 22284 13144
rect 22336 13132 22342 13184
rect 22370 13132 22376 13184
rect 22428 13132 22434 13184
rect 23290 13132 23296 13184
rect 23348 13132 23354 13184
rect 24118 13132 24124 13184
rect 24176 13132 24182 13184
rect 25038 13132 25044 13184
rect 25096 13132 25102 13184
rect 26436 13172 26464 13212
rect 26970 13200 26976 13212
rect 27028 13200 27034 13252
rect 27264 13240 27292 13280
rect 27341 13277 27353 13311
rect 27387 13308 27399 13311
rect 27985 13311 28043 13317
rect 27985 13308 27997 13311
rect 27387 13280 27997 13308
rect 27387 13277 27399 13280
rect 27341 13271 27399 13277
rect 27985 13277 27997 13280
rect 28031 13277 28043 13311
rect 27985 13271 28043 13277
rect 28276 13240 28304 13348
rect 28350 13336 28356 13388
rect 28408 13336 28414 13388
rect 28644 13385 28672 13484
rect 28810 13472 28816 13484
rect 28868 13472 28874 13524
rect 29178 13472 29184 13524
rect 29236 13512 29242 13524
rect 29454 13512 29460 13524
rect 29236 13484 29460 13512
rect 29236 13472 29242 13484
rect 29454 13472 29460 13484
rect 29512 13472 29518 13524
rect 30282 13512 30288 13524
rect 29748 13484 30288 13512
rect 28721 13447 28779 13453
rect 28721 13413 28733 13447
rect 28767 13444 28779 13447
rect 29748 13444 29776 13484
rect 30282 13472 30288 13484
rect 30340 13472 30346 13524
rect 30374 13472 30380 13524
rect 30432 13512 30438 13524
rect 30837 13515 30895 13521
rect 30837 13512 30849 13515
rect 30432 13484 30849 13512
rect 30432 13472 30438 13484
rect 30837 13481 30849 13484
rect 30883 13481 30895 13515
rect 31478 13512 31484 13524
rect 30837 13475 30895 13481
rect 30944 13484 31484 13512
rect 28767 13416 29776 13444
rect 30024 13416 30420 13444
rect 28767 13413 28779 13416
rect 28721 13407 28779 13413
rect 30024 13388 30052 13416
rect 28629 13379 28687 13385
rect 28629 13345 28641 13379
rect 28675 13345 28687 13379
rect 28629 13339 28687 13345
rect 28813 13379 28871 13385
rect 28813 13345 28825 13379
rect 28859 13345 28871 13379
rect 28813 13339 28871 13345
rect 28828 13308 28856 13339
rect 28902 13336 28908 13388
rect 28960 13382 28966 13388
rect 28997 13382 29055 13385
rect 28960 13379 29055 13382
rect 28960 13354 29009 13379
rect 28960 13336 28966 13354
rect 28997 13345 29009 13354
rect 29043 13345 29055 13379
rect 28997 13339 29055 13345
rect 29086 13336 29092 13388
rect 29144 13336 29150 13388
rect 30006 13336 30012 13388
rect 30064 13336 30070 13388
rect 30190 13336 30196 13388
rect 30248 13336 30254 13388
rect 30392 13385 30420 13416
rect 30466 13404 30472 13456
rect 30524 13444 30530 13456
rect 30944 13444 30972 13484
rect 31478 13472 31484 13484
rect 31536 13472 31542 13524
rect 32048 13484 32812 13512
rect 32048 13444 32076 13484
rect 30524 13416 30972 13444
rect 31878 13416 32076 13444
rect 30524 13404 30530 13416
rect 32306 13404 32312 13456
rect 32364 13444 32370 13456
rect 32784 13453 32812 13484
rect 33042 13472 33048 13524
rect 33100 13472 33106 13524
rect 35158 13472 35164 13524
rect 35216 13472 35222 13524
rect 32769 13447 32827 13453
rect 32364 13416 32628 13444
rect 32364 13404 32370 13416
rect 32600 13388 32628 13416
rect 32769 13413 32781 13447
rect 32815 13413 32827 13447
rect 32769 13407 32827 13413
rect 30377 13379 30435 13385
rect 30377 13345 30389 13379
rect 30423 13345 30435 13379
rect 30377 13339 30435 13345
rect 30561 13379 30619 13385
rect 30561 13345 30573 13379
rect 30607 13345 30619 13379
rect 30561 13339 30619 13345
rect 29104 13308 29132 13336
rect 28828 13280 29132 13308
rect 29181 13311 29239 13317
rect 29181 13277 29193 13311
rect 29227 13308 29239 13311
rect 29227 13280 29316 13308
rect 29227 13277 29239 13280
rect 29181 13271 29239 13277
rect 29288 13252 29316 13280
rect 29914 13268 29920 13320
rect 29972 13308 29978 13320
rect 30576 13308 30604 13339
rect 32582 13336 32588 13388
rect 32640 13336 32646 13388
rect 32861 13379 32919 13385
rect 32861 13345 32873 13379
rect 32907 13376 32919 13379
rect 33060 13376 33088 13472
rect 32907 13348 33088 13376
rect 33965 13379 34023 13385
rect 32907 13345 32919 13348
rect 32861 13339 32919 13345
rect 33965 13345 33977 13379
rect 34011 13376 34023 13379
rect 35176 13376 35204 13472
rect 34011 13348 35204 13376
rect 34011 13345 34023 13348
rect 33965 13339 34023 13345
rect 29972 13280 30604 13308
rect 29972 13268 29978 13280
rect 32306 13268 32312 13320
rect 32364 13268 32370 13320
rect 29270 13240 29276 13252
rect 27264 13212 29276 13240
rect 29270 13200 29276 13212
rect 29328 13200 29334 13252
rect 29840 13212 30236 13240
rect 29840 13172 29868 13212
rect 26436 13144 29868 13172
rect 29914 13132 29920 13184
rect 29972 13172 29978 13184
rect 30101 13175 30159 13181
rect 30101 13172 30113 13175
rect 29972 13144 30113 13172
rect 29972 13132 29978 13144
rect 30101 13141 30113 13144
rect 30147 13141 30159 13175
rect 30208 13172 30236 13212
rect 32692 13212 33824 13240
rect 32692 13172 32720 13212
rect 33796 13181 33824 13212
rect 30208 13144 32720 13172
rect 33781 13175 33839 13181
rect 30101 13135 30159 13141
rect 33781 13141 33793 13175
rect 33827 13141 33839 13175
rect 33781 13135 33839 13141
rect 2760 13082 34316 13104
rect 2760 13030 6550 13082
rect 6602 13030 6614 13082
rect 6666 13030 6678 13082
rect 6730 13030 6742 13082
rect 6794 13030 6806 13082
rect 6858 13030 14439 13082
rect 14491 13030 14503 13082
rect 14555 13030 14567 13082
rect 14619 13030 14631 13082
rect 14683 13030 14695 13082
rect 14747 13030 22328 13082
rect 22380 13030 22392 13082
rect 22444 13030 22456 13082
rect 22508 13030 22520 13082
rect 22572 13030 22584 13082
rect 22636 13030 30217 13082
rect 30269 13030 30281 13082
rect 30333 13030 30345 13082
rect 30397 13030 30409 13082
rect 30461 13030 30473 13082
rect 30525 13030 34316 13082
rect 2760 13008 34316 13030
rect 3421 12971 3479 12977
rect 3421 12937 3433 12971
rect 3467 12968 3479 12971
rect 3789 12971 3847 12977
rect 3789 12968 3801 12971
rect 3467 12940 3801 12968
rect 3467 12937 3479 12940
rect 3421 12931 3479 12937
rect 3789 12937 3801 12940
rect 3835 12968 3847 12971
rect 3970 12968 3976 12980
rect 3835 12940 3976 12968
rect 3835 12937 3847 12940
rect 3789 12931 3847 12937
rect 3970 12928 3976 12940
rect 4028 12968 4034 12980
rect 4338 12968 4344 12980
rect 4028 12940 4344 12968
rect 4028 12928 4034 12940
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 6454 12928 6460 12980
rect 6512 12928 6518 12980
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 8938 12968 8944 12980
rect 8628 12940 8944 12968
rect 8628 12928 8634 12940
rect 8938 12928 8944 12940
rect 8996 12968 9002 12980
rect 9953 12971 10011 12977
rect 9953 12968 9965 12971
rect 8996 12940 9965 12968
rect 8996 12928 9002 12940
rect 9953 12937 9965 12940
rect 9999 12937 10011 12971
rect 12434 12968 12440 12980
rect 9953 12931 10011 12937
rect 11348 12940 12440 12968
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 6472 12832 6500 12928
rect 7576 12872 9076 12900
rect 7576 12841 7604 12872
rect 7561 12835 7619 12841
rect 4396 12804 5856 12832
rect 6472 12804 7420 12832
rect 4396 12792 4402 12804
rect 3878 12724 3884 12776
rect 3936 12724 3942 12776
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 5718 12724 5724 12776
rect 5776 12724 5782 12776
rect 5828 12764 5856 12804
rect 5902 12764 5908 12776
rect 5828 12736 5908 12764
rect 5902 12724 5908 12736
rect 5960 12764 5966 12776
rect 7392 12773 7420 12804
rect 7561 12801 7573 12835
rect 7607 12801 7619 12835
rect 7561 12795 7619 12801
rect 8128 12804 8984 12832
rect 8128 12776 8156 12804
rect 7101 12767 7159 12773
rect 5960 12736 6592 12764
rect 5960 12724 5966 12736
rect 5534 12656 5540 12708
rect 5592 12696 5598 12708
rect 5592 12668 6500 12696
rect 5592 12656 5598 12668
rect 6472 12640 6500 12668
rect 4522 12588 4528 12640
rect 4580 12588 4586 12640
rect 5261 12631 5319 12637
rect 5261 12597 5273 12631
rect 5307 12628 5319 12631
rect 5442 12628 5448 12640
rect 5307 12600 5448 12628
rect 5307 12597 5319 12600
rect 5261 12591 5319 12597
rect 5442 12588 5448 12600
rect 5500 12588 5506 12640
rect 6178 12588 6184 12640
rect 6236 12628 6242 12640
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 6236 12600 6377 12628
rect 6236 12588 6242 12600
rect 6365 12597 6377 12600
rect 6411 12597 6423 12631
rect 6365 12591 6423 12597
rect 6454 12588 6460 12640
rect 6512 12588 6518 12640
rect 6564 12628 6592 12736
rect 7101 12733 7113 12767
rect 7147 12733 7159 12767
rect 7101 12727 7159 12733
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 7116 12696 7144 12727
rect 7834 12724 7840 12776
rect 7892 12724 7898 12776
rect 8110 12724 8116 12776
rect 8168 12724 8174 12776
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 8956 12773 8984 12804
rect 8757 12767 8815 12773
rect 8757 12764 8769 12767
rect 8628 12736 8769 12764
rect 8628 12724 8634 12736
rect 8757 12733 8769 12736
rect 8803 12733 8815 12767
rect 8757 12727 8815 12733
rect 8941 12767 8999 12773
rect 8941 12733 8953 12767
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9048 12708 9076 12872
rect 11348 12841 11376 12940
rect 12434 12928 12440 12940
rect 12492 12928 12498 12980
rect 12710 12928 12716 12980
rect 12768 12968 12774 12980
rect 12986 12968 12992 12980
rect 12768 12940 12992 12968
rect 12768 12928 12774 12940
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13814 12928 13820 12980
rect 13872 12928 13878 12980
rect 16209 12971 16267 12977
rect 16209 12937 16221 12971
rect 16255 12968 16267 12971
rect 16298 12968 16304 12980
rect 16255 12940 16304 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16298 12928 16304 12940
rect 16356 12928 16362 12980
rect 16758 12928 16764 12980
rect 16816 12928 16822 12980
rect 16850 12928 16856 12980
rect 16908 12928 16914 12980
rect 17310 12928 17316 12980
rect 17368 12968 17374 12980
rect 17865 12971 17923 12977
rect 17865 12968 17877 12971
rect 17368 12940 17877 12968
rect 17368 12928 17374 12940
rect 17865 12937 17877 12940
rect 17911 12937 17923 12971
rect 17865 12931 17923 12937
rect 18046 12928 18052 12980
rect 18104 12928 18110 12980
rect 18138 12928 18144 12980
rect 18196 12968 18202 12980
rect 18598 12968 18604 12980
rect 18196 12940 18604 12968
rect 18196 12928 18202 12940
rect 18598 12928 18604 12940
rect 18656 12928 18662 12980
rect 19242 12928 19248 12980
rect 19300 12928 19306 12980
rect 20070 12928 20076 12980
rect 20128 12928 20134 12980
rect 20162 12928 20168 12980
rect 20220 12968 20226 12980
rect 20625 12971 20683 12977
rect 20625 12968 20637 12971
rect 20220 12940 20637 12968
rect 20220 12928 20226 12940
rect 20625 12937 20637 12940
rect 20671 12968 20683 12971
rect 22002 12968 22008 12980
rect 20671 12940 22008 12968
rect 20671 12937 20683 12940
rect 20625 12931 20683 12937
rect 22002 12928 22008 12940
rect 22060 12928 22066 12980
rect 22094 12928 22100 12980
rect 22152 12928 22158 12980
rect 22186 12928 22192 12980
rect 22244 12968 22250 12980
rect 22830 12968 22836 12980
rect 22244 12940 22836 12968
rect 22244 12928 22250 12940
rect 22830 12928 22836 12940
rect 22888 12928 22894 12980
rect 23290 12928 23296 12980
rect 23348 12928 23354 12980
rect 25133 12971 25191 12977
rect 25133 12937 25145 12971
rect 25179 12968 25191 12971
rect 25682 12968 25688 12980
rect 25179 12940 25688 12968
rect 25179 12937 25191 12940
rect 25133 12931 25191 12937
rect 25682 12928 25688 12940
rect 25740 12928 25746 12980
rect 26053 12971 26111 12977
rect 26053 12968 26065 12971
rect 25792 12940 26065 12968
rect 15010 12860 15016 12912
rect 15068 12900 15074 12912
rect 16022 12900 16028 12912
rect 15068 12872 16028 12900
rect 15068 12860 15074 12872
rect 16022 12860 16028 12872
rect 16080 12900 16086 12912
rect 17678 12900 17684 12912
rect 16080 12872 17080 12900
rect 16080 12860 16086 12872
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12801 11391 12835
rect 11333 12795 11391 12801
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12832 11575 12835
rect 11698 12832 11704 12844
rect 11563 12804 11704 12832
rect 11563 12801 11575 12804
rect 11517 12795 11575 12801
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12342 12832 12348 12844
rect 11808 12804 12348 12832
rect 9122 12724 9128 12776
rect 9180 12724 9186 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 9646 12736 10333 12764
rect 8294 12696 8300 12708
rect 7116 12668 8300 12696
rect 8294 12656 8300 12668
rect 8352 12656 8358 12708
rect 8849 12699 8907 12705
rect 8849 12665 8861 12699
rect 8895 12665 8907 12699
rect 8849 12659 8907 12665
rect 7193 12631 7251 12637
rect 7193 12628 7205 12631
rect 6564 12600 7205 12628
rect 7193 12597 7205 12600
rect 7239 12597 7251 12631
rect 7193 12591 7251 12597
rect 8478 12588 8484 12640
rect 8536 12588 8542 12640
rect 8570 12588 8576 12640
rect 8628 12588 8634 12640
rect 8864 12628 8892 12659
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 9646 12696 9674 12736
rect 10321 12733 10333 12736
rect 10367 12764 10379 12767
rect 11808 12764 11836 12804
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 13725 12835 13783 12841
rect 13725 12801 13737 12835
rect 13771 12832 13783 12835
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 13771 12804 14381 12832
rect 13771 12801 13783 12804
rect 13725 12795 13783 12801
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 15194 12792 15200 12844
rect 15252 12792 15258 12844
rect 15470 12792 15476 12844
rect 15528 12792 15534 12844
rect 16117 12835 16175 12841
rect 16117 12832 16129 12835
rect 15580 12804 16129 12832
rect 15580 12776 15608 12804
rect 16117 12801 16129 12804
rect 16163 12832 16175 12835
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 16163 12804 16405 12832
rect 16163 12801 16175 12804
rect 16117 12795 16175 12801
rect 16393 12801 16405 12804
rect 16439 12801 16451 12835
rect 16393 12795 16451 12801
rect 16592 12804 16988 12832
rect 16592 12776 16620 12804
rect 16960 12776 16988 12804
rect 10367 12736 11836 12764
rect 11885 12767 11943 12773
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 11885 12733 11897 12767
rect 11931 12733 11943 12767
rect 11885 12727 11943 12733
rect 9088 12668 9674 12696
rect 11900 12696 11928 12727
rect 11974 12724 11980 12776
rect 12032 12724 12038 12776
rect 15562 12724 15568 12776
rect 15620 12724 15626 12776
rect 16022 12724 16028 12776
rect 16080 12724 16086 12776
rect 16298 12724 16304 12776
rect 16356 12764 16362 12776
rect 16485 12767 16543 12773
rect 16485 12764 16497 12767
rect 16356 12736 16497 12764
rect 16356 12724 16362 12736
rect 16485 12733 16497 12736
rect 16531 12733 16543 12767
rect 16485 12727 16543 12733
rect 16574 12724 16580 12776
rect 16632 12724 16638 12776
rect 16758 12724 16764 12776
rect 16816 12724 16822 12776
rect 16942 12724 16948 12776
rect 17000 12724 17006 12776
rect 17052 12773 17080 12872
rect 17393 12872 17684 12900
rect 17393 12773 17421 12872
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 18064 12900 18092 12928
rect 18064 12872 19104 12900
rect 18785 12835 18843 12841
rect 18785 12832 18797 12835
rect 17512 12804 18797 12832
rect 17512 12773 17540 12804
rect 18785 12801 18797 12804
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12733 17095 12767
rect 17393 12767 17463 12773
rect 17393 12736 17417 12767
rect 17037 12727 17095 12733
rect 17405 12733 17417 12736
rect 17451 12733 17463 12767
rect 17405 12727 17463 12733
rect 17497 12767 17555 12773
rect 17497 12733 17509 12767
rect 17543 12733 17555 12767
rect 17497 12727 17555 12733
rect 17586 12724 17592 12776
rect 17644 12724 17650 12776
rect 18966 12724 18972 12776
rect 19024 12724 19030 12776
rect 19076 12773 19104 12872
rect 19260 12832 19288 12928
rect 20088 12841 20116 12928
rect 21453 12903 21511 12909
rect 21453 12869 21465 12903
rect 21499 12900 21511 12903
rect 21634 12900 21640 12912
rect 21499 12872 21640 12900
rect 21499 12869 21511 12872
rect 21453 12863 21511 12869
rect 21634 12860 21640 12872
rect 21692 12900 21698 12912
rect 22112 12900 22140 12928
rect 21692 12872 22140 12900
rect 21692 12860 21698 12872
rect 20073 12835 20131 12841
rect 19260 12804 19748 12832
rect 19061 12767 19119 12773
rect 19061 12733 19073 12767
rect 19107 12733 19119 12767
rect 19061 12727 19119 12733
rect 19337 12767 19395 12773
rect 19337 12733 19349 12767
rect 19383 12764 19395 12767
rect 19518 12764 19524 12776
rect 19383 12736 19524 12764
rect 19383 12733 19395 12736
rect 19337 12727 19395 12733
rect 19518 12724 19524 12736
rect 19576 12724 19582 12776
rect 19720 12773 19748 12804
rect 20073 12801 20085 12835
rect 20119 12801 20131 12835
rect 22848 12832 22876 12928
rect 23308 12900 23336 12928
rect 23308 12872 23520 12900
rect 23385 12835 23443 12841
rect 23385 12832 23397 12835
rect 22848 12804 23397 12832
rect 20073 12795 20131 12801
rect 23385 12801 23397 12804
rect 23431 12801 23443 12835
rect 23492 12832 23520 12872
rect 24670 12860 24676 12912
rect 24728 12900 24734 12912
rect 25792 12900 25820 12940
rect 26053 12937 26065 12940
rect 26099 12937 26111 12971
rect 26053 12931 26111 12937
rect 27706 12928 27712 12980
rect 27764 12928 27770 12980
rect 28810 12928 28816 12980
rect 28868 12968 28874 12980
rect 28997 12971 29055 12977
rect 28997 12968 29009 12971
rect 28868 12940 29009 12968
rect 28868 12928 28874 12940
rect 28997 12937 29009 12940
rect 29043 12937 29055 12971
rect 28997 12931 29055 12937
rect 31849 12971 31907 12977
rect 31849 12937 31861 12971
rect 31895 12968 31907 12971
rect 32306 12968 32312 12980
rect 31895 12940 32312 12968
rect 31895 12937 31907 12940
rect 31849 12931 31907 12937
rect 32306 12928 32312 12940
rect 32364 12928 32370 12980
rect 33781 12903 33839 12909
rect 33781 12900 33793 12903
rect 24728 12872 25820 12900
rect 25884 12872 33793 12900
rect 24728 12860 24734 12872
rect 23661 12835 23719 12841
rect 23661 12832 23673 12835
rect 23492 12804 23673 12832
rect 23385 12795 23443 12801
rect 23661 12801 23673 12804
rect 23707 12801 23719 12835
rect 23661 12795 23719 12801
rect 23750 12792 23756 12844
rect 23808 12832 23814 12844
rect 23808 12804 24900 12832
rect 23808 12792 23814 12804
rect 19613 12767 19671 12773
rect 19613 12733 19625 12767
rect 19659 12733 19671 12767
rect 19613 12727 19671 12733
rect 19705 12767 19763 12773
rect 19705 12733 19717 12767
rect 19751 12733 19763 12767
rect 19705 12727 19763 12733
rect 12158 12696 12164 12708
rect 11900 12668 12164 12696
rect 9088 12656 9094 12668
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 12253 12699 12311 12705
rect 12253 12665 12265 12699
rect 12299 12696 12311 12699
rect 12299 12668 12434 12696
rect 12299 12665 12311 12668
rect 12253 12659 12311 12665
rect 9585 12631 9643 12637
rect 9585 12628 9597 12631
rect 8864 12600 9597 12628
rect 9585 12597 9597 12600
rect 9631 12628 9643 12631
rect 10594 12628 10600 12640
rect 9631 12600 10600 12628
rect 9631 12597 9643 12600
rect 9585 12591 9643 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 10870 12588 10876 12640
rect 10928 12588 10934 12640
rect 11241 12631 11299 12637
rect 11241 12597 11253 12631
rect 11287 12628 11299 12631
rect 11422 12628 11428 12640
rect 11287 12600 11428 12628
rect 11287 12597 11299 12600
rect 11241 12591 11299 12597
rect 11422 12588 11428 12600
rect 11480 12588 11486 12640
rect 11606 12588 11612 12640
rect 11664 12628 11670 12640
rect 11793 12631 11851 12637
rect 11793 12628 11805 12631
rect 11664 12600 11805 12628
rect 11664 12588 11670 12600
rect 11793 12597 11805 12600
rect 11839 12597 11851 12631
rect 12406 12628 12434 12668
rect 12894 12656 12900 12708
rect 12952 12656 12958 12708
rect 14182 12656 14188 12708
rect 14240 12696 14246 12708
rect 15749 12699 15807 12705
rect 15749 12696 15761 12699
rect 14240 12668 15761 12696
rect 14240 12656 14246 12668
rect 15749 12665 15761 12668
rect 15795 12696 15807 12699
rect 15930 12696 15936 12708
rect 15795 12668 15936 12696
rect 15795 12665 15807 12668
rect 15749 12659 15807 12665
rect 15930 12656 15936 12668
rect 15988 12696 15994 12708
rect 17129 12699 17187 12705
rect 17129 12696 17141 12699
rect 15988 12668 17141 12696
rect 15988 12656 15994 12668
rect 17129 12665 17141 12668
rect 17175 12665 17187 12699
rect 17129 12659 17187 12665
rect 17221 12699 17279 12705
rect 17221 12665 17233 12699
rect 17267 12696 17279 12699
rect 17267 12668 17448 12696
rect 17267 12665 17279 12668
rect 17221 12659 17279 12665
rect 17420 12640 17448 12668
rect 17770 12656 17776 12708
rect 17828 12696 17834 12708
rect 18233 12699 18291 12705
rect 18233 12696 18245 12699
rect 17828 12668 18245 12696
rect 17828 12656 17834 12668
rect 18233 12665 18245 12668
rect 18279 12696 18291 12699
rect 18279 12668 19472 12696
rect 18279 12665 18291 12668
rect 18233 12659 18291 12665
rect 13170 12628 13176 12640
rect 12406 12600 13176 12628
rect 11793 12591 11851 12597
rect 13170 12588 13176 12600
rect 13228 12588 13234 12640
rect 14918 12588 14924 12640
rect 14976 12628 14982 12640
rect 15841 12631 15899 12637
rect 15841 12628 15853 12631
rect 14976 12600 15853 12628
rect 14976 12588 14982 12600
rect 15841 12597 15853 12600
rect 15887 12628 15899 12631
rect 17034 12628 17040 12640
rect 15887 12600 17040 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 17034 12588 17040 12600
rect 17092 12628 17098 12640
rect 17402 12628 17408 12640
rect 17092 12600 17408 12628
rect 17092 12588 17098 12600
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 17856 12631 17914 12637
rect 17856 12597 17868 12631
rect 17902 12628 17914 12631
rect 18506 12628 18512 12640
rect 17902 12600 18512 12628
rect 17902 12597 17914 12600
rect 17856 12591 17914 12597
rect 18506 12588 18512 12600
rect 18564 12588 18570 12640
rect 19444 12637 19472 12668
rect 19429 12631 19487 12637
rect 19429 12597 19441 12631
rect 19475 12597 19487 12631
rect 19628 12628 19656 12727
rect 22738 12724 22744 12776
rect 22796 12764 22802 12776
rect 22922 12764 22928 12776
rect 22796 12736 22928 12764
rect 22796 12724 22802 12736
rect 22922 12724 22928 12736
rect 22980 12724 22986 12776
rect 24872 12764 24900 12804
rect 25038 12792 25044 12844
rect 25096 12832 25102 12844
rect 25777 12835 25835 12841
rect 25777 12832 25789 12835
rect 25096 12804 25789 12832
rect 25096 12792 25102 12804
rect 25777 12801 25789 12804
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 25884 12764 25912 12872
rect 33781 12869 33793 12872
rect 33827 12869 33839 12903
rect 33781 12863 33839 12869
rect 26234 12792 26240 12844
rect 26292 12832 26298 12844
rect 27433 12835 27491 12841
rect 27433 12832 27445 12835
rect 26292 12804 27445 12832
rect 26292 12792 26298 12804
rect 27433 12801 27445 12804
rect 27479 12832 27491 12835
rect 28350 12832 28356 12844
rect 27479 12804 28356 12832
rect 27479 12801 27491 12804
rect 27433 12795 27491 12801
rect 28350 12792 28356 12804
rect 28408 12832 28414 12844
rect 28810 12832 28816 12844
rect 28408 12804 28816 12832
rect 28408 12792 28414 12804
rect 28810 12792 28816 12804
rect 28868 12792 28874 12844
rect 31294 12792 31300 12844
rect 31352 12792 31358 12844
rect 24872 12736 25912 12764
rect 26142 12724 26148 12776
rect 26200 12764 26206 12776
rect 26605 12767 26663 12773
rect 26605 12764 26617 12767
rect 26200 12736 26617 12764
rect 26200 12724 26206 12736
rect 26605 12733 26617 12736
rect 26651 12733 26663 12767
rect 26605 12727 26663 12733
rect 27062 12724 27068 12776
rect 27120 12764 27126 12776
rect 27341 12767 27399 12773
rect 27341 12764 27353 12767
rect 27120 12736 27353 12764
rect 27120 12724 27126 12736
rect 27341 12733 27353 12736
rect 27387 12733 27399 12767
rect 27341 12727 27399 12733
rect 27893 12767 27951 12773
rect 27893 12733 27905 12767
rect 27939 12764 27951 12767
rect 27982 12764 27988 12776
rect 27939 12736 27988 12764
rect 27939 12733 27951 12736
rect 27893 12727 27951 12733
rect 27982 12724 27988 12736
rect 28040 12724 28046 12776
rect 29178 12724 29184 12776
rect 29236 12724 29242 12776
rect 29546 12724 29552 12776
rect 29604 12724 29610 12776
rect 30374 12724 30380 12776
rect 30432 12724 30438 12776
rect 33965 12767 34023 12773
rect 33965 12733 33977 12767
rect 34011 12764 34023 12767
rect 34422 12764 34428 12776
rect 34011 12736 34428 12764
rect 34011 12733 34023 12736
rect 33965 12727 34023 12733
rect 34422 12724 34428 12736
rect 34480 12724 34486 12776
rect 19978 12656 19984 12708
rect 20036 12696 20042 12708
rect 20438 12696 20444 12708
rect 20036 12668 20444 12696
rect 20036 12656 20042 12668
rect 20438 12656 20444 12668
rect 20496 12656 20502 12708
rect 21450 12656 21456 12708
rect 21508 12696 21514 12708
rect 21545 12699 21603 12705
rect 21545 12696 21557 12699
rect 21508 12668 21557 12696
rect 21508 12656 21514 12668
rect 21545 12665 21557 12668
rect 21591 12665 21603 12699
rect 21545 12659 21603 12665
rect 23750 12656 23756 12708
rect 23808 12656 23814 12708
rect 23934 12656 23940 12708
rect 23992 12696 23998 12708
rect 23992 12668 24150 12696
rect 23992 12656 23998 12668
rect 26510 12656 26516 12708
rect 26568 12696 26574 12708
rect 27249 12699 27307 12705
rect 27249 12696 27261 12699
rect 26568 12668 27261 12696
rect 26568 12656 26574 12668
rect 27249 12665 27261 12668
rect 27295 12696 27307 12699
rect 27522 12696 27528 12708
rect 27295 12668 27528 12696
rect 27295 12665 27307 12668
rect 27249 12659 27307 12665
rect 27522 12656 27528 12668
rect 27580 12656 27586 12708
rect 28074 12656 28080 12708
rect 28132 12656 28138 12708
rect 19886 12628 19892 12640
rect 19628 12600 19892 12628
rect 19429 12591 19487 12597
rect 19886 12588 19892 12600
rect 19944 12628 19950 12640
rect 23768 12628 23796 12656
rect 19944 12600 23796 12628
rect 19944 12588 19950 12600
rect 24302 12588 24308 12640
rect 24360 12628 24366 12640
rect 25225 12631 25283 12637
rect 25225 12628 25237 12631
rect 24360 12600 25237 12628
rect 24360 12588 24366 12600
rect 25225 12597 25237 12600
rect 25271 12597 25283 12631
rect 25225 12591 25283 12597
rect 26878 12588 26884 12640
rect 26936 12588 26942 12640
rect 30006 12588 30012 12640
rect 30064 12628 30070 12640
rect 30193 12631 30251 12637
rect 30193 12628 30205 12631
rect 30064 12600 30205 12628
rect 30064 12588 30070 12600
rect 30193 12597 30205 12600
rect 30239 12597 30251 12631
rect 30193 12591 30251 12597
rect 31021 12631 31079 12637
rect 31021 12597 31033 12631
rect 31067 12628 31079 12631
rect 31754 12628 31760 12640
rect 31067 12600 31760 12628
rect 31067 12597 31079 12600
rect 31021 12591 31079 12597
rect 31754 12588 31760 12600
rect 31812 12588 31818 12640
rect 2760 12538 34316 12560
rect 2760 12486 7210 12538
rect 7262 12486 7274 12538
rect 7326 12486 7338 12538
rect 7390 12486 7402 12538
rect 7454 12486 7466 12538
rect 7518 12486 15099 12538
rect 15151 12486 15163 12538
rect 15215 12486 15227 12538
rect 15279 12486 15291 12538
rect 15343 12486 15355 12538
rect 15407 12486 22988 12538
rect 23040 12486 23052 12538
rect 23104 12486 23116 12538
rect 23168 12486 23180 12538
rect 23232 12486 23244 12538
rect 23296 12486 30877 12538
rect 30929 12486 30941 12538
rect 30993 12486 31005 12538
rect 31057 12486 31069 12538
rect 31121 12486 31133 12538
rect 31185 12486 34316 12538
rect 2760 12464 34316 12486
rect 3605 12427 3663 12433
rect 3605 12393 3617 12427
rect 3651 12424 3663 12427
rect 3878 12424 3884 12436
rect 3651 12396 3884 12424
rect 3651 12393 3663 12396
rect 3605 12387 3663 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 5534 12424 5540 12436
rect 4019 12396 5540 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 6178 12424 6184 12436
rect 5920 12396 6184 12424
rect 5810 12356 5816 12368
rect 5474 12328 5816 12356
rect 5810 12316 5816 12328
rect 5868 12316 5874 12368
rect 5920 12365 5948 12396
rect 6178 12384 6184 12396
rect 6236 12384 6242 12436
rect 6825 12427 6883 12433
rect 6825 12393 6837 12427
rect 6871 12424 6883 12427
rect 7834 12424 7840 12436
rect 6871 12396 7840 12424
rect 6871 12393 6883 12396
rect 6825 12387 6883 12393
rect 7834 12384 7840 12396
rect 7892 12384 7898 12436
rect 11974 12384 11980 12436
rect 12032 12384 12038 12436
rect 12158 12384 12164 12436
rect 12216 12384 12222 12436
rect 12345 12427 12403 12433
rect 12345 12393 12357 12427
rect 12391 12424 12403 12427
rect 12618 12424 12624 12436
rect 12391 12396 12624 12424
rect 12391 12393 12403 12396
rect 12345 12387 12403 12393
rect 12618 12384 12624 12396
rect 12676 12384 12682 12436
rect 12894 12384 12900 12436
rect 12952 12384 12958 12436
rect 13170 12384 13176 12436
rect 13228 12384 13234 12436
rect 13446 12384 13452 12436
rect 13504 12424 13510 12436
rect 13541 12427 13599 12433
rect 13541 12424 13553 12427
rect 13504 12396 13553 12424
rect 13504 12384 13510 12396
rect 13541 12393 13553 12396
rect 13587 12393 13599 12427
rect 13541 12387 13599 12393
rect 13633 12427 13691 12433
rect 13633 12393 13645 12427
rect 13679 12424 13691 12427
rect 13814 12424 13820 12436
rect 13679 12396 13820 12424
rect 13679 12393 13691 12396
rect 13633 12387 13691 12393
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 14274 12384 14280 12436
rect 14332 12424 14338 12436
rect 14645 12427 14703 12433
rect 14645 12424 14657 12427
rect 14332 12396 14657 12424
rect 14332 12384 14338 12396
rect 14645 12393 14657 12396
rect 14691 12393 14703 12427
rect 17037 12427 17095 12433
rect 14645 12387 14703 12393
rect 14752 12396 16988 12424
rect 5905 12359 5963 12365
rect 5905 12325 5917 12359
rect 5951 12325 5963 12359
rect 5905 12319 5963 12325
rect 6546 12316 6552 12368
rect 6604 12316 6610 12368
rect 8570 12316 8576 12368
rect 8628 12356 8634 12368
rect 8665 12359 8723 12365
rect 8665 12356 8677 12359
rect 8628 12328 8677 12356
rect 8628 12316 8634 12328
rect 8665 12325 8677 12328
rect 8711 12325 8723 12359
rect 8665 12319 8723 12325
rect 10505 12359 10563 12365
rect 10505 12325 10517 12359
rect 10551 12356 10563 12359
rect 10778 12356 10784 12368
rect 10551 12328 10784 12356
rect 10551 12325 10563 12328
rect 10505 12319 10563 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 3329 12291 3387 12297
rect 3329 12257 3341 12291
rect 3375 12288 3387 12291
rect 3375 12260 4752 12288
rect 3375 12257 3387 12260
rect 3329 12251 3387 12257
rect 3970 12180 3976 12232
rect 4028 12180 4034 12232
rect 4062 12180 4068 12232
rect 4120 12180 4126 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4724 12220 4752 12260
rect 6178 12248 6184 12300
rect 6236 12248 6242 12300
rect 6362 12297 6368 12300
rect 6319 12291 6368 12297
rect 6319 12257 6331 12291
rect 6365 12257 6368 12291
rect 6319 12251 6368 12257
rect 6362 12248 6368 12251
rect 6420 12248 6426 12300
rect 6457 12291 6515 12297
rect 6457 12257 6469 12291
rect 6503 12286 6515 12291
rect 6665 12291 6723 12297
rect 6503 12258 6592 12286
rect 6503 12257 6515 12258
rect 6457 12251 6515 12257
rect 5166 12220 5172 12232
rect 4724 12192 5172 12220
rect 4157 12183 4215 12189
rect 3988 12152 4016 12180
rect 4172 12152 4200 12183
rect 5166 12180 5172 12192
rect 5224 12180 5230 12232
rect 5258 12180 5264 12232
rect 5316 12220 5322 12232
rect 6564 12220 6592 12258
rect 6665 12257 6677 12291
rect 6711 12288 6723 12291
rect 8202 12288 8208 12300
rect 6711 12260 6960 12288
rect 6711 12257 6723 12260
rect 6665 12251 6723 12257
rect 6822 12220 6828 12232
rect 5316 12192 6828 12220
rect 5316 12180 5322 12192
rect 6822 12180 6828 12192
rect 6880 12180 6886 12232
rect 3988 12124 4200 12152
rect 6932 12152 6960 12260
rect 7024 12260 8208 12288
rect 7024 12232 7052 12260
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 9766 12248 9772 12300
rect 9824 12248 9830 12300
rect 10226 12248 10232 12300
rect 10284 12248 10290 12300
rect 11606 12248 11612 12300
rect 11664 12248 11670 12300
rect 12176 12288 12204 12384
rect 14752 12356 14780 12396
rect 16114 12356 16120 12368
rect 12912 12328 14780 12356
rect 14844 12328 16120 12356
rect 12805 12291 12863 12297
rect 12805 12288 12817 12291
rect 12176 12260 12817 12288
rect 12805 12257 12817 12260
rect 12851 12257 12863 12291
rect 12805 12251 12863 12257
rect 7006 12180 7012 12232
rect 7064 12180 7070 12232
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 8389 12223 8447 12229
rect 8389 12220 8401 12223
rect 7708 12192 8401 12220
rect 7708 12180 7714 12192
rect 8389 12189 8401 12192
rect 8435 12189 8447 12223
rect 8389 12183 8447 12189
rect 10594 12180 10600 12232
rect 10652 12220 10658 12232
rect 12912 12220 12940 12328
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 14277 12291 14335 12297
rect 14277 12288 14289 12291
rect 13320 12260 14289 12288
rect 13320 12248 13326 12260
rect 14277 12257 14289 12260
rect 14323 12257 14335 12291
rect 14277 12251 14335 12257
rect 14642 12248 14648 12300
rect 14700 12248 14706 12300
rect 14844 12297 14872 12328
rect 16114 12316 16120 12328
rect 16172 12316 16178 12368
rect 16574 12356 16580 12368
rect 16500 12328 16580 12356
rect 14829 12291 14887 12297
rect 14829 12257 14841 12291
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 14921 12291 14979 12297
rect 14921 12257 14933 12291
rect 14967 12257 14979 12291
rect 14921 12251 14979 12257
rect 10652 12192 12940 12220
rect 10652 12180 10658 12192
rect 13722 12180 13728 12232
rect 13780 12180 13786 12232
rect 14936 12220 14964 12251
rect 15010 12248 15016 12300
rect 15068 12248 15074 12300
rect 16022 12288 16028 12300
rect 15304 12260 16028 12288
rect 14844 12192 14964 12220
rect 14844 12164 14872 12192
rect 6932 12124 8432 12152
rect 8404 12096 8432 12124
rect 14826 12112 14832 12164
rect 14884 12112 14890 12164
rect 15028 12152 15056 12248
rect 15304 12229 15332 12260
rect 16022 12248 16028 12260
rect 16080 12288 16086 12300
rect 16500 12297 16528 12328
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 16850 12316 16856 12368
rect 16908 12316 16914 12368
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 16080 12260 16497 12288
rect 16080 12248 16086 12260
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 15470 12180 15476 12232
rect 15528 12180 15534 12232
rect 15746 12180 15752 12232
rect 15804 12180 15810 12232
rect 15838 12180 15844 12232
rect 15896 12220 15902 12232
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 15896 12192 16313 12220
rect 15896 12180 15902 12192
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 16301 12183 16359 12189
rect 15086 12155 15144 12161
rect 15086 12152 15098 12155
rect 15028 12124 15098 12152
rect 15086 12121 15098 12124
rect 15132 12121 15144 12155
rect 15086 12115 15144 12121
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12152 15255 12155
rect 15562 12152 15568 12164
rect 15243 12124 15568 12152
rect 15243 12121 15255 12124
rect 15197 12115 15255 12121
rect 15562 12112 15568 12124
rect 15620 12152 15626 12164
rect 16868 12152 16896 12316
rect 16960 12288 16988 12396
rect 17037 12393 17049 12427
rect 17083 12424 17095 12427
rect 18785 12427 18843 12433
rect 17083 12396 17172 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 17144 12368 17172 12396
rect 17880 12396 18368 12424
rect 17880 12368 17908 12396
rect 17126 12316 17132 12368
rect 17184 12316 17190 12368
rect 17862 12316 17868 12368
rect 17920 12316 17926 12368
rect 18340 12365 18368 12396
rect 18785 12393 18797 12427
rect 18831 12424 18843 12427
rect 18966 12424 18972 12436
rect 18831 12396 18972 12424
rect 18831 12393 18843 12396
rect 18785 12387 18843 12393
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 19150 12384 19156 12436
rect 19208 12424 19214 12436
rect 19254 12427 19312 12433
rect 19254 12424 19266 12427
rect 19208 12396 19266 12424
rect 19208 12384 19214 12396
rect 19254 12393 19266 12396
rect 19300 12393 19312 12427
rect 19254 12387 19312 12393
rect 19518 12384 19524 12436
rect 19576 12424 19582 12436
rect 19797 12427 19855 12433
rect 19797 12424 19809 12427
rect 19576 12396 19809 12424
rect 19576 12384 19582 12396
rect 19797 12393 19809 12396
rect 19843 12393 19855 12427
rect 19797 12387 19855 12393
rect 19886 12384 19892 12436
rect 19944 12424 19950 12436
rect 19944 12396 20024 12424
rect 19944 12384 19950 12396
rect 18325 12359 18383 12365
rect 18325 12325 18337 12359
rect 18371 12325 18383 12359
rect 18325 12319 18383 12325
rect 18598 12316 18604 12368
rect 18656 12356 18662 12368
rect 18877 12359 18935 12365
rect 18877 12356 18889 12359
rect 18656 12328 18889 12356
rect 18656 12316 18662 12328
rect 18877 12325 18889 12328
rect 18923 12325 18935 12359
rect 18877 12319 18935 12325
rect 19518 12288 19524 12300
rect 16960 12260 19524 12288
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 19889 12291 19947 12297
rect 19889 12257 19901 12291
rect 19935 12288 19947 12291
rect 19996 12288 20024 12396
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 20990 12424 20996 12436
rect 20772 12396 20996 12424
rect 20772 12384 20778 12396
rect 20990 12384 20996 12396
rect 21048 12424 21054 12436
rect 21048 12396 21772 12424
rect 21048 12384 21054 12396
rect 19935 12260 20024 12288
rect 19935 12257 19947 12260
rect 19889 12251 19947 12257
rect 20898 12248 20904 12300
rect 20956 12248 20962 12300
rect 20990 12248 20996 12300
rect 21048 12288 21054 12300
rect 21744 12297 21772 12396
rect 23934 12384 23940 12436
rect 23992 12384 23998 12436
rect 25222 12424 25228 12436
rect 24412 12396 25228 12424
rect 23750 12356 23756 12368
rect 23492 12328 23756 12356
rect 23492 12297 23520 12328
rect 23750 12316 23756 12328
rect 23808 12356 23814 12368
rect 23808 12328 24164 12356
rect 23808 12316 23814 12328
rect 24136 12300 24164 12328
rect 21453 12291 21511 12297
rect 21048 12286 21404 12288
rect 21453 12286 21465 12291
rect 21048 12260 21465 12286
rect 21048 12248 21054 12260
rect 21376 12258 21465 12260
rect 21453 12257 21465 12258
rect 21499 12257 21511 12291
rect 21453 12251 21511 12257
rect 21729 12291 21787 12297
rect 21729 12257 21741 12291
rect 21775 12257 21787 12291
rect 21729 12251 21787 12257
rect 23477 12291 23535 12297
rect 23477 12257 23489 12291
rect 23523 12257 23535 12291
rect 23477 12251 23535 12257
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18104 12192 18736 12220
rect 18104 12180 18110 12192
rect 17218 12152 17224 12164
rect 15620 12124 15792 12152
rect 16868 12124 17224 12152
rect 15620 12112 15626 12124
rect 15764 12096 15792 12124
rect 17218 12112 17224 12124
rect 17276 12152 17282 12164
rect 18601 12155 18659 12161
rect 18601 12152 18613 12155
rect 17276 12124 18613 12152
rect 17276 12112 17282 12124
rect 18601 12121 18613 12124
rect 18647 12121 18659 12155
rect 18708 12152 18736 12192
rect 18874 12180 18880 12232
rect 18932 12220 18938 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 18932 12192 20269 12220
rect 18932 12180 18938 12192
rect 20257 12189 20269 12192
rect 20303 12220 20315 12223
rect 20806 12220 20812 12232
rect 20303 12192 20812 12220
rect 20303 12189 20315 12192
rect 20257 12183 20315 12189
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 21082 12180 21088 12232
rect 21140 12180 21146 12232
rect 21266 12152 21272 12164
rect 18708 12124 21272 12152
rect 18601 12115 18659 12121
rect 21266 12112 21272 12124
rect 21324 12112 21330 12164
rect 3418 12044 3424 12096
rect 3476 12044 3482 12096
rect 4430 12044 4436 12096
rect 4488 12044 4494 12096
rect 5902 12044 5908 12096
rect 5960 12084 5966 12096
rect 6546 12084 6552 12096
rect 5960 12056 6552 12084
rect 5960 12044 5966 12056
rect 6546 12044 6552 12056
rect 6604 12084 6610 12096
rect 6917 12087 6975 12093
rect 6917 12084 6929 12087
rect 6604 12056 6929 12084
rect 6604 12044 6610 12056
rect 6917 12053 6929 12056
rect 6963 12053 6975 12087
rect 6917 12047 6975 12053
rect 8110 12044 8116 12096
rect 8168 12044 8174 12096
rect 8386 12044 8392 12096
rect 8444 12044 8450 12096
rect 10134 12044 10140 12096
rect 10192 12044 10198 12096
rect 12710 12044 12716 12096
rect 12768 12044 12774 12096
rect 12894 12044 12900 12096
rect 12952 12084 12958 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 12952 12056 14381 12084
rect 12952 12044 12958 12056
rect 14369 12053 14381 12056
rect 14415 12084 14427 12087
rect 14918 12084 14924 12096
rect 14415 12056 14924 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15746 12044 15752 12096
rect 15804 12044 15810 12096
rect 16298 12044 16304 12096
rect 16356 12084 16362 12096
rect 16853 12087 16911 12093
rect 16853 12084 16865 12087
rect 16356 12056 16865 12084
rect 16356 12044 16362 12056
rect 16853 12053 16865 12056
rect 16899 12084 16911 12087
rect 17862 12084 17868 12096
rect 16899 12056 17868 12084
rect 16899 12053 16911 12056
rect 16853 12047 16911 12053
rect 17862 12044 17868 12056
rect 17920 12084 17926 12096
rect 18782 12084 18788 12096
rect 17920 12056 18788 12084
rect 17920 12044 17926 12056
rect 18782 12044 18788 12056
rect 18840 12084 18846 12096
rect 19245 12087 19303 12093
rect 19245 12084 19257 12087
rect 18840 12056 19257 12084
rect 18840 12044 18846 12056
rect 19245 12053 19257 12056
rect 19291 12053 19303 12087
rect 19245 12047 19303 12053
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 19978 12084 19984 12096
rect 19484 12056 19984 12084
rect 19484 12044 19490 12056
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 21542 12044 21548 12096
rect 21600 12084 21606 12096
rect 21744 12084 21772 12251
rect 23566 12248 23572 12300
rect 23624 12248 23630 12300
rect 23845 12291 23903 12297
rect 23845 12257 23857 12291
rect 23891 12257 23903 12291
rect 23845 12251 23903 12257
rect 22002 12180 22008 12232
rect 22060 12220 22066 12232
rect 22281 12223 22339 12229
rect 22281 12220 22293 12223
rect 22060 12192 22293 12220
rect 22060 12180 22066 12192
rect 22281 12189 22293 12192
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 22557 12223 22615 12229
rect 22557 12189 22569 12223
rect 22603 12220 22615 12223
rect 23584 12220 23612 12248
rect 22603 12192 23612 12220
rect 23860 12220 23888 12251
rect 24118 12248 24124 12300
rect 24176 12248 24182 12300
rect 24412 12297 24440 12396
rect 25222 12384 25228 12396
rect 25280 12384 25286 12436
rect 26237 12427 26295 12433
rect 26237 12393 26249 12427
rect 26283 12424 26295 12427
rect 26418 12424 26424 12436
rect 26283 12396 26424 12424
rect 26283 12393 26295 12396
rect 26237 12387 26295 12393
rect 26418 12384 26424 12396
rect 26476 12384 26482 12436
rect 26513 12427 26571 12433
rect 26513 12393 26525 12427
rect 26559 12424 26571 12427
rect 26694 12424 26700 12436
rect 26559 12396 26700 12424
rect 26559 12393 26571 12396
rect 26513 12387 26571 12393
rect 26694 12384 26700 12396
rect 26752 12384 26758 12436
rect 27890 12384 27896 12436
rect 27948 12424 27954 12436
rect 28629 12427 28687 12433
rect 28629 12424 28641 12427
rect 27948 12396 28641 12424
rect 27948 12384 27954 12396
rect 28629 12393 28641 12396
rect 28675 12393 28687 12427
rect 28902 12424 28908 12436
rect 28629 12387 28687 12393
rect 28736 12396 28908 12424
rect 26881 12359 26939 12365
rect 26881 12325 26893 12359
rect 26927 12356 26939 12359
rect 28736 12356 28764 12396
rect 28902 12384 28908 12396
rect 28960 12384 28966 12436
rect 29270 12384 29276 12436
rect 29328 12384 29334 12436
rect 29457 12427 29515 12433
rect 29457 12393 29469 12427
rect 29503 12424 29515 12427
rect 29546 12424 29552 12436
rect 29503 12396 29552 12424
rect 29503 12393 29515 12396
rect 29457 12387 29515 12393
rect 29546 12384 29552 12396
rect 29604 12384 29610 12436
rect 30098 12384 30104 12436
rect 30156 12424 30162 12436
rect 30285 12427 30343 12433
rect 30285 12424 30297 12427
rect 30156 12396 30297 12424
rect 30156 12384 30162 12396
rect 30285 12393 30297 12396
rect 30331 12393 30343 12427
rect 30285 12387 30343 12393
rect 33502 12384 33508 12436
rect 33560 12384 33566 12436
rect 26927 12328 28764 12356
rect 28813 12359 28871 12365
rect 26927 12325 26939 12328
rect 26881 12319 26939 12325
rect 28813 12325 28825 12359
rect 28859 12356 28871 12359
rect 29288 12356 29316 12384
rect 28859 12328 29316 12356
rect 28859 12325 28871 12328
rect 28813 12319 28871 12325
rect 24397 12291 24455 12297
rect 24397 12257 24409 12291
rect 24443 12257 24455 12291
rect 24397 12251 24455 12257
rect 24578 12248 24584 12300
rect 24636 12248 24642 12300
rect 26418 12288 26424 12300
rect 26160 12260 26424 12288
rect 24946 12220 24952 12232
rect 23860 12192 24952 12220
rect 22603 12189 22615 12192
rect 22557 12183 22615 12189
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 25314 12180 25320 12232
rect 25372 12180 25378 12232
rect 25498 12229 25504 12232
rect 25455 12223 25504 12229
rect 25455 12189 25467 12223
rect 25501 12189 25504 12223
rect 25455 12183 25504 12189
rect 25498 12180 25504 12183
rect 25556 12180 25562 12232
rect 25593 12223 25651 12229
rect 25593 12189 25605 12223
rect 25639 12220 25651 12223
rect 26160 12220 26188 12260
rect 26418 12248 26424 12260
rect 26476 12288 26482 12300
rect 26697 12291 26755 12297
rect 26697 12288 26709 12291
rect 26476 12260 26709 12288
rect 26476 12248 26482 12260
rect 26697 12257 26709 12260
rect 26743 12257 26755 12291
rect 26697 12251 26755 12257
rect 25639 12192 26188 12220
rect 25639 12189 25651 12192
rect 25593 12183 25651 12189
rect 26234 12180 26240 12232
rect 26292 12180 26298 12232
rect 26712 12220 26740 12251
rect 26970 12248 26976 12300
rect 27028 12248 27034 12300
rect 28994 12248 29000 12300
rect 29052 12248 29058 12300
rect 29196 12297 29224 12328
rect 29730 12316 29736 12368
rect 29788 12316 29794 12368
rect 29825 12359 29883 12365
rect 29825 12325 29837 12359
rect 29871 12356 29883 12359
rect 30006 12356 30012 12368
rect 29871 12328 30012 12356
rect 29871 12325 29883 12328
rect 29825 12319 29883 12325
rect 30006 12316 30012 12328
rect 30064 12316 30070 12368
rect 31294 12316 31300 12368
rect 31352 12316 31358 12368
rect 31754 12316 31760 12368
rect 31812 12316 31818 12368
rect 29181 12291 29239 12297
rect 29181 12257 29193 12291
rect 29227 12257 29239 12291
rect 29181 12251 29239 12257
rect 29270 12248 29276 12300
rect 29328 12248 29334 12300
rect 29549 12291 29607 12297
rect 29549 12257 29561 12291
rect 29595 12257 29607 12291
rect 29549 12251 29607 12257
rect 29917 12291 29975 12297
rect 29917 12257 29929 12291
rect 29963 12288 29975 12291
rect 32033 12291 32091 12297
rect 29963 12260 30604 12288
rect 29963 12257 29975 12260
rect 29917 12251 29975 12257
rect 27062 12220 27068 12232
rect 26712 12192 27068 12220
rect 27062 12180 27068 12192
rect 27120 12220 27126 12232
rect 29564 12220 29592 12251
rect 27120 12192 29960 12220
rect 27120 12180 27126 12192
rect 25041 12155 25099 12161
rect 25041 12121 25053 12155
rect 25087 12121 25099 12155
rect 25041 12115 25099 12121
rect 21600 12056 21772 12084
rect 21600 12044 21606 12056
rect 22738 12044 22744 12096
rect 22796 12084 22802 12096
rect 23382 12084 23388 12096
rect 22796 12056 23388 12084
rect 22796 12044 22802 12056
rect 23382 12044 23388 12056
rect 23440 12084 23446 12096
rect 23661 12087 23719 12093
rect 23661 12084 23673 12087
rect 23440 12056 23673 12084
rect 23440 12044 23446 12056
rect 23661 12053 23673 12056
rect 23707 12053 23719 12087
rect 25056 12084 25084 12115
rect 26252 12084 26280 12180
rect 29932 12164 29960 12192
rect 30374 12180 30380 12232
rect 30432 12180 30438 12232
rect 30576 12220 30604 12260
rect 32033 12257 32045 12291
rect 32079 12288 32091 12291
rect 32582 12288 32588 12300
rect 32079 12260 32588 12288
rect 32079 12257 32091 12260
rect 32033 12251 32091 12257
rect 32582 12248 32588 12260
rect 32640 12248 32646 12300
rect 31202 12220 31208 12232
rect 30576 12192 31208 12220
rect 31202 12180 31208 12192
rect 31260 12180 31266 12232
rect 32674 12180 32680 12232
rect 32732 12180 32738 12232
rect 29914 12112 29920 12164
rect 29972 12112 29978 12164
rect 30101 12155 30159 12161
rect 30101 12121 30113 12155
rect 30147 12152 30159 12155
rect 30392 12152 30420 12180
rect 30147 12124 30420 12152
rect 30147 12121 30159 12124
rect 30101 12115 30159 12121
rect 25056 12056 26280 12084
rect 23661 12047 23719 12053
rect 27062 12044 27068 12096
rect 27120 12044 27126 12096
rect 32122 12044 32128 12096
rect 32180 12044 32186 12096
rect 33042 12044 33048 12096
rect 33100 12044 33106 12096
rect 2760 11994 34316 12016
rect 2760 11942 6550 11994
rect 6602 11942 6614 11994
rect 6666 11942 6678 11994
rect 6730 11942 6742 11994
rect 6794 11942 6806 11994
rect 6858 11942 14439 11994
rect 14491 11942 14503 11994
rect 14555 11942 14567 11994
rect 14619 11942 14631 11994
rect 14683 11942 14695 11994
rect 14747 11942 22328 11994
rect 22380 11942 22392 11994
rect 22444 11942 22456 11994
rect 22508 11942 22520 11994
rect 22572 11942 22584 11994
rect 22636 11942 30217 11994
rect 30269 11942 30281 11994
rect 30333 11942 30345 11994
rect 30397 11942 30409 11994
rect 30461 11942 30473 11994
rect 30525 11942 34316 11994
rect 2760 11920 34316 11942
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 4062 11880 4068 11892
rect 3099 11852 4068 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 5166 11840 5172 11892
rect 5224 11840 5230 11892
rect 5258 11840 5264 11892
rect 5316 11840 5322 11892
rect 5445 11883 5503 11889
rect 5445 11849 5457 11883
rect 5491 11880 5503 11883
rect 5718 11880 5724 11892
rect 5491 11852 5724 11880
rect 5491 11849 5503 11852
rect 5445 11843 5503 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 5868 11852 6377 11880
rect 5868 11840 5874 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6733 11883 6791 11889
rect 6733 11849 6745 11883
rect 6779 11880 6791 11883
rect 7466 11880 7472 11892
rect 6779 11852 7472 11880
rect 6779 11849 6791 11852
rect 6733 11843 6791 11849
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 8386 11840 8392 11892
rect 8444 11880 8450 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8444 11852 8769 11880
rect 8444 11840 8450 11852
rect 8757 11849 8769 11852
rect 8803 11880 8815 11883
rect 8938 11880 8944 11892
rect 8803 11852 8944 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 9585 11883 9643 11889
rect 9585 11849 9597 11883
rect 9631 11880 9643 11883
rect 9766 11880 9772 11892
rect 9631 11852 9772 11880
rect 9631 11849 9643 11852
rect 9585 11843 9643 11849
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12526 11880 12532 11892
rect 12483 11852 12532 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 12710 11840 12716 11892
rect 12768 11880 12774 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 12768 11852 13001 11880
rect 12768 11840 12774 11852
rect 12989 11849 13001 11852
rect 13035 11849 13047 11883
rect 12989 11843 13047 11849
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 13412 11852 14105 11880
rect 13412 11840 13418 11852
rect 14093 11849 14105 11852
rect 14139 11849 14151 11883
rect 14093 11843 14151 11849
rect 14369 11883 14427 11889
rect 14369 11849 14381 11883
rect 14415 11880 14427 11883
rect 14826 11880 14832 11892
rect 14415 11852 14832 11880
rect 14415 11849 14427 11852
rect 14369 11843 14427 11849
rect 14826 11840 14832 11852
rect 14884 11840 14890 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15562 11880 15568 11892
rect 15252 11852 15568 11880
rect 15252 11840 15258 11852
rect 15562 11840 15568 11852
rect 15620 11880 15626 11892
rect 15620 11852 17540 11880
rect 15620 11840 15626 11852
rect 5184 11812 5212 11840
rect 7006 11812 7012 11824
rect 5184 11784 7012 11812
rect 4522 11704 4528 11756
rect 4580 11704 4586 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5592 11716 6009 11744
rect 5592 11704 5598 11716
rect 5997 11713 6009 11716
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 3418 11636 3424 11688
rect 3476 11636 3482 11688
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11676 4859 11679
rect 6178 11676 6184 11688
rect 4847 11648 6184 11676
rect 4847 11645 4859 11648
rect 4801 11639 4859 11645
rect 4816 11608 4844 11639
rect 6178 11636 6184 11648
rect 6236 11636 6242 11688
rect 6472 11685 6500 11784
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 10134 11772 10140 11824
rect 10192 11772 10198 11824
rect 12805 11815 12863 11821
rect 12805 11781 12817 11815
rect 12851 11812 12863 11815
rect 13096 11812 13124 11840
rect 15749 11815 15807 11821
rect 15749 11812 15761 11815
rect 12851 11784 13124 11812
rect 13188 11784 15761 11812
rect 12851 11781 12863 11784
rect 12805 11775 12863 11781
rect 7650 11704 7656 11756
rect 7708 11744 7714 11756
rect 8481 11747 8539 11753
rect 8481 11744 8493 11747
rect 7708 11716 8493 11744
rect 7708 11704 7714 11716
rect 8481 11713 8493 11716
rect 8527 11713 8539 11747
rect 10152 11744 10180 11772
rect 10152 11716 13032 11744
rect 8481 11707 8539 11713
rect 6457 11679 6515 11685
rect 6457 11645 6469 11679
rect 6503 11645 6515 11679
rect 6457 11639 6515 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 10042 11676 10048 11688
rect 9723 11648 10048 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 10042 11636 10048 11648
rect 10100 11636 10106 11688
rect 11146 11636 11152 11688
rect 11204 11676 11210 11688
rect 11514 11676 11520 11688
rect 11204 11648 11520 11676
rect 11204 11636 11210 11648
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 11664 11648 11989 11676
rect 11664 11636 11670 11648
rect 11977 11645 11989 11648
rect 12023 11676 12035 11679
rect 12894 11676 12900 11688
rect 12023 11648 12900 11676
rect 12023 11645 12035 11648
rect 11977 11639 12035 11645
rect 12894 11636 12900 11648
rect 12952 11636 12958 11688
rect 4632 11580 4844 11608
rect 4632 11552 4660 11580
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 5905 11611 5963 11617
rect 5905 11608 5917 11611
rect 5500 11580 5917 11608
rect 5500 11568 5506 11580
rect 5905 11577 5917 11580
rect 5951 11577 5963 11611
rect 5905 11571 5963 11577
rect 6914 11568 6920 11620
rect 6972 11568 6978 11620
rect 8110 11608 8116 11620
rect 7774 11580 8116 11608
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 8205 11611 8263 11617
rect 8205 11577 8217 11611
rect 8251 11608 8263 11611
rect 8478 11608 8484 11620
rect 8251 11580 8484 11608
rect 8251 11577 8263 11580
rect 8205 11571 8263 11577
rect 8478 11568 8484 11580
rect 8536 11568 8542 11620
rect 12158 11608 12164 11620
rect 9646 11580 12164 11608
rect 4614 11500 4620 11552
rect 4672 11500 4678 11552
rect 5810 11500 5816 11552
rect 5868 11500 5874 11552
rect 6932 11540 6960 11568
rect 9646 11540 9674 11580
rect 12158 11568 12164 11580
rect 12216 11568 12222 11620
rect 6932 11512 9674 11540
rect 10778 11500 10784 11552
rect 10836 11540 10842 11552
rect 10962 11540 10968 11552
rect 10836 11512 10968 11540
rect 10836 11500 10842 11512
rect 10962 11500 10968 11512
rect 11020 11540 11026 11552
rect 11241 11543 11299 11549
rect 11241 11540 11253 11543
rect 11020 11512 11253 11540
rect 11020 11500 11026 11512
rect 11241 11509 11253 11512
rect 11287 11540 11299 11543
rect 12894 11540 12900 11552
rect 11287 11512 12900 11540
rect 11287 11509 11299 11512
rect 11241 11503 11299 11509
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13004 11540 13032 11716
rect 13188 11685 13216 11784
rect 15749 11781 15761 11784
rect 15795 11812 15807 11815
rect 15838 11812 15844 11824
rect 15795 11784 15844 11812
rect 15795 11781 15807 11784
rect 15749 11775 15807 11781
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 16298 11812 16304 11824
rect 16132 11784 16304 11812
rect 13446 11704 13452 11756
rect 13504 11704 13510 11756
rect 14182 11704 14188 11756
rect 14240 11744 14246 11756
rect 14240 11716 14504 11744
rect 14240 11704 14246 11716
rect 14476 11685 14504 11716
rect 15010 11704 15016 11756
rect 15068 11704 15074 11756
rect 15194 11704 15200 11756
rect 15252 11704 15258 11756
rect 15654 11704 15660 11756
rect 15712 11744 15718 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 15712 11716 15945 11744
rect 15712 11704 15718 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 16022 11704 16028 11756
rect 16080 11704 16086 11756
rect 16132 11753 16160 11784
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 16577 11815 16635 11821
rect 16577 11781 16589 11815
rect 16623 11812 16635 11815
rect 17313 11815 17371 11821
rect 17313 11812 17325 11815
rect 16623 11784 17325 11812
rect 16623 11781 16635 11784
rect 16577 11775 16635 11781
rect 17313 11781 17325 11784
rect 17359 11812 17371 11815
rect 17402 11812 17408 11824
rect 17359 11784 17408 11812
rect 17359 11781 17371 11784
rect 17313 11775 17371 11781
rect 16117 11747 16175 11753
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11676 13415 11679
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 13403 11648 14289 11676
rect 13403 11645 13415 11648
rect 13357 11639 13415 11645
rect 14277 11645 14289 11648
rect 14323 11645 14335 11679
rect 14277 11639 14335 11645
rect 14461 11679 14519 11685
rect 14461 11645 14473 11679
rect 14507 11645 14519 11679
rect 15028 11676 15056 11704
rect 14461 11639 14519 11645
rect 14568 11648 15056 11676
rect 15565 11679 15623 11685
rect 14292 11608 14320 11639
rect 14568 11608 14596 11648
rect 15565 11645 15577 11679
rect 15611 11676 15623 11679
rect 16592 11676 16620 11775
rect 17402 11772 17408 11784
rect 17460 11772 17466 11824
rect 17512 11812 17540 11852
rect 18506 11840 18512 11892
rect 18564 11840 18570 11892
rect 18690 11840 18696 11892
rect 18748 11840 18754 11892
rect 19242 11840 19248 11892
rect 19300 11880 19306 11892
rect 19334 11880 19340 11892
rect 19300 11852 19340 11880
rect 19300 11840 19306 11852
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 20714 11880 20720 11892
rect 19444 11852 20720 11880
rect 19444 11812 19472 11852
rect 20714 11840 20720 11852
rect 20772 11840 20778 11892
rect 21361 11883 21419 11889
rect 21361 11849 21373 11883
rect 21407 11880 21419 11883
rect 21910 11880 21916 11892
rect 21407 11852 21916 11880
rect 21407 11849 21419 11852
rect 21361 11843 21419 11849
rect 21910 11840 21916 11852
rect 21968 11840 21974 11892
rect 22646 11840 22652 11892
rect 22704 11840 22710 11892
rect 27062 11889 27068 11892
rect 27052 11883 27068 11889
rect 27052 11849 27064 11883
rect 27052 11843 27068 11849
rect 27062 11840 27068 11843
rect 27120 11840 27126 11892
rect 28537 11883 28595 11889
rect 28537 11849 28549 11883
rect 28583 11880 28595 11883
rect 29270 11880 29276 11892
rect 28583 11852 29276 11880
rect 28583 11849 28595 11852
rect 28537 11843 28595 11849
rect 29270 11840 29276 11852
rect 29328 11840 29334 11892
rect 31294 11840 31300 11892
rect 31352 11840 31358 11892
rect 31938 11840 31944 11892
rect 31996 11840 32002 11892
rect 32125 11883 32183 11889
rect 32125 11849 32137 11883
rect 32171 11880 32183 11883
rect 32674 11880 32680 11892
rect 32171 11852 32680 11880
rect 32171 11849 32183 11852
rect 32125 11843 32183 11849
rect 32674 11840 32680 11852
rect 32732 11840 32738 11892
rect 17512 11784 19472 11812
rect 25685 11815 25743 11821
rect 25685 11781 25697 11815
rect 25731 11812 25743 11815
rect 26050 11812 26056 11824
rect 25731 11784 26056 11812
rect 25731 11781 25743 11784
rect 25685 11775 25743 11781
rect 26050 11772 26056 11784
rect 26108 11772 26114 11824
rect 26418 11772 26424 11824
rect 26476 11772 26482 11824
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11744 17003 11747
rect 17034 11744 17040 11756
rect 16991 11716 17040 11744
rect 16991 11713 17003 11716
rect 16945 11707 17003 11713
rect 17034 11704 17040 11716
rect 17092 11704 17098 11756
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11744 18843 11747
rect 19150 11744 19156 11756
rect 18831 11716 19156 11744
rect 18831 11713 18843 11716
rect 18785 11707 18843 11713
rect 19150 11704 19156 11716
rect 19208 11704 19214 11756
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11744 19395 11747
rect 19383 11716 21680 11744
rect 19383 11713 19395 11716
rect 19337 11707 19395 11713
rect 15611 11648 16620 11676
rect 17129 11679 17187 11685
rect 15611 11645 15623 11648
rect 15565 11639 15623 11645
rect 17129 11645 17141 11679
rect 17175 11676 17187 11679
rect 17218 11676 17224 11688
rect 17175 11648 17224 11676
rect 17175 11645 17187 11648
rect 17129 11639 17187 11645
rect 17218 11636 17224 11648
rect 17276 11636 17282 11688
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11676 18935 11679
rect 18966 11676 18972 11688
rect 18923 11648 18972 11676
rect 18923 11645 18935 11648
rect 18877 11639 18935 11645
rect 18966 11636 18972 11648
rect 19024 11636 19030 11688
rect 19426 11636 19432 11688
rect 19484 11636 19490 11688
rect 19610 11636 19616 11688
rect 19668 11636 19674 11688
rect 19334 11608 19340 11620
rect 14292 11580 14596 11608
rect 14844 11580 19340 11608
rect 14844 11540 14872 11580
rect 19334 11568 19340 11580
rect 19392 11568 19398 11620
rect 13004 11512 14872 11540
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 17681 11543 17739 11549
rect 17681 11540 17693 11543
rect 17552 11512 17693 11540
rect 17552 11500 17558 11512
rect 17681 11509 17693 11512
rect 17727 11509 17739 11543
rect 17681 11503 17739 11509
rect 19150 11500 19156 11552
rect 19208 11540 19214 11552
rect 19720 11540 19748 11716
rect 21652 11688 21680 11716
rect 22830 11704 22836 11756
rect 22888 11744 22894 11756
rect 22925 11747 22983 11753
rect 22925 11744 22937 11747
rect 22888 11716 22937 11744
rect 22888 11704 22894 11716
rect 22925 11713 22937 11716
rect 22971 11713 22983 11747
rect 22925 11707 22983 11713
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11744 23259 11747
rect 24210 11744 24216 11756
rect 23247 11716 24216 11744
rect 23247 11713 23259 11716
rect 23201 11707 23259 11713
rect 24210 11704 24216 11716
rect 24268 11704 24274 11756
rect 26436 11744 26464 11772
rect 25700 11716 26464 11744
rect 26789 11747 26847 11753
rect 19886 11636 19892 11688
rect 19944 11676 19950 11688
rect 20073 11679 20131 11685
rect 20073 11676 20085 11679
rect 19944 11648 20085 11676
rect 19944 11636 19950 11648
rect 20073 11645 20085 11648
rect 20119 11676 20131 11679
rect 20898 11676 20904 11688
rect 20119 11648 20904 11676
rect 20119 11645 20131 11648
rect 20073 11639 20131 11645
rect 20898 11636 20904 11648
rect 20956 11676 20962 11688
rect 20993 11679 21051 11685
rect 20993 11676 21005 11679
rect 20956 11648 21005 11676
rect 20956 11636 20962 11648
rect 20993 11645 21005 11648
rect 21039 11645 21051 11679
rect 20993 11639 21051 11645
rect 21634 11636 21640 11688
rect 21692 11636 21698 11688
rect 21821 11679 21879 11685
rect 21821 11645 21833 11679
rect 21867 11676 21879 11679
rect 22094 11676 22100 11688
rect 21867 11648 22100 11676
rect 21867 11645 21879 11648
rect 21821 11639 21879 11645
rect 19208 11512 19748 11540
rect 19208 11500 19214 11512
rect 20530 11500 20536 11552
rect 20588 11540 20594 11552
rect 20717 11543 20775 11549
rect 20717 11540 20729 11543
rect 20588 11512 20729 11540
rect 20588 11500 20594 11512
rect 20717 11509 20729 11512
rect 20763 11509 20775 11543
rect 20717 11503 20775 11509
rect 20806 11500 20812 11552
rect 20864 11540 20870 11552
rect 21836 11540 21864 11639
rect 22094 11636 22100 11648
rect 22152 11636 22158 11688
rect 24946 11636 24952 11688
rect 25004 11636 25010 11688
rect 25700 11685 25728 11716
rect 26789 11713 26801 11747
rect 26835 11744 26847 11747
rect 27798 11744 27804 11756
rect 26835 11716 27804 11744
rect 26835 11713 26847 11716
rect 26789 11707 26847 11713
rect 27798 11704 27804 11716
rect 27856 11704 27862 11756
rect 28258 11704 28264 11756
rect 28316 11744 28322 11756
rect 32769 11747 32827 11753
rect 28316 11716 31984 11744
rect 28316 11704 28322 11716
rect 25685 11679 25743 11685
rect 25685 11645 25697 11679
rect 25731 11645 25743 11679
rect 25685 11639 25743 11645
rect 25869 11679 25927 11685
rect 25869 11645 25881 11679
rect 25915 11676 25927 11679
rect 26602 11676 26608 11688
rect 25915 11648 26608 11676
rect 25915 11645 25927 11648
rect 25869 11639 25927 11645
rect 26602 11636 26608 11648
rect 26660 11636 26666 11688
rect 28166 11636 28172 11688
rect 28224 11636 28230 11688
rect 29178 11636 29184 11688
rect 29236 11636 29242 11688
rect 30561 11679 30619 11685
rect 30561 11645 30573 11679
rect 30607 11676 30619 11679
rect 30650 11676 30656 11688
rect 30607 11648 30656 11676
rect 30607 11645 30619 11648
rect 30561 11639 30619 11645
rect 30650 11636 30656 11648
rect 30708 11636 30714 11688
rect 31389 11679 31447 11685
rect 31389 11676 31401 11679
rect 31220 11648 31401 11676
rect 24857 11611 24915 11617
rect 24857 11608 24869 11611
rect 24426 11580 24869 11608
rect 24857 11577 24869 11580
rect 24903 11577 24915 11611
rect 24857 11571 24915 11577
rect 26142 11568 26148 11620
rect 26200 11568 26206 11620
rect 28902 11568 28908 11620
rect 28960 11608 28966 11620
rect 29917 11611 29975 11617
rect 29917 11608 29929 11611
rect 28960 11580 29929 11608
rect 28960 11568 28966 11580
rect 29917 11577 29929 11580
rect 29963 11577 29975 11611
rect 29917 11571 29975 11577
rect 20864 11512 21864 11540
rect 24673 11543 24731 11549
rect 20864 11500 20870 11512
rect 24673 11509 24685 11543
rect 24719 11540 24731 11543
rect 26160 11540 26188 11568
rect 31220 11552 31248 11648
rect 31389 11645 31401 11648
rect 31435 11645 31447 11679
rect 31956 11676 31984 11716
rect 32769 11713 32781 11747
rect 32815 11744 32827 11747
rect 33502 11744 33508 11756
rect 32815 11716 33508 11744
rect 32815 11713 32827 11716
rect 32769 11707 32827 11713
rect 33502 11704 33508 11716
rect 33560 11704 33566 11756
rect 33042 11676 33048 11688
rect 31956 11648 33048 11676
rect 31389 11639 31447 11645
rect 33042 11636 33048 11648
rect 33100 11636 33106 11688
rect 31938 11568 31944 11620
rect 31996 11608 32002 11620
rect 32493 11611 32551 11617
rect 32493 11608 32505 11611
rect 31996 11580 32505 11608
rect 31996 11568 32002 11580
rect 32493 11577 32505 11580
rect 32539 11577 32551 11611
rect 32493 11571 32551 11577
rect 24719 11512 26188 11540
rect 24719 11509 24731 11512
rect 24673 11503 24731 11509
rect 29638 11500 29644 11552
rect 29696 11540 29702 11552
rect 29825 11543 29883 11549
rect 29825 11540 29837 11543
rect 29696 11512 29837 11540
rect 29696 11500 29702 11512
rect 29825 11509 29837 11512
rect 29871 11509 29883 11543
rect 29825 11503 29883 11509
rect 31202 11500 31208 11552
rect 31260 11500 31266 11552
rect 32582 11500 32588 11552
rect 32640 11500 32646 11552
rect 2760 11450 34316 11472
rect 2760 11398 7210 11450
rect 7262 11398 7274 11450
rect 7326 11398 7338 11450
rect 7390 11398 7402 11450
rect 7454 11398 7466 11450
rect 7518 11398 15099 11450
rect 15151 11398 15163 11450
rect 15215 11398 15227 11450
rect 15279 11398 15291 11450
rect 15343 11398 15355 11450
rect 15407 11398 22988 11450
rect 23040 11398 23052 11450
rect 23104 11398 23116 11450
rect 23168 11398 23180 11450
rect 23232 11398 23244 11450
rect 23296 11398 30877 11450
rect 30929 11398 30941 11450
rect 30993 11398 31005 11450
rect 31057 11398 31069 11450
rect 31121 11398 31133 11450
rect 31185 11398 34316 11450
rect 2760 11376 34316 11398
rect 4890 11296 4896 11348
rect 4948 11336 4954 11348
rect 4948 11308 7788 11336
rect 4948 11296 4954 11308
rect 1302 11228 1308 11280
rect 1360 11268 1366 11280
rect 3237 11271 3295 11277
rect 3237 11268 3249 11271
rect 1360 11240 3249 11268
rect 1360 11228 1366 11240
rect 3237 11237 3249 11240
rect 3283 11237 3295 11271
rect 3237 11231 3295 11237
rect 4430 11160 4436 11212
rect 4488 11160 4494 11212
rect 5460 11209 5488 11308
rect 7760 11280 7788 11308
rect 8294 11296 8300 11348
rect 8352 11336 8358 11348
rect 8849 11339 8907 11345
rect 8849 11336 8861 11339
rect 8352 11308 8861 11336
rect 8352 11296 8358 11308
rect 8849 11305 8861 11308
rect 8895 11305 8907 11339
rect 8849 11299 8907 11305
rect 9950 11296 9956 11348
rect 10008 11296 10014 11348
rect 10962 11296 10968 11348
rect 11020 11336 11026 11348
rect 11333 11339 11391 11345
rect 11333 11336 11345 11339
rect 11020 11308 11345 11336
rect 11020 11296 11026 11308
rect 11333 11305 11345 11308
rect 11379 11336 11391 11339
rect 11379 11308 12480 11336
rect 11379 11305 11391 11308
rect 11333 11299 11391 11305
rect 6086 11228 6092 11280
rect 6144 11228 6150 11280
rect 6178 11228 6184 11280
rect 6236 11268 6242 11280
rect 7374 11268 7380 11280
rect 6236 11240 7380 11268
rect 6236 11228 6242 11240
rect 7374 11228 7380 11240
rect 7432 11268 7438 11280
rect 7650 11268 7656 11280
rect 7432 11240 7656 11268
rect 7432 11228 7438 11240
rect 7650 11228 7656 11240
rect 7708 11228 7714 11280
rect 7742 11228 7748 11280
rect 7800 11228 7806 11280
rect 9858 11228 9864 11280
rect 9916 11228 9922 11280
rect 9968 11268 9996 11296
rect 11149 11271 11207 11277
rect 11149 11268 11161 11271
rect 9968 11240 11161 11268
rect 11149 11237 11161 11240
rect 11195 11237 11207 11271
rect 11149 11231 11207 11237
rect 5445 11203 5503 11209
rect 5445 11169 5457 11203
rect 5491 11169 5503 11203
rect 5445 11163 5503 11169
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 3970 11024 3976 11076
rect 4028 11064 4034 11076
rect 6104 11064 6132 11228
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 8573 11203 8631 11209
rect 8573 11200 8585 11203
rect 6972 11172 8585 11200
rect 6972 11160 6978 11172
rect 8573 11169 8585 11172
rect 8619 11169 8631 11203
rect 8573 11163 8631 11169
rect 10778 11160 10784 11212
rect 10836 11160 10842 11212
rect 12452 11209 12480 11308
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 13412 11308 13645 11336
rect 13412 11296 13418 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 13722 11296 13728 11348
rect 13780 11296 13786 11348
rect 15562 11336 15568 11348
rect 14844 11308 15568 11336
rect 12618 11228 12624 11280
rect 12676 11268 12682 11280
rect 12989 11271 13047 11277
rect 12989 11268 13001 11271
rect 12676 11240 13001 11268
rect 12676 11228 12682 11240
rect 12989 11237 13001 11240
rect 13035 11268 13047 11271
rect 13740 11268 13768 11296
rect 13035 11240 13768 11268
rect 13035 11237 13047 11240
rect 12989 11231 13047 11237
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 12526 11160 12532 11212
rect 12584 11160 12590 11212
rect 13078 11160 13084 11212
rect 13136 11200 13142 11212
rect 13541 11203 13599 11209
rect 13541 11200 13553 11203
rect 13136 11172 13553 11200
rect 13136 11160 13142 11172
rect 13541 11169 13553 11172
rect 13587 11169 13599 11203
rect 13541 11163 13599 11169
rect 13648 11172 13860 11200
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 8021 11135 8079 11141
rect 8021 11132 8033 11135
rect 6328 11104 8033 11132
rect 6328 11092 6334 11104
rect 8021 11101 8033 11104
rect 8067 11101 8079 11135
rect 8021 11095 8079 11101
rect 10318 11092 10324 11144
rect 10376 11092 10382 11144
rect 10594 11092 10600 11144
rect 10652 11092 10658 11144
rect 11330 11092 11336 11144
rect 11388 11132 11394 11144
rect 12069 11135 12127 11141
rect 12069 11132 12081 11135
rect 11388 11104 12081 11132
rect 11388 11092 11394 11104
rect 12069 11101 12081 11104
rect 12115 11101 12127 11135
rect 12069 11095 12127 11101
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 13648 11132 13676 11172
rect 12952 11104 13676 11132
rect 12952 11092 12958 11104
rect 13722 11092 13728 11144
rect 13780 11092 13786 11144
rect 13832 11132 13860 11172
rect 14182 11160 14188 11212
rect 14240 11160 14246 11212
rect 14734 11160 14740 11212
rect 14792 11200 14798 11212
rect 14844 11200 14872 11308
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 15838 11296 15844 11348
rect 15896 11336 15902 11348
rect 15896 11308 17724 11336
rect 15896 11296 15902 11308
rect 15930 11268 15936 11280
rect 15212 11240 15936 11268
rect 15212 11209 15240 11240
rect 15930 11228 15936 11240
rect 15988 11268 15994 11280
rect 16301 11271 16359 11277
rect 16301 11268 16313 11271
rect 15988 11240 16313 11268
rect 15988 11228 15994 11240
rect 16301 11237 16313 11240
rect 16347 11237 16359 11271
rect 16301 11231 16359 11237
rect 16666 11228 16672 11280
rect 16724 11228 16730 11280
rect 16761 11271 16819 11277
rect 16761 11237 16773 11271
rect 16807 11268 16819 11271
rect 16807 11240 17540 11268
rect 16807 11237 16819 11240
rect 16761 11231 16819 11237
rect 17512 11212 17540 11240
rect 14792 11172 14872 11200
rect 15197 11203 15255 11209
rect 14792 11160 14798 11172
rect 15197 11169 15209 11203
rect 15243 11169 15255 11203
rect 15197 11163 15255 11169
rect 16853 11203 16911 11209
rect 16853 11169 16865 11203
rect 16899 11200 16911 11203
rect 17402 11200 17408 11212
rect 16899 11172 17408 11200
rect 16899 11169 16911 11172
rect 16853 11163 16911 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17494 11160 17500 11212
rect 17552 11160 17558 11212
rect 17586 11160 17592 11212
rect 17644 11160 17650 11212
rect 17696 11209 17724 11308
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 19245 11339 19303 11345
rect 19245 11336 19257 11339
rect 18380 11308 19257 11336
rect 18380 11296 18386 11308
rect 19245 11305 19257 11308
rect 19291 11305 19303 11339
rect 19245 11299 19303 11305
rect 19978 11296 19984 11348
rect 20036 11296 20042 11348
rect 20990 11296 20996 11348
rect 21048 11296 21054 11348
rect 22922 11296 22928 11348
rect 22980 11336 22986 11348
rect 23382 11336 23388 11348
rect 22980 11308 23388 11336
rect 22980 11296 22986 11308
rect 23382 11296 23388 11308
rect 23440 11296 23446 11348
rect 26053 11339 26111 11345
rect 26053 11305 26065 11339
rect 26099 11336 26111 11339
rect 26326 11336 26332 11348
rect 26099 11308 26332 11336
rect 26099 11305 26111 11308
rect 26053 11299 26111 11305
rect 26326 11296 26332 11308
rect 26384 11296 26390 11348
rect 28166 11296 28172 11348
rect 28224 11296 28230 11348
rect 28997 11339 29055 11345
rect 28997 11305 29009 11339
rect 29043 11336 29055 11339
rect 29178 11336 29184 11348
rect 29043 11308 29184 11336
rect 29043 11305 29055 11308
rect 28997 11299 29055 11305
rect 29178 11296 29184 11308
rect 29236 11296 29242 11348
rect 30650 11296 30656 11348
rect 30708 11336 30714 11348
rect 30837 11339 30895 11345
rect 30837 11336 30849 11339
rect 30708 11308 30849 11336
rect 30708 11296 30714 11308
rect 30837 11305 30849 11308
rect 30883 11305 30895 11339
rect 30837 11299 30895 11305
rect 30926 11296 30932 11348
rect 30984 11336 30990 11348
rect 30984 11308 34008 11336
rect 30984 11296 30990 11308
rect 19705 11271 19763 11277
rect 17880 11240 19472 11268
rect 17880 11209 17908 11240
rect 19444 11212 19472 11240
rect 19705 11237 19717 11271
rect 19751 11268 19763 11271
rect 21008 11268 21036 11296
rect 19751 11240 21036 11268
rect 22373 11271 22431 11277
rect 19751 11237 19763 11240
rect 19705 11231 19763 11237
rect 17681 11203 17739 11209
rect 17681 11169 17693 11203
rect 17727 11169 17739 11203
rect 17681 11163 17739 11169
rect 17865 11203 17923 11209
rect 17865 11169 17877 11203
rect 17911 11169 17923 11203
rect 17865 11163 17923 11169
rect 19153 11203 19211 11209
rect 19153 11169 19165 11203
rect 19199 11169 19211 11203
rect 19153 11163 19211 11169
rect 19337 11203 19395 11209
rect 19337 11169 19349 11203
rect 19383 11169 19395 11203
rect 19337 11163 19395 11169
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 13832 11104 16129 11132
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 11606 11064 11612 11076
rect 4028 11036 6040 11064
rect 6104 11036 8248 11064
rect 4028 11024 4034 11036
rect 4706 10956 4712 11008
rect 4764 10996 4770 11008
rect 5534 10996 5540 11008
rect 4764 10968 5540 10996
rect 4764 10956 4770 10968
rect 5534 10956 5540 10968
rect 5592 10996 5598 11008
rect 5905 10999 5963 11005
rect 5905 10996 5917 10999
rect 5592 10968 5917 10996
rect 5592 10956 5598 10968
rect 5905 10965 5917 10968
rect 5951 10965 5963 10999
rect 6012 10996 6040 11036
rect 7650 10996 7656 11008
rect 6012 10968 7656 10996
rect 5905 10959 5963 10965
rect 7650 10956 7656 10968
rect 7708 10956 7714 11008
rect 8220 10996 8248 11036
rect 11072 11036 11612 11064
rect 8294 10996 8300 11008
rect 8220 10968 8300 10996
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 9674 10956 9680 11008
rect 9732 10996 9738 11008
rect 11072 10996 11100 11036
rect 11606 11024 11612 11036
rect 11664 11064 11670 11076
rect 12253 11067 12311 11073
rect 12253 11064 12265 11067
rect 11664 11036 12265 11064
rect 11664 11024 11670 11036
rect 12253 11033 12265 11036
rect 12299 11033 12311 11067
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 12253 11027 12311 11033
rect 13004 11036 14105 11064
rect 13004 11008 13032 11036
rect 14093 11033 14105 11036
rect 14139 11033 14151 11067
rect 16132 11064 16160 11095
rect 17310 11092 17316 11144
rect 17368 11132 17374 11144
rect 17880 11132 17908 11163
rect 17368 11104 17908 11132
rect 17368 11092 17374 11104
rect 16132 11036 18644 11064
rect 14093 11027 14151 11033
rect 9732 10968 11100 10996
rect 9732 10956 9738 10968
rect 11146 10956 11152 11008
rect 11204 10956 11210 11008
rect 11514 10956 11520 11008
rect 11572 10956 11578 11008
rect 12986 10956 12992 11008
rect 13044 10956 13050 11008
rect 13170 10956 13176 11008
rect 13228 10956 13234 11008
rect 13998 10956 14004 11008
rect 14056 10996 14062 11008
rect 14553 10999 14611 11005
rect 14553 10996 14565 10999
rect 14056 10968 14565 10996
rect 14056 10956 14062 10968
rect 14553 10965 14565 10968
rect 14599 10996 14611 10999
rect 15654 10996 15660 11008
rect 14599 10968 15660 10996
rect 14599 10965 14611 10968
rect 14553 10959 14611 10965
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 15930 10956 15936 11008
rect 15988 10956 15994 11008
rect 17034 10956 17040 11008
rect 17092 10956 17098 11008
rect 17218 10956 17224 11008
rect 17276 10996 17282 11008
rect 17497 10999 17555 11005
rect 17497 10996 17509 10999
rect 17276 10968 17509 10996
rect 17276 10956 17282 10968
rect 17497 10965 17509 10968
rect 17543 10996 17555 10999
rect 17681 10999 17739 11005
rect 17681 10996 17693 10999
rect 17543 10968 17693 10996
rect 17543 10965 17555 10968
rect 17497 10959 17555 10965
rect 17681 10965 17693 10968
rect 17727 10965 17739 10999
rect 17681 10959 17739 10965
rect 18046 10956 18052 11008
rect 18104 10956 18110 11008
rect 18616 11005 18644 11036
rect 18690 11024 18696 11076
rect 18748 11064 18754 11076
rect 19168 11064 19196 11163
rect 19352 11132 19380 11163
rect 19426 11160 19432 11212
rect 19484 11160 19490 11212
rect 19628 11172 19840 11200
rect 19628 11132 19656 11172
rect 19352 11104 19656 11132
rect 19812 11132 19840 11172
rect 19886 11160 19892 11212
rect 19944 11160 19950 11212
rect 20070 11132 20076 11144
rect 19812 11104 20076 11132
rect 20070 11092 20076 11104
rect 20128 11132 20134 11144
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 20128 11104 20361 11132
rect 20128 11092 20134 11104
rect 20349 11101 20361 11104
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 20456 11064 20484 11240
rect 22373 11237 22385 11271
rect 22419 11268 22431 11271
rect 24121 11271 24179 11277
rect 24121 11268 24133 11271
rect 22419 11240 24133 11268
rect 22419 11237 22431 11240
rect 22373 11231 22431 11237
rect 24121 11237 24133 11240
rect 24167 11268 24179 11271
rect 25593 11271 25651 11277
rect 25593 11268 25605 11271
rect 24167 11240 25605 11268
rect 24167 11237 24179 11240
rect 24121 11231 24179 11237
rect 25593 11237 25605 11240
rect 25639 11237 25651 11271
rect 25593 11231 25651 11237
rect 27798 11228 27804 11280
rect 27856 11268 27862 11280
rect 29365 11271 29423 11277
rect 27856 11240 29132 11268
rect 27856 11228 27862 11240
rect 29104 11212 29132 11240
rect 29365 11237 29377 11271
rect 29411 11268 29423 11271
rect 29638 11268 29644 11280
rect 29411 11240 29644 11268
rect 29411 11237 29423 11240
rect 29365 11231 29423 11237
rect 29638 11228 29644 11240
rect 29696 11228 29702 11280
rect 31021 11271 31079 11277
rect 31021 11268 31033 11271
rect 30590 11240 31033 11268
rect 31021 11237 31033 11240
rect 31067 11237 31079 11271
rect 31021 11231 31079 11237
rect 32122 11228 32128 11280
rect 32180 11228 32186 11280
rect 33873 11271 33931 11277
rect 33873 11268 33885 11271
rect 33350 11240 33885 11268
rect 33873 11237 33885 11240
rect 33919 11237 33931 11271
rect 33873 11231 33931 11237
rect 22465 11203 22523 11209
rect 22465 11169 22477 11203
rect 22511 11200 22523 11203
rect 22511 11172 22692 11200
rect 22511 11169 22523 11172
rect 22465 11163 22523 11169
rect 22664 11144 22692 11172
rect 23014 11160 23020 11212
rect 23072 11200 23078 11212
rect 23109 11203 23167 11209
rect 23109 11200 23121 11203
rect 23072 11172 23121 11200
rect 23072 11160 23078 11172
rect 23109 11169 23121 11172
rect 23155 11200 23167 11203
rect 23290 11200 23296 11212
rect 23155 11172 23296 11200
rect 23155 11169 23167 11172
rect 23109 11163 23167 11169
rect 23290 11160 23296 11172
rect 23348 11160 23354 11212
rect 23658 11200 23664 11212
rect 23400 11172 23664 11200
rect 21913 11135 21971 11141
rect 21913 11101 21925 11135
rect 21959 11132 21971 11135
rect 22557 11135 22615 11141
rect 21959 11104 22048 11132
rect 21959 11101 21971 11104
rect 21913 11095 21971 11101
rect 22020 11073 22048 11104
rect 22557 11101 22569 11135
rect 22603 11101 22615 11135
rect 22557 11095 22615 11101
rect 18748 11036 20484 11064
rect 22005 11067 22063 11073
rect 18748 11024 18754 11036
rect 22005 11033 22017 11067
rect 22051 11033 22063 11067
rect 22572 11064 22600 11095
rect 22646 11092 22652 11144
rect 22704 11092 22710 11144
rect 23400 11132 23428 11172
rect 23658 11160 23664 11172
rect 23716 11200 23722 11212
rect 25685 11203 25743 11209
rect 23716 11172 24532 11200
rect 23716 11160 23722 11172
rect 24504 11144 24532 11172
rect 25685 11169 25697 11203
rect 25731 11200 25743 11203
rect 27249 11203 27307 11209
rect 25731 11172 26556 11200
rect 25731 11169 25743 11172
rect 25685 11163 25743 11169
rect 22756 11104 23428 11132
rect 22756 11064 22784 11104
rect 23474 11092 23480 11144
rect 23532 11092 23538 11144
rect 24486 11092 24492 11144
rect 24544 11092 24550 11144
rect 24854 11092 24860 11144
rect 24912 11092 24918 11144
rect 25501 11135 25559 11141
rect 25501 11101 25513 11135
rect 25547 11132 25559 11135
rect 26234 11132 26240 11144
rect 25547 11104 26240 11132
rect 25547 11101 25559 11104
rect 25501 11095 25559 11101
rect 26234 11092 26240 11104
rect 26292 11092 26298 11144
rect 26418 11092 26424 11144
rect 26476 11092 26482 11144
rect 22572 11036 22784 11064
rect 23201 11067 23259 11073
rect 22005 11027 22063 11033
rect 23201 11033 23213 11067
rect 23247 11064 23259 11067
rect 26528 11064 26556 11172
rect 27249 11169 27261 11203
rect 27295 11200 27307 11203
rect 28261 11203 28319 11209
rect 28261 11200 28273 11203
rect 27295 11172 28273 11200
rect 27295 11169 27307 11172
rect 27249 11163 27307 11169
rect 28261 11169 28273 11172
rect 28307 11200 28319 11203
rect 28534 11200 28540 11212
rect 28307 11172 28540 11200
rect 28307 11169 28319 11172
rect 28261 11163 28319 11169
rect 28534 11160 28540 11172
rect 28592 11160 28598 11212
rect 28629 11203 28687 11209
rect 28629 11169 28641 11203
rect 28675 11200 28687 11203
rect 28718 11200 28724 11212
rect 28675 11172 28724 11200
rect 28675 11169 28687 11172
rect 28629 11163 28687 11169
rect 28718 11160 28724 11172
rect 28776 11160 28782 11212
rect 28813 11203 28871 11209
rect 28813 11169 28825 11203
rect 28859 11200 28871 11203
rect 28902 11200 28908 11212
rect 28859 11172 28908 11200
rect 28859 11169 28871 11172
rect 28813 11163 28871 11169
rect 28902 11160 28908 11172
rect 28960 11160 28966 11212
rect 29086 11160 29092 11212
rect 29144 11160 29150 11212
rect 31113 11203 31171 11209
rect 31113 11169 31125 11203
rect 31159 11200 31171 11203
rect 31202 11200 31208 11212
rect 31159 11172 31208 11200
rect 31159 11169 31171 11172
rect 31113 11163 31171 11169
rect 26970 11092 26976 11144
rect 27028 11132 27034 11144
rect 27893 11135 27951 11141
rect 27893 11132 27905 11135
rect 27028 11104 27905 11132
rect 27028 11092 27034 11104
rect 27893 11101 27905 11104
rect 27939 11101 27951 11135
rect 28552 11132 28580 11160
rect 31128 11132 31156 11163
rect 31202 11160 31208 11172
rect 31260 11160 31266 11212
rect 33781 11203 33839 11209
rect 33781 11169 33793 11203
rect 33827 11200 33839 11203
rect 33980 11200 34008 11308
rect 33827 11172 34008 11200
rect 33827 11169 33839 11172
rect 33781 11163 33839 11169
rect 28552 11104 31156 11132
rect 27893 11095 27951 11101
rect 31662 11092 31668 11144
rect 31720 11132 31726 11144
rect 31849 11135 31907 11141
rect 31849 11132 31861 11135
rect 31720 11104 31861 11132
rect 31720 11092 31726 11104
rect 31849 11101 31861 11104
rect 31895 11101 31907 11135
rect 31849 11095 31907 11101
rect 32582 11092 32588 11144
rect 32640 11132 32646 11144
rect 33597 11135 33655 11141
rect 33597 11132 33609 11135
rect 32640 11104 33609 11132
rect 32640 11092 32646 11104
rect 33597 11101 33609 11104
rect 33643 11101 33655 11135
rect 33597 11095 33655 11101
rect 23247 11036 23980 11064
rect 26528 11036 27384 11064
rect 23247 11033 23259 11036
rect 23201 11027 23259 11033
rect 23952 11008 23980 11036
rect 27356 11008 27384 11036
rect 18601 10999 18659 11005
rect 18601 10965 18613 10999
rect 18647 10996 18659 10999
rect 19242 10996 19248 11008
rect 18647 10968 19248 10996
rect 18647 10965 18659 10968
rect 18601 10959 18659 10965
rect 19242 10956 19248 10968
rect 19300 10956 19306 11008
rect 20990 10956 20996 11008
rect 21048 10956 21054 11008
rect 21266 10956 21272 11008
rect 21324 10956 21330 11008
rect 23934 10956 23940 11008
rect 23992 10956 23998 11008
rect 24210 10956 24216 11008
rect 24268 10956 24274 11008
rect 27338 10956 27344 11008
rect 27396 10956 27402 11008
rect 2760 10906 34316 10928
rect 2760 10854 6550 10906
rect 6602 10854 6614 10906
rect 6666 10854 6678 10906
rect 6730 10854 6742 10906
rect 6794 10854 6806 10906
rect 6858 10854 14439 10906
rect 14491 10854 14503 10906
rect 14555 10854 14567 10906
rect 14619 10854 14631 10906
rect 14683 10854 14695 10906
rect 14747 10854 22328 10906
rect 22380 10854 22392 10906
rect 22444 10854 22456 10906
rect 22508 10854 22520 10906
rect 22572 10854 22584 10906
rect 22636 10854 30217 10906
rect 30269 10854 30281 10906
rect 30333 10854 30345 10906
rect 30397 10854 30409 10906
rect 30461 10854 30473 10906
rect 30525 10854 34316 10906
rect 2760 10832 34316 10854
rect 4543 10795 4601 10801
rect 4543 10761 4555 10795
rect 4589 10792 4601 10795
rect 6270 10792 6276 10804
rect 4589 10764 6276 10792
rect 4589 10761 4601 10764
rect 4543 10755 4601 10761
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 8849 10795 8907 10801
rect 8849 10792 8861 10795
rect 6748 10764 8861 10792
rect 6181 10727 6239 10733
rect 4724 10696 5764 10724
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4724 10656 4752 10696
rect 4212 10628 4752 10656
rect 4212 10616 4218 10628
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 5736 10665 5764 10696
rect 6181 10693 6193 10727
rect 6227 10724 6239 10727
rect 6638 10724 6644 10736
rect 6227 10696 6644 10724
rect 6227 10693 6239 10696
rect 6181 10687 6239 10693
rect 6638 10684 6644 10696
rect 6696 10684 6702 10736
rect 5721 10659 5779 10665
rect 5721 10625 5733 10659
rect 5767 10625 5779 10659
rect 5721 10619 5779 10625
rect 5074 10597 5080 10600
rect 4801 10591 4859 10597
rect 4801 10557 4813 10591
rect 4847 10557 4859 10591
rect 5069 10588 5080 10597
rect 4801 10551 4859 10557
rect 4908 10560 5080 10588
rect 3510 10480 3516 10532
rect 3568 10480 3574 10532
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 4816 10520 4844 10551
rect 4672 10492 4844 10520
rect 4672 10480 4678 10492
rect 3053 10455 3111 10461
rect 3053 10421 3065 10455
rect 3099 10452 3111 10455
rect 4154 10452 4160 10464
rect 3099 10424 4160 10452
rect 3099 10421 3111 10424
rect 3053 10415 3111 10421
rect 4154 10412 4160 10424
rect 4212 10412 4218 10464
rect 4430 10412 4436 10464
rect 4488 10452 4494 10464
rect 4908 10452 4936 10560
rect 5069 10551 5080 10560
rect 5074 10548 5080 10551
rect 5132 10548 5138 10600
rect 6748 10588 6776 10764
rect 8849 10761 8861 10764
rect 8895 10761 8907 10795
rect 8849 10755 8907 10761
rect 9769 10795 9827 10801
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 10318 10792 10324 10804
rect 9815 10764 10324 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 11330 10752 11336 10804
rect 11388 10752 11394 10804
rect 11688 10795 11746 10801
rect 11688 10761 11700 10795
rect 11734 10792 11746 10795
rect 13170 10792 13176 10804
rect 11734 10764 13176 10792
rect 11734 10761 11746 10764
rect 11688 10755 11746 10761
rect 13170 10752 13176 10764
rect 13228 10752 13234 10804
rect 16666 10752 16672 10804
rect 16724 10752 16730 10804
rect 16942 10752 16948 10804
rect 17000 10752 17006 10804
rect 18874 10752 18880 10804
rect 18932 10752 18938 10804
rect 23109 10795 23167 10801
rect 23109 10761 23121 10795
rect 23155 10792 23167 10795
rect 23474 10792 23480 10804
rect 23155 10764 23480 10792
rect 23155 10761 23167 10764
rect 23109 10755 23167 10761
rect 23474 10752 23480 10764
rect 23532 10752 23538 10804
rect 24949 10795 25007 10801
rect 24949 10761 24961 10795
rect 24995 10792 25007 10795
rect 25314 10792 25320 10804
rect 24995 10764 25320 10792
rect 24995 10761 25007 10764
rect 24949 10755 25007 10761
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 26053 10795 26111 10801
rect 26053 10761 26065 10795
rect 26099 10792 26111 10795
rect 26970 10792 26976 10804
rect 26099 10764 26976 10792
rect 26099 10761 26111 10764
rect 26053 10755 26111 10761
rect 26970 10752 26976 10764
rect 27028 10752 27034 10804
rect 28074 10752 28080 10804
rect 28132 10792 28138 10804
rect 28353 10795 28411 10801
rect 28353 10792 28365 10795
rect 28132 10764 28365 10792
rect 28132 10752 28138 10764
rect 28353 10761 28365 10764
rect 28399 10761 28411 10795
rect 28353 10755 28411 10761
rect 8110 10684 8116 10736
rect 8168 10724 8174 10736
rect 8168 10696 8616 10724
rect 8168 10684 8174 10696
rect 7374 10616 7380 10668
rect 7432 10656 7438 10668
rect 8021 10659 8079 10665
rect 8021 10656 8033 10659
rect 7432 10628 8033 10656
rect 7432 10616 7438 10628
rect 8021 10625 8033 10628
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 8386 10616 8392 10668
rect 8444 10616 8450 10668
rect 6670 10560 6776 10588
rect 8297 10591 8355 10597
rect 8297 10557 8309 10591
rect 8343 10588 8355 10591
rect 8404 10588 8432 10616
rect 8343 10560 8432 10588
rect 8481 10591 8539 10597
rect 8343 10557 8355 10560
rect 8297 10551 8355 10557
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8588 10588 8616 10696
rect 8956 10696 9812 10724
rect 8527 10560 8616 10588
rect 8665 10591 8723 10597
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8665 10557 8677 10591
rect 8711 10588 8723 10591
rect 8754 10588 8760 10600
rect 8711 10560 8760 10588
rect 8711 10557 8723 10560
rect 8665 10551 8723 10557
rect 8754 10548 8760 10560
rect 8812 10548 8818 10600
rect 8956 10597 8984 10696
rect 9674 10656 9680 10668
rect 9416 10628 9680 10656
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8864 10560 8953 10588
rect 8864 10532 8892 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 9416 10597 9444 10628
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 9217 10591 9275 10597
rect 9217 10588 9229 10591
rect 9180 10560 9229 10588
rect 9180 10548 9186 10560
rect 9217 10557 9229 10560
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9582 10548 9588 10600
rect 9640 10588 9646 10600
rect 9784 10588 9812 10696
rect 9858 10684 9864 10736
rect 9916 10724 9922 10736
rect 9953 10727 10011 10733
rect 9953 10724 9965 10727
rect 9916 10696 9965 10724
rect 9916 10684 9922 10696
rect 9953 10693 9965 10696
rect 9999 10693 10011 10727
rect 9953 10687 10011 10693
rect 14553 10727 14611 10733
rect 14553 10693 14565 10727
rect 14599 10693 14611 10727
rect 14553 10687 14611 10693
rect 11425 10659 11483 10665
rect 11425 10625 11437 10659
rect 11471 10656 11483 10659
rect 11790 10656 11796 10668
rect 11471 10628 11796 10656
rect 11471 10625 11483 10628
rect 11425 10619 11483 10625
rect 11790 10616 11796 10628
rect 11848 10656 11854 10668
rect 14274 10656 14280 10668
rect 11848 10628 14280 10656
rect 11848 10616 11854 10628
rect 14274 10616 14280 10628
rect 14332 10656 14338 10668
rect 14568 10656 14596 10687
rect 14918 10684 14924 10736
rect 14976 10724 14982 10736
rect 16684 10724 16712 10752
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 14976 10696 16344 10724
rect 16684 10696 17785 10724
rect 14976 10684 14982 10696
rect 16206 10656 16212 10668
rect 14332 10628 14596 10656
rect 15304 10628 16212 10656
rect 14332 10616 14338 10628
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9640 10548 9674 10588
rect 9784 10560 10057 10588
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 10781 10591 10839 10597
rect 10781 10557 10793 10591
rect 10827 10588 10839 10591
rect 10870 10588 10876 10600
rect 10827 10560 10876 10588
rect 10827 10557 10839 10560
rect 10781 10551 10839 10557
rect 10870 10548 10876 10560
rect 10928 10548 10934 10600
rect 10962 10548 10968 10600
rect 11020 10548 11026 10600
rect 11149 10591 11207 10597
rect 11149 10557 11161 10591
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 7745 10523 7803 10529
rect 7745 10489 7757 10523
rect 7791 10489 7803 10523
rect 7745 10483 7803 10489
rect 4488 10424 4936 10452
rect 4488 10412 4494 10424
rect 5166 10412 5172 10464
rect 5224 10412 5230 10464
rect 5813 10455 5871 10461
rect 5813 10421 5825 10455
rect 5859 10452 5871 10455
rect 6086 10452 6092 10464
rect 5859 10424 6092 10452
rect 5859 10421 5871 10424
rect 5813 10415 5871 10421
rect 6086 10412 6092 10424
rect 6144 10412 6150 10464
rect 6273 10455 6331 10461
rect 6273 10421 6285 10455
rect 6319 10452 6331 10455
rect 6454 10452 6460 10464
rect 6319 10424 6460 10452
rect 6319 10421 6331 10424
rect 6273 10415 6331 10421
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 7760 10452 7788 10483
rect 8202 10480 8208 10532
rect 8260 10520 8266 10532
rect 8389 10523 8447 10529
rect 8389 10520 8401 10523
rect 8260 10492 8401 10520
rect 8260 10480 8266 10492
rect 8389 10489 8401 10492
rect 8435 10489 8447 10523
rect 8389 10483 8447 10489
rect 8846 10480 8852 10532
rect 8904 10480 8910 10532
rect 9493 10523 9551 10529
rect 9493 10489 9505 10523
rect 9539 10489 9551 10523
rect 9493 10483 9551 10489
rect 8113 10455 8171 10461
rect 8113 10452 8125 10455
rect 7760 10424 8125 10452
rect 8113 10421 8125 10424
rect 8159 10421 8171 10455
rect 8113 10415 8171 10421
rect 8478 10412 8484 10464
rect 8536 10452 8542 10464
rect 9508 10452 9536 10483
rect 8536 10424 9536 10452
rect 9646 10452 9674 10548
rect 11057 10523 11115 10529
rect 11057 10489 11069 10523
rect 11103 10489 11115 10523
rect 11164 10520 11192 10551
rect 13446 10548 13452 10600
rect 13504 10548 13510 10600
rect 14182 10548 14188 10600
rect 14240 10588 14246 10600
rect 15304 10597 15332 10628
rect 16206 10616 16212 10628
rect 16264 10616 16270 10668
rect 16316 10656 16344 10696
rect 17773 10693 17785 10696
rect 17819 10724 17831 10727
rect 18417 10727 18475 10733
rect 18417 10724 18429 10727
rect 17819 10696 18429 10724
rect 17819 10693 17831 10696
rect 17773 10687 17831 10693
rect 18417 10693 18429 10696
rect 18463 10693 18475 10727
rect 18417 10687 18475 10693
rect 16482 10656 16488 10668
rect 16316 10628 16488 10656
rect 16482 10616 16488 10628
rect 16540 10656 16546 10668
rect 16540 10628 17816 10656
rect 16540 10616 16546 10628
rect 17788 10600 17816 10628
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14240 10560 15301 10588
rect 14240 10548 14246 10560
rect 15289 10557 15301 10560
rect 15335 10557 15347 10591
rect 15289 10551 15347 10557
rect 15746 10548 15752 10600
rect 15804 10548 15810 10600
rect 15930 10548 15936 10600
rect 15988 10548 15994 10600
rect 16298 10548 16304 10600
rect 16356 10548 16362 10600
rect 17037 10591 17095 10597
rect 17037 10557 17049 10591
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 11698 10520 11704 10532
rect 11164 10492 11704 10520
rect 11057 10483 11115 10489
rect 10321 10455 10379 10461
rect 10321 10452 10333 10455
rect 9646 10424 10333 10452
rect 8536 10412 8542 10424
rect 10321 10421 10333 10424
rect 10367 10421 10379 10455
rect 11072 10452 11100 10483
rect 11698 10480 11704 10492
rect 11756 10480 11762 10532
rect 12986 10520 12992 10532
rect 12926 10492 12992 10520
rect 12986 10480 12992 10492
rect 13044 10480 13050 10532
rect 13078 10480 13084 10532
rect 13136 10520 13142 10532
rect 13265 10523 13323 10529
rect 13265 10520 13277 10523
rect 13136 10492 13277 10520
rect 13136 10480 13142 10492
rect 13265 10489 13277 10492
rect 13311 10489 13323 10523
rect 13265 10483 13323 10489
rect 12526 10452 12532 10464
rect 11072 10424 12532 10452
rect 10321 10415 10379 10421
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 13173 10455 13231 10461
rect 13173 10421 13185 10455
rect 13219 10452 13231 10455
rect 13464 10452 13492 10548
rect 15948 10520 15976 10548
rect 17052 10520 17080 10551
rect 17402 10548 17408 10600
rect 17460 10548 17466 10600
rect 17770 10548 17776 10600
rect 17828 10548 17834 10600
rect 18432 10588 18460 10687
rect 18892 10656 18920 10752
rect 23014 10724 23020 10736
rect 22756 10696 23020 10724
rect 19613 10659 19671 10665
rect 18892 10628 19288 10656
rect 18966 10588 18972 10600
rect 18432 10560 18972 10588
rect 18966 10548 18972 10560
rect 19024 10588 19030 10600
rect 19150 10588 19156 10600
rect 19024 10560 19156 10588
rect 19024 10548 19030 10560
rect 19150 10548 19156 10560
rect 19208 10548 19214 10600
rect 19260 10597 19288 10628
rect 19613 10625 19625 10659
rect 19659 10656 19671 10659
rect 19702 10656 19708 10668
rect 19659 10628 19708 10656
rect 19659 10625 19671 10628
rect 19613 10619 19671 10625
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 22756 10656 22784 10696
rect 23014 10684 23020 10696
rect 23072 10684 23078 10736
rect 20548 10628 22784 10656
rect 19245 10591 19303 10597
rect 19245 10557 19257 10591
rect 19291 10557 19303 10591
rect 19245 10551 19303 10557
rect 20438 10548 20444 10600
rect 20496 10588 20502 10600
rect 20548 10597 20576 10628
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 23201 10659 23259 10665
rect 23201 10656 23213 10659
rect 22888 10628 23213 10656
rect 22888 10616 22894 10628
rect 23201 10625 23213 10628
rect 23247 10625 23259 10659
rect 23201 10619 23259 10625
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10656 23535 10659
rect 24210 10656 24216 10668
rect 23523 10628 24216 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 24210 10616 24216 10628
rect 24268 10616 24274 10668
rect 25332 10656 25360 10752
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 25332 10628 25605 10656
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 28810 10616 28816 10668
rect 28868 10656 28874 10668
rect 28905 10659 28963 10665
rect 28905 10656 28917 10659
rect 28868 10628 28917 10656
rect 28868 10616 28874 10628
rect 28905 10625 28917 10628
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 33781 10659 33839 10665
rect 33781 10625 33793 10659
rect 33827 10656 33839 10659
rect 34882 10656 34888 10668
rect 33827 10628 34888 10656
rect 33827 10625 33839 10628
rect 33781 10619 33839 10625
rect 34882 10616 34888 10628
rect 34940 10616 34946 10668
rect 20533 10591 20591 10597
rect 20533 10588 20545 10591
rect 20496 10560 20545 10588
rect 20496 10548 20502 10560
rect 20533 10557 20545 10560
rect 20579 10557 20591 10591
rect 20533 10551 20591 10557
rect 20901 10591 20959 10597
rect 20901 10557 20913 10591
rect 20947 10588 20959 10591
rect 20990 10588 20996 10600
rect 20947 10560 20996 10588
rect 20947 10557 20959 10560
rect 20901 10551 20959 10557
rect 20990 10548 20996 10560
rect 21048 10548 21054 10600
rect 21361 10591 21419 10597
rect 21361 10588 21373 10591
rect 21192 10560 21373 10588
rect 15764 10492 17080 10520
rect 17313 10523 17371 10529
rect 15764 10464 15792 10492
rect 17313 10489 17325 10523
rect 17359 10489 17371 10523
rect 17420 10520 17448 10548
rect 19705 10523 19763 10529
rect 17420 10492 19104 10520
rect 17313 10483 17371 10489
rect 13219 10424 13492 10452
rect 15381 10455 15439 10461
rect 13219 10421 13231 10424
rect 13173 10415 13231 10421
rect 15381 10421 15393 10455
rect 15427 10452 15439 10455
rect 15562 10452 15568 10464
rect 15427 10424 15568 10452
rect 15427 10421 15439 10424
rect 15381 10415 15439 10421
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 15746 10412 15752 10464
rect 15804 10412 15810 10464
rect 15838 10412 15844 10464
rect 15896 10412 15902 10464
rect 17328 10452 17356 10483
rect 17586 10452 17592 10464
rect 17328 10424 17592 10452
rect 17586 10412 17592 10424
rect 17644 10412 17650 10464
rect 19076 10452 19104 10492
rect 19705 10489 19717 10523
rect 19751 10520 19763 10523
rect 19886 10520 19892 10532
rect 19751 10492 19892 10520
rect 19751 10489 19763 10492
rect 19705 10483 19763 10489
rect 19720 10452 19748 10483
rect 19886 10480 19892 10492
rect 19944 10520 19950 10532
rect 19944 10492 21128 10520
rect 19944 10480 19950 10492
rect 19076 10424 19748 10452
rect 20622 10412 20628 10464
rect 20680 10412 20686 10464
rect 21100 10461 21128 10492
rect 21192 10464 21220 10560
rect 21361 10557 21373 10560
rect 21407 10557 21419 10591
rect 21361 10551 21419 10557
rect 22738 10548 22744 10600
rect 22796 10548 22802 10600
rect 27798 10548 27804 10600
rect 27856 10548 27862 10600
rect 28721 10591 28779 10597
rect 28721 10557 28733 10591
rect 28767 10588 28779 10591
rect 28994 10588 29000 10600
rect 28767 10560 29000 10588
rect 28767 10557 28779 10560
rect 28721 10551 28779 10557
rect 28994 10548 29000 10560
rect 29052 10548 29058 10600
rect 29362 10548 29368 10600
rect 29420 10588 29426 10600
rect 29733 10591 29791 10597
rect 29733 10588 29745 10591
rect 29420 10560 29745 10588
rect 29420 10548 29426 10560
rect 29733 10557 29745 10560
rect 29779 10557 29791 10591
rect 29733 10551 29791 10557
rect 29914 10548 29920 10600
rect 29972 10548 29978 10600
rect 30006 10548 30012 10600
rect 30064 10588 30070 10600
rect 30745 10591 30803 10597
rect 30745 10588 30757 10591
rect 30064 10560 30757 10588
rect 30064 10548 30070 10560
rect 30745 10557 30757 10560
rect 30791 10557 30803 10591
rect 30745 10551 30803 10557
rect 30837 10591 30895 10597
rect 30837 10557 30849 10591
rect 30883 10588 30895 10591
rect 30926 10588 30932 10600
rect 30883 10560 30932 10588
rect 30883 10557 30895 10560
rect 30837 10551 30895 10557
rect 21266 10480 21272 10532
rect 21324 10520 21330 10532
rect 21637 10523 21695 10529
rect 21637 10520 21649 10523
rect 21324 10492 21649 10520
rect 21324 10480 21330 10492
rect 21637 10489 21649 10492
rect 21683 10489 21695 10523
rect 21637 10483 21695 10489
rect 23934 10480 23940 10532
rect 23992 10480 23998 10532
rect 25958 10480 25964 10532
rect 26016 10520 26022 10532
rect 27525 10523 27583 10529
rect 26016 10492 26358 10520
rect 26016 10480 26022 10492
rect 27525 10489 27537 10523
rect 27571 10520 27583 10523
rect 29181 10523 29239 10529
rect 29181 10520 29193 10523
rect 27571 10492 29193 10520
rect 27571 10489 27583 10492
rect 27525 10483 27583 10489
rect 29181 10489 29193 10492
rect 29227 10489 29239 10523
rect 30852 10520 30880 10551
rect 30926 10548 30932 10560
rect 30984 10548 30990 10600
rect 32582 10548 32588 10600
rect 32640 10548 32646 10600
rect 29181 10483 29239 10489
rect 30668 10492 30880 10520
rect 30668 10464 30696 10492
rect 21085 10455 21143 10461
rect 21085 10421 21097 10455
rect 21131 10421 21143 10455
rect 21085 10415 21143 10421
rect 21174 10412 21180 10464
rect 21232 10412 21238 10464
rect 25038 10412 25044 10464
rect 25096 10412 25102 10464
rect 28813 10455 28871 10461
rect 28813 10421 28825 10455
rect 28859 10452 28871 10455
rect 28902 10452 28908 10464
rect 28859 10424 28908 10452
rect 28859 10421 28871 10424
rect 28813 10415 28871 10421
rect 28902 10412 28908 10424
rect 28960 10412 28966 10464
rect 30190 10412 30196 10464
rect 30248 10452 30254 10464
rect 30561 10455 30619 10461
rect 30561 10452 30573 10455
rect 30248 10424 30573 10452
rect 30248 10412 30254 10424
rect 30561 10421 30573 10424
rect 30607 10421 30619 10455
rect 30561 10415 30619 10421
rect 30650 10412 30656 10464
rect 30708 10412 30714 10464
rect 2760 10362 34316 10384
rect 2760 10310 7210 10362
rect 7262 10310 7274 10362
rect 7326 10310 7338 10362
rect 7390 10310 7402 10362
rect 7454 10310 7466 10362
rect 7518 10310 15099 10362
rect 15151 10310 15163 10362
rect 15215 10310 15227 10362
rect 15279 10310 15291 10362
rect 15343 10310 15355 10362
rect 15407 10310 22988 10362
rect 23040 10310 23052 10362
rect 23104 10310 23116 10362
rect 23168 10310 23180 10362
rect 23232 10310 23244 10362
rect 23296 10310 30877 10362
rect 30929 10310 30941 10362
rect 30993 10310 31005 10362
rect 31057 10310 31069 10362
rect 31121 10310 31133 10362
rect 31185 10310 34316 10362
rect 2760 10288 34316 10310
rect 3510 10208 3516 10260
rect 3568 10248 3574 10260
rect 3605 10251 3663 10257
rect 3605 10248 3617 10251
rect 3568 10220 3617 10248
rect 3568 10208 3574 10220
rect 3605 10217 3617 10220
rect 3651 10217 3663 10251
rect 5350 10248 5356 10260
rect 3605 10211 3663 10217
rect 4172 10220 5356 10248
rect 4172 10189 4200 10220
rect 5350 10208 5356 10220
rect 5408 10208 5414 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5592 10220 6040 10248
rect 5592 10208 5598 10220
rect 3421 10183 3479 10189
rect 3421 10149 3433 10183
rect 3467 10180 3479 10183
rect 4065 10183 4123 10189
rect 3467 10152 4016 10180
rect 3467 10149 3479 10152
rect 3421 10143 3479 10149
rect 3988 10124 4016 10152
rect 4065 10149 4077 10183
rect 4111 10149 4123 10183
rect 4065 10143 4123 10149
rect 4157 10183 4215 10189
rect 4157 10149 4169 10183
rect 4203 10149 4215 10183
rect 4614 10180 4620 10192
rect 4157 10143 4215 10149
rect 4448 10152 4620 10180
rect 3513 10115 3571 10121
rect 3513 10081 3525 10115
rect 3559 10081 3571 10115
rect 3513 10075 3571 10081
rect 3528 9976 3556 10075
rect 3970 10072 3976 10124
rect 4028 10072 4034 10124
rect 4080 10044 4108 10143
rect 4338 10072 4344 10124
rect 4396 10072 4402 10124
rect 4448 10121 4476 10152
rect 4614 10140 4620 10152
rect 4672 10140 4678 10192
rect 4706 10140 4712 10192
rect 4764 10140 4770 10192
rect 5166 10140 5172 10192
rect 5224 10140 5230 10192
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10081 4491 10115
rect 6012 10112 6040 10220
rect 6086 10208 6092 10260
rect 6144 10248 6150 10260
rect 6273 10251 6331 10257
rect 6273 10248 6285 10251
rect 6144 10220 6285 10248
rect 6144 10208 6150 10220
rect 6273 10217 6285 10220
rect 6319 10217 6331 10251
rect 6273 10211 6331 10217
rect 6362 10208 6368 10260
rect 6420 10248 6426 10260
rect 8202 10248 8208 10260
rect 6420 10220 8208 10248
rect 6420 10208 6426 10220
rect 8202 10208 8208 10220
rect 8260 10208 8266 10260
rect 8294 10208 8300 10260
rect 8352 10208 8358 10260
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 8444 10220 8708 10248
rect 8444 10208 8450 10220
rect 6546 10140 6552 10192
rect 6604 10180 6610 10192
rect 8478 10180 8484 10192
rect 6604 10152 8484 10180
rect 6604 10140 6610 10152
rect 8478 10140 8484 10152
rect 8536 10140 8542 10192
rect 8680 10180 8708 10220
rect 8754 10208 8760 10260
rect 8812 10248 8818 10260
rect 9309 10251 9367 10257
rect 9309 10248 9321 10251
rect 8812 10220 9321 10248
rect 8812 10208 8818 10220
rect 9309 10217 9321 10220
rect 9355 10248 9367 10251
rect 10870 10248 10876 10260
rect 9355 10220 10876 10248
rect 9355 10217 9367 10220
rect 9309 10211 9367 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12526 10208 12532 10260
rect 12584 10248 12590 10260
rect 13538 10248 13544 10260
rect 12584 10220 13544 10248
rect 12584 10208 12590 10220
rect 13538 10208 13544 10220
rect 13596 10248 13602 10260
rect 14001 10251 14059 10257
rect 14001 10248 14013 10251
rect 13596 10220 14013 10248
rect 13596 10208 13602 10220
rect 14001 10217 14013 10220
rect 14047 10217 14059 10251
rect 14001 10211 14059 10217
rect 16025 10251 16083 10257
rect 16025 10217 16037 10251
rect 16071 10248 16083 10251
rect 16298 10248 16304 10260
rect 16071 10220 16304 10248
rect 16071 10217 16083 10220
rect 16025 10211 16083 10217
rect 16298 10208 16304 10220
rect 16356 10208 16362 10260
rect 17034 10208 17040 10260
rect 17092 10208 17098 10260
rect 17313 10251 17371 10257
rect 17313 10217 17325 10251
rect 17359 10248 17371 10251
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17359 10220 17693 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 17681 10211 17739 10217
rect 18046 10208 18052 10260
rect 18104 10208 18110 10260
rect 18141 10251 18199 10257
rect 18141 10217 18153 10251
rect 18187 10248 18199 10251
rect 18187 10220 18644 10248
rect 18187 10217 18199 10220
rect 18141 10211 18199 10217
rect 8941 10183 8999 10189
rect 8941 10180 8953 10183
rect 8680 10152 8953 10180
rect 8941 10149 8953 10152
rect 8987 10149 8999 10183
rect 8941 10143 8999 10149
rect 7193 10115 7251 10121
rect 7193 10112 7205 10115
rect 6012 10084 7205 10112
rect 4433 10075 4491 10081
rect 7193 10081 7205 10084
rect 7239 10112 7251 10115
rect 8662 10112 8668 10124
rect 7239 10084 8668 10112
rect 7239 10081 7251 10084
rect 7193 10075 7251 10081
rect 8662 10072 8668 10084
rect 8720 10072 8726 10124
rect 8956 10112 8984 10143
rect 9122 10140 9128 10192
rect 9180 10180 9186 10192
rect 9861 10183 9919 10189
rect 9861 10180 9873 10183
rect 9180 10152 9873 10180
rect 9180 10140 9186 10152
rect 9861 10149 9873 10152
rect 9907 10149 9919 10183
rect 9861 10143 9919 10149
rect 11514 10140 11520 10192
rect 11572 10140 11578 10192
rect 13262 10180 13268 10192
rect 12742 10152 13268 10180
rect 13262 10140 13268 10152
rect 13320 10140 13326 10192
rect 14553 10183 14611 10189
rect 14553 10149 14565 10183
rect 14599 10180 14611 10183
rect 14826 10180 14832 10192
rect 14599 10152 14832 10180
rect 14599 10149 14611 10152
rect 14553 10143 14611 10149
rect 14826 10140 14832 10152
rect 14884 10140 14890 10192
rect 15562 10140 15568 10192
rect 15620 10140 15626 10192
rect 16945 10183 17003 10189
rect 16945 10149 16957 10183
rect 16991 10180 17003 10183
rect 17218 10180 17224 10192
rect 16991 10152 17224 10180
rect 16991 10149 17003 10152
rect 16945 10143 17003 10149
rect 17218 10140 17224 10152
rect 17276 10180 17282 10192
rect 18064 10180 18092 10208
rect 18616 10189 18644 10220
rect 20070 10208 20076 10260
rect 20128 10208 20134 10260
rect 20622 10208 20628 10260
rect 20680 10208 20686 10260
rect 22738 10208 22744 10260
rect 22796 10248 22802 10260
rect 23109 10251 23167 10257
rect 23109 10248 23121 10251
rect 22796 10220 23121 10248
rect 22796 10208 22802 10220
rect 23109 10217 23121 10220
rect 23155 10217 23167 10251
rect 23109 10211 23167 10217
rect 23937 10251 23995 10257
rect 23937 10217 23949 10251
rect 23983 10248 23995 10251
rect 25038 10248 25044 10260
rect 23983 10220 25044 10248
rect 23983 10217 23995 10220
rect 23937 10211 23995 10217
rect 25038 10208 25044 10220
rect 25096 10208 25102 10260
rect 25958 10208 25964 10260
rect 26016 10208 26022 10260
rect 26513 10251 26571 10257
rect 26513 10217 26525 10251
rect 26559 10248 26571 10251
rect 27338 10248 27344 10260
rect 26559 10220 27344 10248
rect 26559 10217 26571 10220
rect 26513 10211 26571 10217
rect 27338 10208 27344 10220
rect 27396 10208 27402 10260
rect 29086 10208 29092 10260
rect 29144 10248 29150 10260
rect 29730 10248 29736 10260
rect 29144 10220 29736 10248
rect 29144 10208 29150 10220
rect 29730 10208 29736 10220
rect 29788 10248 29794 10260
rect 31202 10248 31208 10260
rect 29788 10220 31208 10248
rect 29788 10208 29794 10220
rect 17276 10152 18092 10180
rect 18601 10183 18659 10189
rect 17276 10140 17282 10152
rect 18601 10149 18613 10183
rect 18647 10149 18659 10183
rect 18601 10143 18659 10149
rect 19334 10140 19340 10192
rect 19392 10140 19398 10192
rect 20640 10180 20668 10208
rect 20640 10152 21206 10180
rect 26418 10140 26424 10192
rect 26476 10140 26482 10192
rect 30006 10180 30012 10192
rect 29670 10152 30012 10180
rect 30006 10140 30012 10152
rect 30064 10140 30070 10192
rect 30101 10183 30159 10189
rect 30101 10149 30113 10183
rect 30147 10180 30159 10183
rect 30190 10180 30196 10192
rect 30147 10152 30196 10180
rect 30147 10149 30159 10152
rect 30101 10143 30159 10149
rect 30190 10140 30196 10152
rect 30248 10140 30254 10192
rect 9306 10112 9312 10124
rect 8956 10084 9312 10112
rect 9306 10072 9312 10084
rect 9364 10112 9370 10124
rect 9582 10112 9588 10124
rect 9364 10084 9588 10112
rect 9364 10072 9370 10084
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 10594 10072 10600 10124
rect 10652 10112 10658 10124
rect 11241 10115 11299 10121
rect 11241 10112 11253 10115
rect 10652 10084 11253 10112
rect 10652 10072 10658 10084
rect 11241 10081 11253 10084
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 14274 10072 14280 10124
rect 14332 10072 14338 10124
rect 16577 10115 16635 10121
rect 16577 10081 16589 10115
rect 16623 10112 16635 10115
rect 17773 10115 17831 10121
rect 17773 10112 17785 10115
rect 16623 10084 16988 10112
rect 16623 10081 16635 10084
rect 16577 10075 16635 10081
rect 16960 10056 16988 10084
rect 17420 10084 17785 10112
rect 4246 10044 4252 10056
rect 4080 10016 4252 10044
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10044 6239 10047
rect 6825 10047 6883 10053
rect 6825 10044 6837 10047
rect 6227 10016 6837 10044
rect 6227 10013 6239 10016
rect 6181 10007 6239 10013
rect 6825 10013 6837 10016
rect 6871 10013 6883 10047
rect 6825 10007 6883 10013
rect 8202 10004 8208 10056
rect 8260 10044 8266 10056
rect 8846 10044 8852 10056
rect 8260 10016 8852 10044
rect 8260 10004 8266 10016
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 11146 10004 11152 10056
rect 11204 10044 11210 10056
rect 12526 10044 12532 10056
rect 11204 10016 12532 10044
rect 11204 10004 11210 10016
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10044 13047 10047
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 13035 10016 13369 10044
rect 13035 10013 13047 10016
rect 12989 10007 13047 10013
rect 13357 10013 13369 10016
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 15746 10004 15752 10056
rect 15804 10044 15810 10056
rect 16301 10047 16359 10053
rect 16301 10044 16313 10047
rect 15804 10016 16313 10044
rect 15804 10004 15810 10016
rect 16301 10013 16313 10016
rect 16347 10013 16359 10047
rect 16301 10007 16359 10013
rect 16669 10047 16727 10053
rect 16669 10013 16681 10047
rect 16715 10044 16727 10047
rect 16850 10044 16856 10056
rect 16715 10016 16856 10044
rect 16715 10013 16727 10016
rect 16669 10007 16727 10013
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 16942 10004 16948 10056
rect 17000 10004 17006 10056
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 17154 10047 17212 10053
rect 17154 10044 17166 10047
rect 17092 10016 17166 10044
rect 17092 10004 17098 10016
rect 17154 10013 17166 10016
rect 17200 10013 17212 10047
rect 17154 10007 17212 10013
rect 17420 9988 17448 10084
rect 17773 10081 17785 10084
rect 17819 10081 17831 10115
rect 17773 10075 17831 10081
rect 18322 10072 18328 10124
rect 18380 10072 18386 10124
rect 22094 10072 22100 10124
rect 22152 10112 22158 10124
rect 22738 10112 22744 10124
rect 22152 10084 22744 10112
rect 22152 10072 22158 10084
rect 22738 10072 22744 10084
rect 22796 10072 22802 10124
rect 23201 10115 23259 10121
rect 23201 10081 23213 10115
rect 23247 10112 23259 10115
rect 23247 10084 23428 10112
rect 23247 10081 23259 10084
rect 23201 10075 23259 10081
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 17678 10044 17684 10056
rect 17635 10016 17684 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 20441 10047 20499 10053
rect 18248 10016 19748 10044
rect 4430 9976 4436 9988
rect 3528 9948 4436 9976
rect 4430 9936 4436 9948
rect 4488 9936 4494 9988
rect 7653 9979 7711 9985
rect 7653 9945 7665 9979
rect 7699 9976 7711 9979
rect 7742 9976 7748 9988
rect 7699 9948 7748 9976
rect 7699 9945 7711 9948
rect 7653 9939 7711 9945
rect 7742 9936 7748 9948
rect 7800 9976 7806 9988
rect 7800 9948 9628 9976
rect 7800 9936 7806 9948
rect 9600 9920 9628 9948
rect 17402 9936 17408 9988
rect 17460 9936 17466 9988
rect 3789 9911 3847 9917
rect 3789 9877 3801 9911
rect 3835 9908 3847 9911
rect 5350 9908 5356 9920
rect 3835 9880 5356 9908
rect 3835 9877 3847 9880
rect 3789 9871 3847 9877
rect 5350 9868 5356 9880
rect 5408 9868 5414 9920
rect 8570 9868 8576 9920
rect 8628 9868 8634 9920
rect 9582 9868 9588 9920
rect 9640 9868 9646 9920
rect 10870 9868 10876 9920
rect 10928 9908 10934 9920
rect 11149 9911 11207 9917
rect 11149 9908 11161 9911
rect 10928 9880 11161 9908
rect 10928 9868 10934 9880
rect 11149 9877 11161 9880
rect 11195 9908 11207 9911
rect 18248 9908 18276 10016
rect 19720 9988 19748 10016
rect 20441 10013 20453 10047
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 19702 9936 19708 9988
rect 19760 9936 19766 9988
rect 11195 9880 18276 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 18322 9868 18328 9920
rect 18380 9908 18386 9920
rect 20456 9908 20484 10007
rect 20714 10004 20720 10056
rect 20772 10004 20778 10056
rect 22189 10047 22247 10053
rect 22189 10013 22201 10047
rect 22235 10044 22247 10047
rect 22281 10047 22339 10053
rect 22281 10044 22293 10047
rect 22235 10016 22293 10044
rect 22235 10013 22247 10016
rect 22189 10007 22247 10013
rect 22281 10013 22293 10016
rect 22327 10013 22339 10047
rect 22281 10007 22339 10013
rect 23400 9988 23428 10084
rect 23934 10072 23940 10124
rect 23992 10112 23998 10124
rect 24949 10115 25007 10121
rect 24949 10112 24961 10115
rect 23992 10084 24961 10112
rect 23992 10072 23998 10084
rect 24949 10081 24961 10084
rect 24995 10081 25007 10115
rect 24949 10075 25007 10081
rect 26053 10115 26111 10121
rect 26053 10081 26065 10115
rect 26099 10112 26111 10115
rect 26436 10112 26464 10140
rect 26970 10112 26976 10124
rect 26099 10084 26976 10112
rect 26099 10081 26111 10084
rect 26053 10075 26111 10081
rect 26970 10072 26976 10084
rect 27028 10072 27034 10124
rect 27430 10072 27436 10124
rect 27488 10072 27494 10124
rect 27525 10115 27583 10121
rect 27525 10081 27537 10115
rect 27571 10112 27583 10115
rect 28810 10112 28816 10124
rect 27571 10084 28816 10112
rect 27571 10081 27583 10084
rect 27525 10075 27583 10081
rect 28810 10072 28816 10084
rect 28868 10072 28874 10124
rect 30392 10121 30420 10220
rect 31202 10208 31208 10220
rect 31260 10248 31266 10260
rect 31662 10248 31668 10260
rect 31260 10220 31668 10248
rect 31260 10208 31266 10220
rect 31662 10208 31668 10220
rect 31720 10248 31726 10260
rect 31757 10251 31815 10257
rect 31757 10248 31769 10251
rect 31720 10220 31769 10248
rect 31720 10208 31726 10220
rect 31757 10217 31769 10220
rect 31803 10217 31815 10251
rect 31757 10211 31815 10217
rect 30377 10115 30435 10121
rect 30377 10081 30389 10115
rect 30423 10081 30435 10115
rect 30377 10075 30435 10081
rect 30469 10115 30527 10121
rect 30469 10081 30481 10115
rect 30515 10112 30527 10115
rect 31386 10112 31392 10124
rect 30515 10084 31392 10112
rect 30515 10081 30527 10084
rect 30469 10075 30527 10081
rect 31386 10072 31392 10084
rect 31444 10072 31450 10124
rect 33965 10115 34023 10121
rect 33965 10081 33977 10115
rect 34011 10081 34023 10115
rect 33965 10075 34023 10081
rect 23658 10004 23664 10056
rect 23716 10004 23722 10056
rect 23750 10004 23756 10056
rect 23808 10044 23814 10056
rect 23845 10047 23903 10053
rect 23845 10044 23857 10047
rect 23808 10016 23857 10044
rect 23808 10004 23814 10016
rect 23845 10013 23857 10016
rect 23891 10044 23903 10047
rect 24397 10047 24455 10053
rect 24397 10044 24409 10047
rect 23891 10016 24409 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24397 10013 24409 10016
rect 24443 10013 24455 10047
rect 24397 10007 24455 10013
rect 25682 10004 25688 10056
rect 25740 10004 25746 10056
rect 26234 10004 26240 10056
rect 26292 10004 26298 10056
rect 26418 10004 26424 10056
rect 26476 10004 26482 10056
rect 26510 10004 26516 10056
rect 26568 10044 26574 10056
rect 27617 10047 27675 10053
rect 27617 10044 27629 10047
rect 26568 10016 27629 10044
rect 26568 10004 26574 10016
rect 27617 10013 27629 10016
rect 27663 10013 27675 10047
rect 29362 10044 29368 10056
rect 27617 10007 27675 10013
rect 28276 10016 29368 10044
rect 21818 9936 21824 9988
rect 21876 9976 21882 9988
rect 22094 9976 22100 9988
rect 21876 9948 22100 9976
rect 21876 9936 21882 9948
rect 22094 9936 22100 9948
rect 22152 9936 22158 9988
rect 23382 9936 23388 9988
rect 23440 9936 23446 9988
rect 24305 9979 24363 9985
rect 24305 9945 24317 9979
rect 24351 9976 24363 9979
rect 24854 9976 24860 9988
rect 24351 9948 24860 9976
rect 24351 9945 24363 9948
rect 24305 9939 24363 9945
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 26528 9976 26556 10004
rect 24964 9948 26556 9976
rect 26881 9979 26939 9985
rect 21174 9908 21180 9920
rect 18380 9880 21180 9908
rect 18380 9868 18386 9880
rect 21174 9868 21180 9880
rect 21232 9868 21238 9920
rect 22646 9868 22652 9920
rect 22704 9908 22710 9920
rect 22922 9908 22928 9920
rect 22704 9880 22928 9908
rect 22704 9868 22710 9880
rect 22922 9868 22928 9880
rect 22980 9868 22986 9920
rect 23290 9868 23296 9920
rect 23348 9908 23354 9920
rect 24964 9908 24992 9948
rect 26881 9945 26893 9979
rect 26927 9976 26939 9979
rect 28276 9976 28304 10016
rect 29362 10004 29368 10016
rect 29420 10004 29426 10056
rect 33980 10044 34008 10075
rect 34422 10044 34428 10056
rect 33980 10016 34428 10044
rect 34422 10004 34428 10016
rect 34480 10004 34486 10056
rect 26927 9948 28304 9976
rect 26927 9945 26939 9948
rect 26881 9939 26939 9945
rect 23348 9880 24992 9908
rect 23348 9868 23354 9880
rect 25130 9868 25136 9920
rect 25188 9868 25194 9920
rect 27065 9911 27123 9917
rect 27065 9877 27077 9911
rect 27111 9908 27123 9911
rect 27154 9908 27160 9920
rect 27111 9880 27160 9908
rect 27111 9877 27123 9880
rect 27065 9871 27123 9877
rect 27154 9868 27160 9880
rect 27212 9868 27218 9920
rect 28629 9911 28687 9917
rect 28629 9877 28641 9911
rect 28675 9908 28687 9911
rect 29086 9908 29092 9920
rect 28675 9880 29092 9908
rect 28675 9877 28687 9880
rect 28629 9871 28687 9877
rect 29086 9868 29092 9880
rect 29144 9868 29150 9920
rect 33778 9868 33784 9920
rect 33836 9868 33842 9920
rect 2760 9818 34316 9840
rect 2760 9766 6550 9818
rect 6602 9766 6614 9818
rect 6666 9766 6678 9818
rect 6730 9766 6742 9818
rect 6794 9766 6806 9818
rect 6858 9766 14439 9818
rect 14491 9766 14503 9818
rect 14555 9766 14567 9818
rect 14619 9766 14631 9818
rect 14683 9766 14695 9818
rect 14747 9766 22328 9818
rect 22380 9766 22392 9818
rect 22444 9766 22456 9818
rect 22508 9766 22520 9818
rect 22572 9766 22584 9818
rect 22636 9766 30217 9818
rect 30269 9766 30281 9818
rect 30333 9766 30345 9818
rect 30397 9766 30409 9818
rect 30461 9766 30473 9818
rect 30525 9766 34316 9818
rect 2760 9744 34316 9766
rect 3970 9664 3976 9716
rect 4028 9704 4034 9716
rect 4028 9676 6040 9704
rect 4028 9664 4034 9676
rect 4706 9596 4712 9648
rect 4764 9596 4770 9648
rect 5445 9639 5503 9645
rect 5445 9605 5457 9639
rect 5491 9605 5503 9639
rect 5445 9599 5503 9605
rect 6012 9636 6040 9676
rect 11698 9664 11704 9716
rect 11756 9664 11762 9716
rect 13262 9664 13268 9716
rect 13320 9664 13326 9716
rect 14826 9664 14832 9716
rect 14884 9664 14890 9716
rect 15746 9664 15752 9716
rect 15804 9704 15810 9716
rect 16853 9707 16911 9713
rect 16853 9704 16865 9707
rect 15804 9676 16865 9704
rect 15804 9664 15810 9676
rect 16853 9673 16865 9676
rect 16899 9673 16911 9707
rect 16853 9667 16911 9673
rect 17034 9664 17040 9716
rect 17092 9664 17098 9716
rect 19334 9664 19340 9716
rect 19392 9664 19398 9716
rect 22480 9676 22692 9704
rect 7101 9639 7159 9645
rect 7101 9636 7113 9639
rect 6012 9608 6224 9636
rect 1302 9528 1308 9580
rect 1360 9568 1366 9580
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 1360 9540 3249 9568
rect 1360 9528 1366 9540
rect 3237 9537 3249 9540
rect 3283 9537 3295 9571
rect 3237 9531 3295 9537
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 4724 9568 4752 9596
rect 4663 9540 4752 9568
rect 5261 9571 5319 9577
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 5261 9537 5273 9571
rect 5307 9568 5319 9571
rect 5460 9568 5488 9599
rect 6012 9577 6040 9608
rect 6196 9580 6224 9608
rect 7024 9608 7113 9636
rect 5307 9540 5488 9568
rect 5997 9571 6055 9577
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6086 9528 6092 9580
rect 6144 9528 6150 9580
rect 6178 9528 6184 9580
rect 6236 9528 6242 9580
rect 7024 9577 7052 9608
rect 7101 9605 7113 9608
rect 7147 9605 7159 9639
rect 8570 9636 8576 9648
rect 7101 9599 7159 9605
rect 7392 9608 8576 9636
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 4154 9460 4160 9512
rect 4212 9500 4218 9512
rect 4249 9503 4307 9509
rect 4249 9500 4261 9503
rect 4212 9472 4261 9500
rect 4212 9460 4218 9472
rect 4249 9469 4261 9472
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5644 9432 5672 9463
rect 5718 9460 5724 9512
rect 5776 9460 5782 9512
rect 7392 9500 7420 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 14645 9639 14703 9645
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 15378 9636 15384 9648
rect 14691 9608 15384 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 8386 9568 8392 9580
rect 7708 9540 8392 9568
rect 7708 9528 7714 9540
rect 8386 9528 8392 9540
rect 8444 9568 8450 9580
rect 8849 9571 8907 9577
rect 8849 9568 8861 9571
rect 8444 9540 8861 9568
rect 8444 9528 8450 9540
rect 8849 9537 8861 9540
rect 8895 9537 8907 9571
rect 8849 9531 8907 9537
rect 6012 9472 7420 9500
rect 7469 9503 7527 9509
rect 6012 9432 6040 9472
rect 7469 9469 7481 9503
rect 7515 9500 7527 9503
rect 7558 9500 7564 9512
rect 7515 9472 7564 9500
rect 7515 9469 7527 9472
rect 7469 9463 7527 9469
rect 7558 9460 7564 9472
rect 7616 9460 7622 9512
rect 8018 9460 8024 9512
rect 8076 9500 8082 9512
rect 8481 9503 8539 9509
rect 8481 9500 8493 9503
rect 8076 9472 8493 9500
rect 8076 9460 8082 9472
rect 8481 9469 8493 9472
rect 8527 9469 8539 9503
rect 8864 9500 8892 9531
rect 12066 9528 12072 9580
rect 12124 9568 12130 9580
rect 14200 9568 14228 9596
rect 12124 9540 14228 9568
rect 12124 9528 12130 9540
rect 13372 9509 13400 9540
rect 13357 9503 13415 9509
rect 8864 9472 12434 9500
rect 8481 9463 8539 9469
rect 10686 9432 10692 9444
rect 5644 9404 6040 9432
rect 6104 9404 10692 9432
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 6104 9364 6132 9404
rect 10686 9392 10692 9404
rect 10744 9392 10750 9444
rect 12406 9432 12434 9472
rect 13357 9469 13369 9503
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9500 13875 9503
rect 13906 9500 13912 9512
rect 13863 9472 13912 9500
rect 13863 9469 13875 9472
rect 13817 9463 13875 9469
rect 13832 9432 13860 9463
rect 13906 9460 13912 9472
rect 13964 9460 13970 9512
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9500 14243 9503
rect 14660 9500 14688 9599
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 17678 9636 17684 9648
rect 15488 9608 17684 9636
rect 15488 9577 15516 9608
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 18785 9639 18843 9645
rect 18785 9605 18797 9639
rect 18831 9636 18843 9639
rect 19352 9636 19380 9664
rect 20806 9636 20812 9648
rect 18831 9608 19380 9636
rect 20088 9608 20812 9636
rect 18831 9605 18843 9608
rect 18785 9599 18843 9605
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9537 15531 9571
rect 15473 9531 15531 9537
rect 15838 9528 15844 9580
rect 15896 9528 15902 9580
rect 16574 9528 16580 9580
rect 16632 9528 16638 9580
rect 20088 9568 20116 9608
rect 20806 9596 20812 9608
rect 20864 9596 20870 9648
rect 22480 9636 22508 9676
rect 21468 9608 22508 9636
rect 22557 9639 22615 9645
rect 16684 9540 20116 9568
rect 20165 9571 20223 9577
rect 14231 9472 14688 9500
rect 15289 9503 15347 9509
rect 14231 9469 14243 9472
rect 14185 9463 14243 9469
rect 15289 9469 15301 9503
rect 15335 9500 15347 9503
rect 15856 9500 15884 9528
rect 15335 9472 15884 9500
rect 15335 9469 15347 9472
rect 15289 9463 15347 9469
rect 16684 9432 16712 9540
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 20530 9568 20536 9580
rect 20211 9540 20536 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 21468 9577 21496 9608
rect 22557 9605 22569 9639
rect 22603 9605 22615 9639
rect 22557 9599 22615 9605
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9568 22523 9571
rect 22572 9568 22600 9599
rect 22511 9540 22600 9568
rect 22664 9568 22692 9676
rect 25130 9664 25136 9716
rect 25188 9664 25194 9716
rect 28718 9704 28724 9716
rect 26252 9676 28724 9704
rect 22830 9568 22836 9580
rect 22664 9540 22836 9568
rect 22511 9537 22523 9540
rect 22465 9531 22523 9537
rect 22830 9528 22836 9540
rect 22888 9568 22894 9580
rect 23106 9568 23112 9580
rect 22888 9540 23112 9568
rect 22888 9528 22894 9540
rect 23106 9528 23112 9540
rect 23164 9528 23170 9580
rect 24121 9571 24179 9577
rect 24121 9537 24133 9571
rect 24167 9568 24179 9571
rect 25148 9568 25176 9664
rect 26252 9648 26280 9676
rect 28718 9664 28724 9676
rect 28776 9704 28782 9716
rect 28994 9704 29000 9716
rect 28776 9676 29000 9704
rect 28776 9664 28782 9676
rect 28994 9664 29000 9676
rect 29052 9664 29058 9716
rect 29549 9707 29607 9713
rect 29549 9673 29561 9707
rect 29595 9704 29607 9707
rect 29914 9704 29920 9716
rect 29595 9676 29920 9704
rect 29595 9673 29607 9676
rect 29549 9667 29607 9673
rect 29914 9664 29920 9676
rect 29972 9664 29978 9716
rect 31386 9664 31392 9716
rect 31444 9664 31450 9716
rect 25222 9596 25228 9648
rect 25280 9636 25286 9648
rect 25498 9636 25504 9648
rect 25280 9608 25504 9636
rect 25280 9596 25286 9608
rect 25498 9596 25504 9608
rect 25556 9636 25562 9648
rect 26053 9639 26111 9645
rect 26053 9636 26065 9639
rect 25556 9608 26065 9636
rect 25556 9596 25562 9608
rect 26053 9605 26065 9608
rect 26099 9605 26111 9639
rect 26053 9599 26111 9605
rect 26234 9596 26240 9648
rect 26292 9596 26298 9648
rect 33962 9636 33968 9648
rect 28644 9608 33968 9636
rect 24167 9540 25176 9568
rect 25593 9571 25651 9577
rect 24167 9537 24179 9540
rect 24121 9531 24179 9537
rect 25593 9537 25605 9571
rect 25639 9568 25651 9571
rect 26605 9571 26663 9577
rect 26605 9568 26617 9571
rect 25639 9540 26617 9568
rect 25639 9537 25651 9540
rect 25593 9531 25651 9537
rect 26605 9537 26617 9540
rect 26651 9537 26663 9571
rect 26605 9531 26663 9537
rect 26973 9571 27031 9577
rect 26973 9537 26985 9571
rect 27019 9568 27031 9571
rect 27798 9568 27804 9580
rect 27019 9540 27804 9568
rect 27019 9537 27031 9540
rect 26973 9531 27031 9537
rect 27798 9528 27804 9540
rect 27856 9528 27862 9580
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9500 17279 9503
rect 17402 9500 17408 9512
rect 17267 9472 17408 9500
rect 17267 9469 17279 9472
rect 17221 9463 17279 9469
rect 17402 9460 17408 9472
rect 17460 9460 17466 9512
rect 17497 9503 17555 9509
rect 17497 9469 17509 9503
rect 17543 9500 17555 9503
rect 17586 9500 17592 9512
rect 17543 9472 17592 9500
rect 17543 9469 17555 9472
rect 17497 9463 17555 9469
rect 17586 9460 17592 9472
rect 17644 9460 17650 9512
rect 18693 9503 18751 9509
rect 18693 9469 18705 9503
rect 18739 9469 18751 9503
rect 18693 9463 18751 9469
rect 12406 9404 13860 9432
rect 14476 9404 16712 9432
rect 3200 9336 6132 9364
rect 3200 9324 3206 9336
rect 6362 9324 6368 9376
rect 6420 9324 6426 9376
rect 7561 9367 7619 9373
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 7929 9367 7987 9373
rect 7929 9364 7941 9367
rect 7607 9336 7941 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 7929 9333 7941 9336
rect 7975 9333 7987 9367
rect 7929 9327 7987 9333
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10778 9364 10784 9376
rect 10008 9336 10784 9364
rect 10008 9324 10014 9336
rect 10778 9324 10784 9336
rect 10836 9324 10842 9376
rect 13078 9324 13084 9376
rect 13136 9324 13142 9376
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 14476 9364 14504 9404
rect 16758 9392 16764 9444
rect 16816 9432 16822 9444
rect 18049 9435 18107 9441
rect 18049 9432 18061 9435
rect 16816 9404 18061 9432
rect 16816 9392 16822 9404
rect 18049 9401 18061 9404
rect 18095 9401 18107 9435
rect 18049 9395 18107 9401
rect 18138 9392 18144 9444
rect 18196 9432 18202 9444
rect 18233 9435 18291 9441
rect 18233 9432 18245 9435
rect 18196 9404 18245 9432
rect 18196 9392 18202 9404
rect 18233 9401 18245 9404
rect 18279 9432 18291 9435
rect 18598 9432 18604 9444
rect 18279 9404 18604 9432
rect 18279 9401 18291 9404
rect 18233 9395 18291 9401
rect 18598 9392 18604 9404
rect 18656 9392 18662 9444
rect 18708 9432 18736 9463
rect 19242 9460 19248 9512
rect 19300 9500 19306 9512
rect 19705 9503 19763 9509
rect 19705 9500 19717 9503
rect 19300 9472 19717 9500
rect 19300 9460 19306 9472
rect 19705 9469 19717 9472
rect 19751 9469 19763 9503
rect 19705 9463 19763 9469
rect 20346 9460 20352 9512
rect 20404 9460 20410 9512
rect 22922 9500 22928 9512
rect 21652 9472 22928 9500
rect 20533 9435 20591 9441
rect 18708 9404 20484 9432
rect 20456 9376 20484 9404
rect 20533 9401 20545 9435
rect 20579 9432 20591 9435
rect 21269 9435 21327 9441
rect 21269 9432 21281 9435
rect 20579 9404 21281 9432
rect 20579 9401 20591 9404
rect 20533 9395 20591 9401
rect 21269 9401 21281 9404
rect 21315 9401 21327 9435
rect 21269 9395 21327 9401
rect 13320 9336 14504 9364
rect 15197 9367 15255 9373
rect 13320 9324 13326 9336
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15746 9364 15752 9376
rect 15243 9336 15752 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15746 9324 15752 9336
rect 15804 9364 15810 9376
rect 15933 9367 15991 9373
rect 15933 9364 15945 9367
rect 15804 9336 15945 9364
rect 15804 9324 15810 9336
rect 15933 9333 15945 9336
rect 15979 9333 15991 9367
rect 15933 9327 15991 9333
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 17405 9367 17463 9373
rect 17405 9364 17417 9367
rect 16724 9336 17417 9364
rect 16724 9324 16730 9336
rect 17405 9333 17417 9336
rect 17451 9333 17463 9367
rect 17405 9327 17463 9333
rect 17586 9324 17592 9376
rect 17644 9364 17650 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17644 9336 17785 9364
rect 17644 9324 17650 9336
rect 17773 9333 17785 9336
rect 17819 9364 17831 9367
rect 18509 9367 18567 9373
rect 18509 9364 18521 9367
rect 17819 9336 18521 9364
rect 17819 9333 17831 9336
rect 17773 9327 17831 9333
rect 18509 9333 18521 9336
rect 18555 9364 18567 9367
rect 19153 9367 19211 9373
rect 19153 9364 19165 9367
rect 18555 9336 19165 9364
rect 18555 9333 18567 9336
rect 18509 9327 18567 9333
rect 19153 9333 19165 9336
rect 19199 9364 19211 9367
rect 19334 9364 19340 9376
rect 19199 9336 19340 9364
rect 19199 9333 19211 9336
rect 19153 9327 19211 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 20438 9324 20444 9376
rect 20496 9324 20502 9376
rect 20898 9324 20904 9376
rect 20956 9324 20962 9376
rect 21361 9367 21419 9373
rect 21361 9333 21373 9367
rect 21407 9364 21419 9367
rect 21652 9364 21680 9472
rect 22922 9460 22928 9472
rect 22980 9460 22986 9512
rect 23017 9503 23075 9509
rect 23017 9469 23029 9503
rect 23063 9500 23075 9503
rect 23750 9500 23756 9512
rect 23063 9472 23756 9500
rect 23063 9469 23075 9472
rect 23017 9463 23075 9469
rect 23750 9460 23756 9472
rect 23808 9460 23814 9512
rect 23842 9460 23848 9512
rect 23900 9460 23906 9512
rect 21726 9392 21732 9444
rect 21784 9432 21790 9444
rect 22186 9432 22192 9444
rect 21784 9404 22192 9432
rect 21784 9392 21790 9404
rect 22186 9392 22192 9404
rect 22244 9432 22250 9444
rect 25406 9432 25412 9444
rect 22244 9404 24532 9432
rect 25346 9404 25412 9432
rect 22244 9392 22250 9404
rect 21407 9336 21680 9364
rect 21407 9333 21419 9336
rect 21361 9327 21419 9333
rect 21818 9324 21824 9376
rect 21876 9324 21882 9376
rect 22646 9324 22652 9376
rect 22704 9364 22710 9376
rect 22925 9367 22983 9373
rect 22925 9364 22937 9367
rect 22704 9336 22937 9364
rect 22704 9324 22710 9336
rect 22925 9333 22937 9336
rect 22971 9333 22983 9367
rect 24504 9364 24532 9404
rect 25406 9392 25412 9404
rect 25464 9392 25470 9444
rect 27154 9392 27160 9444
rect 27212 9432 27218 9444
rect 27249 9435 27307 9441
rect 27249 9432 27261 9435
rect 27212 9404 27261 9432
rect 27212 9392 27218 9404
rect 27249 9401 27261 9404
rect 27295 9401 27307 9435
rect 28534 9432 28540 9444
rect 28474 9404 28540 9432
rect 27249 9395 27307 9401
rect 28534 9392 28540 9404
rect 28592 9392 28598 9444
rect 26326 9364 26332 9376
rect 24504 9336 26332 9364
rect 22925 9327 22983 9333
rect 26326 9324 26332 9336
rect 26384 9324 26390 9376
rect 26786 9324 26792 9376
rect 26844 9364 26850 9376
rect 28644 9364 28672 9608
rect 33962 9596 33968 9608
rect 34020 9596 34026 9648
rect 28994 9528 29000 9580
rect 29052 9528 29058 9580
rect 29546 9528 29552 9580
rect 29604 9568 29610 9580
rect 30929 9571 30987 9577
rect 30929 9568 30941 9571
rect 29604 9540 30941 9568
rect 29604 9528 29610 9540
rect 30929 9537 30941 9540
rect 30975 9537 30987 9571
rect 30929 9531 30987 9537
rect 29086 9460 29092 9512
rect 29144 9500 29150 9512
rect 30193 9503 30251 9509
rect 30193 9500 30205 9503
rect 29144 9472 30205 9500
rect 29144 9460 29150 9472
rect 30193 9469 30205 9472
rect 30239 9469 30251 9503
rect 30193 9463 30251 9469
rect 29181 9435 29239 9441
rect 29181 9401 29193 9435
rect 29227 9432 29239 9435
rect 29641 9435 29699 9441
rect 29641 9432 29653 9435
rect 29227 9404 29653 9432
rect 29227 9401 29239 9404
rect 29181 9395 29239 9401
rect 29641 9401 29653 9404
rect 29687 9401 29699 9435
rect 29641 9395 29699 9401
rect 26844 9336 28672 9364
rect 26844 9324 26850 9336
rect 28718 9324 28724 9376
rect 28776 9324 28782 9376
rect 28810 9324 28816 9376
rect 28868 9364 28874 9376
rect 29089 9367 29147 9373
rect 29089 9364 29101 9367
rect 28868 9336 29101 9364
rect 28868 9324 28874 9336
rect 29089 9333 29101 9336
rect 29135 9364 29147 9367
rect 30377 9367 30435 9373
rect 30377 9364 30389 9367
rect 29135 9336 30389 9364
rect 29135 9333 29147 9336
rect 29089 9327 29147 9333
rect 30377 9333 30389 9336
rect 30423 9333 30435 9367
rect 30377 9327 30435 9333
rect 2760 9274 34316 9296
rect 2760 9222 7210 9274
rect 7262 9222 7274 9274
rect 7326 9222 7338 9274
rect 7390 9222 7402 9274
rect 7454 9222 7466 9274
rect 7518 9222 15099 9274
rect 15151 9222 15163 9274
rect 15215 9222 15227 9274
rect 15279 9222 15291 9274
rect 15343 9222 15355 9274
rect 15407 9222 22988 9274
rect 23040 9222 23052 9274
rect 23104 9222 23116 9274
rect 23168 9222 23180 9274
rect 23232 9222 23244 9274
rect 23296 9222 30877 9274
rect 30929 9222 30941 9274
rect 30993 9222 31005 9274
rect 31057 9222 31069 9274
rect 31121 9222 31133 9274
rect 31185 9222 34316 9274
rect 2760 9200 34316 9222
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 4617 9163 4675 9169
rect 4617 9160 4629 9163
rect 4304 9132 4629 9160
rect 4304 9120 4310 9132
rect 4617 9129 4629 9132
rect 4663 9129 4675 9163
rect 7006 9160 7012 9172
rect 4617 9123 4675 9129
rect 6104 9132 7012 9160
rect 3234 9052 3240 9104
rect 3292 9092 3298 9104
rect 5994 9092 6000 9104
rect 3292 9064 6000 9092
rect 3292 9052 3298 9064
rect 5994 9052 6000 9064
rect 6052 9052 6058 9104
rect 4430 8984 4436 9036
rect 4488 9024 4494 9036
rect 4525 9027 4583 9033
rect 4525 9024 4537 9027
rect 4488 8996 4537 9024
rect 4488 8984 4494 8996
rect 4525 8993 4537 8996
rect 4571 8993 4583 9027
rect 4525 8987 4583 8993
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4540 8888 4568 8987
rect 5350 8984 5356 9036
rect 5408 8984 5414 9036
rect 6104 9033 6132 9132
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 9677 9163 9735 9169
rect 9677 9129 9689 9163
rect 9723 9160 9735 9163
rect 9723 9132 9812 9160
rect 9723 9129 9735 9132
rect 9677 9123 9735 9129
rect 9784 9104 9812 9132
rect 10226 9120 10232 9172
rect 10284 9120 10290 9172
rect 10410 9120 10416 9172
rect 10468 9169 10474 9172
rect 10468 9163 10517 9169
rect 10468 9129 10471 9163
rect 10505 9129 10517 9163
rect 10468 9123 10517 9129
rect 10468 9120 10474 9123
rect 10686 9120 10692 9172
rect 10744 9160 10750 9172
rect 13262 9160 13268 9172
rect 10744 9132 13268 9160
rect 10744 9120 10750 9132
rect 13262 9120 13268 9132
rect 13320 9120 13326 9172
rect 17752 9163 17810 9169
rect 17752 9160 17764 9163
rect 17696 9132 17764 9160
rect 8113 9095 8171 9101
rect 8113 9092 8125 9095
rect 7590 9064 8125 9092
rect 8113 9061 8125 9064
rect 8159 9061 8171 9095
rect 8113 9055 8171 9061
rect 9766 9052 9772 9104
rect 9824 9052 9830 9104
rect 6089 9027 6147 9033
rect 6089 8993 6101 9027
rect 6135 8993 6147 9027
rect 6089 8987 6147 8993
rect 8202 8984 8208 9036
rect 8260 8984 8266 9036
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8536 8996 9229 9024
rect 8536 8984 8542 8996
rect 9217 8993 9229 8996
rect 9263 9024 9275 9027
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 9263 8996 9873 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 9861 8993 9873 8996
rect 9907 9024 9919 9027
rect 10244 9024 10272 9120
rect 11514 9052 11520 9104
rect 11572 9052 11578 9104
rect 14182 9052 14188 9104
rect 14240 9052 14246 9104
rect 14366 9052 14372 9104
rect 14424 9092 14430 9104
rect 14424 9064 14964 9092
rect 14424 9052 14430 9064
rect 14936 9036 14964 9064
rect 9907 8996 10272 9024
rect 11885 9027 11943 9033
rect 9907 8993 9919 8996
rect 9861 8987 9919 8993
rect 11885 8993 11897 9027
rect 11931 9024 11943 9027
rect 11931 8996 13492 9024
rect 11931 8993 11943 8996
rect 11885 8987 11943 8993
rect 5258 8916 5264 8968
rect 5316 8916 5322 8968
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 9493 8959 9551 8965
rect 9493 8925 9505 8959
rect 9539 8956 9551 8959
rect 9950 8956 9956 8968
rect 9539 8928 9956 8956
rect 9539 8925 9551 8928
rect 9493 8919 9551 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 12250 8916 12256 8968
rect 12308 8916 12314 8968
rect 13464 8956 13492 8996
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 17129 9027 17187 9033
rect 17129 8993 17141 9027
rect 17175 9024 17187 9027
rect 17586 9024 17592 9036
rect 17175 8996 17592 9024
rect 17175 8993 17187 8996
rect 17129 8987 17187 8993
rect 17586 8984 17592 8996
rect 17644 9024 17650 9036
rect 17696 9024 17724 9132
rect 17752 9129 17764 9132
rect 17798 9129 17810 9163
rect 17752 9123 17810 9129
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 18104 9132 20300 9160
rect 18104 9120 18110 9132
rect 17862 9052 17868 9104
rect 17920 9092 17926 9104
rect 17957 9095 18015 9101
rect 17957 9092 17969 9095
rect 17920 9064 17969 9092
rect 17920 9052 17926 9064
rect 17957 9061 17969 9064
rect 18003 9061 18015 9095
rect 20272 9092 20300 9132
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 20404 9132 20453 9160
rect 20404 9120 20410 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 20809 9163 20867 9169
rect 20809 9160 20821 9163
rect 20772 9132 20821 9160
rect 20772 9120 20778 9132
rect 20809 9129 20821 9132
rect 20855 9129 20867 9163
rect 24857 9163 24915 9169
rect 20809 9123 20867 9129
rect 22066 9132 23520 9160
rect 22066 9092 22094 9132
rect 23492 9101 23520 9132
rect 24857 9129 24869 9163
rect 24903 9160 24915 9163
rect 25130 9160 25136 9172
rect 24903 9132 25136 9160
rect 24903 9129 24915 9132
rect 24857 9123 24915 9129
rect 25130 9120 25136 9132
rect 25188 9120 25194 9172
rect 25225 9163 25283 9169
rect 25225 9129 25237 9163
rect 25271 9160 25283 9163
rect 25682 9160 25688 9172
rect 25271 9132 25688 9160
rect 25271 9129 25283 9132
rect 25225 9123 25283 9129
rect 25682 9120 25688 9132
rect 25740 9120 25746 9172
rect 26234 9160 26240 9172
rect 25884 9132 26240 9160
rect 20272 9064 22094 9092
rect 23477 9095 23535 9101
rect 17957 9055 18015 9061
rect 23477 9061 23489 9095
rect 23523 9061 23535 9095
rect 25884 9092 25912 9132
rect 26234 9120 26240 9132
rect 26292 9120 26298 9172
rect 26326 9120 26332 9172
rect 26384 9160 26390 9172
rect 27890 9160 27896 9172
rect 26384 9132 27896 9160
rect 26384 9120 26390 9132
rect 27890 9120 27896 9132
rect 27948 9120 27954 9172
rect 28718 9120 28724 9172
rect 28776 9120 28782 9172
rect 29546 9120 29552 9172
rect 29604 9120 29610 9172
rect 29730 9120 29736 9172
rect 29788 9120 29794 9172
rect 23477 9055 23535 9061
rect 24688 9064 25912 9092
rect 28736 9092 28764 9120
rect 29748 9092 29776 9120
rect 31573 9095 31631 9101
rect 31573 9092 31585 9095
rect 28736 9064 28948 9092
rect 17644 8996 17724 9024
rect 17644 8984 17650 8996
rect 18782 8984 18788 9036
rect 18840 8984 18846 9036
rect 19610 8984 19616 9036
rect 19668 9033 19674 9036
rect 19668 9027 19696 9033
rect 19684 8993 19696 9027
rect 19668 8987 19696 8993
rect 19668 8984 19674 8987
rect 20898 8984 20904 9036
rect 20956 8984 20962 9036
rect 21545 9027 21603 9033
rect 21545 9024 21557 9027
rect 21192 8996 21557 9024
rect 14550 8956 14556 8968
rect 13464 8928 14556 8956
rect 14550 8916 14556 8928
rect 14608 8916 14614 8968
rect 14645 8959 14703 8965
rect 14645 8925 14657 8959
rect 14691 8956 14703 8959
rect 16761 8959 16819 8965
rect 14691 8928 14872 8956
rect 14691 8925 14703 8928
rect 14645 8919 14703 8925
rect 4540 8860 5396 8888
rect 5368 8832 5396 8860
rect 14844 8832 14872 8928
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 16942 8956 16948 8968
rect 16807 8928 16948 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 16942 8916 16948 8928
rect 17000 8956 17006 8968
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 17000 8928 17509 8956
rect 17000 8916 17006 8928
rect 17497 8925 17509 8928
rect 17543 8956 17555 8959
rect 17543 8928 18000 8956
rect 17543 8925 17555 8928
rect 17497 8919 17555 8925
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 17126 8888 17132 8900
rect 16908 8860 17132 8888
rect 16908 8848 16914 8860
rect 17126 8848 17132 8860
rect 17184 8888 17190 8900
rect 17589 8891 17647 8897
rect 17589 8888 17601 8891
rect 17184 8860 17601 8888
rect 17184 8848 17190 8860
rect 17589 8857 17601 8860
rect 17635 8857 17647 8891
rect 17972 8888 18000 8928
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 18564 8928 18613 8956
rect 18564 8916 18570 8928
rect 18601 8925 18613 8928
rect 18647 8925 18659 8959
rect 18601 8919 18659 8925
rect 19150 8916 19156 8968
rect 19208 8916 19214 8968
rect 19518 8916 19524 8968
rect 19576 8916 19582 8968
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8956 19855 8959
rect 19843 8928 20208 8956
rect 19843 8925 19855 8928
rect 19797 8919 19855 8925
rect 19168 8888 19196 8916
rect 17972 8860 19196 8888
rect 19245 8891 19303 8897
rect 17589 8851 17647 8857
rect 19245 8857 19257 8891
rect 19291 8888 19303 8891
rect 19334 8888 19340 8900
rect 19291 8860 19340 8888
rect 19291 8857 19303 8860
rect 19245 8851 19303 8857
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 3605 8823 3663 8829
rect 3605 8820 3617 8823
rect 3476 8792 3617 8820
rect 3476 8780 3482 8792
rect 3605 8789 3617 8792
rect 3651 8789 3663 8823
rect 3605 8783 3663 8789
rect 4430 8780 4436 8832
rect 4488 8780 4494 8832
rect 5350 8780 5356 8832
rect 5408 8780 5414 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5960 8792 6009 8820
rect 5960 8780 5966 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 7837 8823 7895 8829
rect 7837 8789 7849 8823
rect 7883 8820 7895 8823
rect 8018 8820 8024 8832
rect 7883 8792 8024 8820
rect 7883 8789 7895 8792
rect 7837 8783 7895 8789
rect 8018 8780 8024 8792
rect 8076 8780 8082 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 9306 8820 9312 8832
rect 8619 8792 9312 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 9306 8780 9312 8792
rect 9364 8780 9370 8832
rect 9490 8780 9496 8832
rect 9548 8780 9554 8832
rect 13173 8823 13231 8829
rect 13173 8789 13185 8823
rect 13219 8820 13231 8823
rect 13906 8820 13912 8832
rect 13219 8792 13912 8820
rect 13219 8789 13231 8792
rect 13173 8783 13231 8789
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 14826 8780 14832 8832
rect 14884 8780 14890 8832
rect 15473 8823 15531 8829
rect 15473 8789 15485 8823
rect 15519 8820 15531 8823
rect 15930 8820 15936 8832
rect 15519 8792 15936 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 15930 8780 15936 8792
rect 15988 8780 15994 8832
rect 16574 8780 16580 8832
rect 16632 8820 16638 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 16632 8792 17785 8820
rect 16632 8780 16638 8792
rect 17773 8789 17785 8792
rect 17819 8820 17831 8823
rect 18138 8820 18144 8832
rect 17819 8792 18144 8820
rect 17819 8789 17831 8792
rect 17773 8783 17831 8789
rect 18138 8780 18144 8792
rect 18196 8780 18202 8832
rect 18966 8780 18972 8832
rect 19024 8820 19030 8832
rect 20180 8820 20208 8928
rect 20916 8888 20944 8984
rect 21192 8968 21220 8996
rect 21545 8993 21557 8996
rect 21591 8993 21603 9027
rect 23566 9024 23572 9036
rect 22954 8996 23572 9024
rect 21545 8987 21603 8993
rect 23566 8984 23572 8996
rect 23624 8984 23630 9036
rect 21174 8916 21180 8968
rect 21232 8916 21238 8968
rect 21361 8959 21419 8965
rect 21361 8925 21373 8959
rect 21407 8925 21419 8959
rect 21361 8919 21419 8925
rect 21376 8888 21404 8919
rect 21818 8916 21824 8968
rect 21876 8916 21882 8968
rect 24688 8965 24716 9064
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 24912 8996 25084 9024
rect 24912 8984 24918 8996
rect 24121 8959 24179 8965
rect 24121 8925 24133 8959
rect 24167 8925 24179 8959
rect 24121 8919 24179 8925
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8925 24731 8959
rect 24673 8919 24731 8925
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8956 24823 8959
rect 24946 8956 24952 8968
rect 24811 8928 24952 8956
rect 24811 8925 24823 8928
rect 24765 8919 24823 8925
rect 20916 8860 21404 8888
rect 23293 8891 23351 8897
rect 23293 8857 23305 8891
rect 23339 8888 23351 8891
rect 23934 8888 23940 8900
rect 23339 8860 23940 8888
rect 23339 8857 23351 8860
rect 23293 8851 23351 8857
rect 23934 8848 23940 8860
rect 23992 8848 23998 8900
rect 22002 8820 22008 8832
rect 19024 8792 22008 8820
rect 19024 8780 19030 8792
rect 22002 8780 22008 8792
rect 22060 8780 22066 8832
rect 24136 8820 24164 8919
rect 24946 8916 24952 8928
rect 25004 8916 25010 8968
rect 25056 8956 25084 8996
rect 25222 8984 25228 9036
rect 25280 9024 25286 9036
rect 25317 9027 25375 9033
rect 25317 9024 25329 9027
rect 25280 8996 25329 9024
rect 25280 8984 25286 8996
rect 25317 8993 25329 8996
rect 25363 8993 25375 9027
rect 25317 8987 25375 8993
rect 25406 8984 25412 9036
rect 25464 8984 25470 9036
rect 26786 9033 26792 9036
rect 26743 9027 26792 9033
rect 26743 8993 26755 9027
rect 26789 8993 26792 9027
rect 26743 8987 26792 8993
rect 26786 8984 26792 8987
rect 26844 8984 26850 9036
rect 28920 9033 28948 9064
rect 29656 9064 29776 9092
rect 31142 9064 31585 9092
rect 29656 9033 29684 9064
rect 31573 9061 31585 9064
rect 31619 9061 31631 9095
rect 31573 9055 31631 9061
rect 28813 9027 28871 9033
rect 28813 8993 28825 9027
rect 28859 8993 28871 9027
rect 28813 8987 28871 8993
rect 28905 9027 28963 9033
rect 28905 8993 28917 9027
rect 28951 8993 28963 9027
rect 28905 8987 28963 8993
rect 29641 9027 29699 9033
rect 29641 8993 29653 9027
rect 29687 8993 29699 9027
rect 31665 9027 31723 9033
rect 31665 9024 31677 9027
rect 29641 8987 29699 8993
rect 31128 8996 31677 9024
rect 25682 8956 25688 8968
rect 25056 8928 25688 8956
rect 25682 8916 25688 8928
rect 25740 8916 25746 8968
rect 25866 8916 25872 8968
rect 25924 8916 25930 8968
rect 26602 8916 26608 8968
rect 26660 8916 26666 8968
rect 26878 8916 26884 8968
rect 26936 8916 26942 8968
rect 28442 8916 28448 8968
rect 28500 8916 28506 8968
rect 28534 8916 28540 8968
rect 28592 8956 28598 8968
rect 28721 8959 28779 8965
rect 28721 8956 28733 8959
rect 28592 8928 28733 8956
rect 28592 8916 28598 8928
rect 28721 8925 28733 8928
rect 28767 8925 28779 8959
rect 28721 8919 28779 8925
rect 25314 8848 25320 8900
rect 25372 8888 25378 8900
rect 26329 8891 26387 8897
rect 26329 8888 26341 8891
rect 25372 8860 26341 8888
rect 25372 8848 25378 8860
rect 26329 8857 26341 8860
rect 26375 8857 26387 8891
rect 27801 8891 27859 8897
rect 27801 8888 27813 8891
rect 26329 8851 26387 8857
rect 27264 8860 27813 8888
rect 27264 8820 27292 8860
rect 27801 8857 27813 8860
rect 27847 8857 27859 8891
rect 27801 8851 27859 8857
rect 24136 8792 27292 8820
rect 27522 8780 27528 8832
rect 27580 8780 27586 8832
rect 27614 8780 27620 8832
rect 27672 8820 27678 8832
rect 28828 8820 28856 8987
rect 29914 8916 29920 8968
rect 29972 8916 29978 8968
rect 30650 8820 30656 8832
rect 27672 8792 30656 8820
rect 27672 8780 27678 8792
rect 30650 8780 30656 8792
rect 30708 8820 30714 8832
rect 31128 8820 31156 8996
rect 31665 8993 31677 8996
rect 31711 8993 31723 9027
rect 31665 8987 31723 8993
rect 32582 8916 32588 8968
rect 32640 8916 32646 8968
rect 31389 8891 31447 8897
rect 31389 8857 31401 8891
rect 31435 8888 31447 8891
rect 33410 8888 33416 8900
rect 31435 8860 33416 8888
rect 31435 8857 31447 8860
rect 31389 8851 31447 8857
rect 33410 8848 33416 8860
rect 33468 8848 33474 8900
rect 30708 8792 31156 8820
rect 30708 8780 30714 8792
rect 32030 8780 32036 8832
rect 32088 8780 32094 8832
rect 2760 8730 34316 8752
rect 2760 8678 6550 8730
rect 6602 8678 6614 8730
rect 6666 8678 6678 8730
rect 6730 8678 6742 8730
rect 6794 8678 6806 8730
rect 6858 8678 14439 8730
rect 14491 8678 14503 8730
rect 14555 8678 14567 8730
rect 14619 8678 14631 8730
rect 14683 8678 14695 8730
rect 14747 8678 22328 8730
rect 22380 8678 22392 8730
rect 22444 8678 22456 8730
rect 22508 8678 22520 8730
rect 22572 8678 22584 8730
rect 22636 8678 30217 8730
rect 30269 8678 30281 8730
rect 30333 8678 30345 8730
rect 30397 8678 30409 8730
rect 30461 8678 30473 8730
rect 30525 8678 34316 8730
rect 2760 8656 34316 8678
rect 3316 8619 3374 8625
rect 3316 8585 3328 8619
rect 3362 8616 3374 8619
rect 3418 8616 3424 8628
rect 3362 8588 3424 8616
rect 3362 8585 3374 8588
rect 3316 8579 3374 8585
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 5074 8576 5080 8628
rect 5132 8576 5138 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5316 8588 5457 8616
rect 5316 8576 5322 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 5445 8579 5503 8585
rect 5902 8576 5908 8628
rect 5960 8616 5966 8628
rect 6929 8619 6987 8625
rect 6929 8616 6941 8619
rect 5960 8588 6941 8616
rect 5960 8576 5966 8588
rect 6929 8585 6941 8588
rect 6975 8585 6987 8619
rect 6929 8579 6987 8585
rect 7098 8576 7104 8628
rect 7156 8576 7162 8628
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 10781 8619 10839 8625
rect 10781 8616 10793 8619
rect 8352 8588 10793 8616
rect 8352 8576 8358 8588
rect 10781 8585 10793 8588
rect 10827 8616 10839 8619
rect 13078 8616 13084 8628
rect 10827 8588 13084 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 13078 8576 13084 8588
rect 13136 8616 13142 8628
rect 13722 8616 13728 8628
rect 13136 8588 13728 8616
rect 13136 8576 13142 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 14182 8576 14188 8628
rect 14240 8576 14246 8628
rect 14645 8619 14703 8625
rect 14645 8585 14657 8619
rect 14691 8616 14703 8619
rect 14826 8616 14832 8628
rect 14691 8588 14832 8616
rect 14691 8585 14703 8588
rect 14645 8579 14703 8585
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15381 8619 15439 8625
rect 15381 8585 15393 8619
rect 15427 8616 15439 8619
rect 18509 8619 18567 8625
rect 15427 8585 15440 8616
rect 15381 8579 15440 8585
rect 18509 8585 18521 8619
rect 18555 8616 18567 8619
rect 18874 8616 18880 8628
rect 18555 8588 18880 8616
rect 18555 8585 18567 8588
rect 18509 8579 18567 8585
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 4338 8480 4344 8492
rect 3099 8452 4344 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 7116 8480 7144 8576
rect 11514 8508 11520 8560
rect 11572 8508 11578 8560
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 12158 8548 12164 8560
rect 11848 8520 12164 8548
rect 11848 8508 11854 8520
rect 12158 8508 12164 8520
rect 12216 8548 12222 8560
rect 12253 8551 12311 8557
rect 12253 8548 12265 8551
rect 12216 8520 12265 8548
rect 12216 8508 12222 8520
rect 12253 8517 12265 8520
rect 12299 8517 12311 8551
rect 12253 8511 12311 8517
rect 13909 8551 13967 8557
rect 13909 8517 13921 8551
rect 13955 8548 13967 8551
rect 13955 8520 14044 8548
rect 13955 8517 13967 8520
rect 13909 8511 13967 8517
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 7116 8452 7205 8480
rect 7193 8449 7205 8452
rect 7239 8480 7251 8483
rect 7377 8483 7435 8489
rect 7377 8480 7389 8483
rect 7239 8452 7389 8480
rect 7239 8449 7251 8452
rect 7193 8443 7251 8449
rect 7377 8449 7389 8452
rect 7423 8449 7435 8483
rect 7377 8443 7435 8449
rect 9122 8440 9128 8492
rect 9180 8480 9186 8492
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9180 8452 9781 8480
rect 9180 8440 9186 8452
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 13081 8483 13139 8489
rect 13081 8449 13093 8483
rect 13127 8480 13139 8483
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 13127 8452 13369 8480
rect 13127 8449 13139 8452
rect 13081 8443 13139 8449
rect 13357 8449 13369 8452
rect 13403 8480 13415 8483
rect 13814 8480 13820 8492
rect 13403 8452 13820 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14016 8489 14044 8520
rect 14001 8483 14059 8489
rect 14001 8449 14013 8483
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 14200 8480 14228 8576
rect 14829 8483 14887 8489
rect 14829 8480 14841 8483
rect 14200 8452 14841 8480
rect 14829 8449 14841 8452
rect 14875 8449 14887 8483
rect 14829 8443 14887 8449
rect 4430 8372 4436 8424
rect 4488 8372 4494 8424
rect 5810 8372 5816 8424
rect 5868 8372 5874 8424
rect 9674 8412 9680 8424
rect 8786 8384 9680 8412
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8412 11667 8415
rect 12066 8412 12072 8424
rect 11655 8384 12072 8412
rect 11655 8381 11667 8384
rect 11609 8375 11667 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 13538 8372 13544 8424
rect 13596 8372 13602 8424
rect 14108 8412 14136 8440
rect 14921 8415 14979 8421
rect 14921 8412 14933 8415
rect 14108 8384 14933 8412
rect 14921 8381 14933 8384
rect 14967 8381 14979 8415
rect 15412 8412 15440 8579
rect 18874 8576 18880 8588
rect 18932 8576 18938 8628
rect 19245 8619 19303 8625
rect 19245 8585 19257 8619
rect 19291 8616 19303 8619
rect 19334 8616 19340 8628
rect 19291 8588 19340 8616
rect 19291 8585 19303 8588
rect 19245 8579 19303 8585
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 19610 8576 19616 8628
rect 19668 8616 19674 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 19668 8588 20545 8616
rect 19668 8576 19674 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 21726 8616 21732 8628
rect 20533 8579 20591 8585
rect 20732 8588 21732 8616
rect 16942 8548 16948 8560
rect 16776 8520 16948 8548
rect 15930 8440 15936 8492
rect 15988 8480 15994 8492
rect 16666 8480 16672 8492
rect 15988 8452 16672 8480
rect 15988 8440 15994 8452
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16776 8489 16804 8520
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17405 8551 17463 8557
rect 17405 8517 17417 8551
rect 17451 8517 17463 8551
rect 18966 8548 18972 8560
rect 17405 8511 17463 8517
rect 17788 8520 18972 8548
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8449 16819 8483
rect 16761 8443 16819 8449
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 17218 8412 17224 8424
rect 17276 8421 17282 8424
rect 17276 8415 17304 8421
rect 15412 8384 17224 8412
rect 14921 8375 14979 8381
rect 17218 8372 17224 8384
rect 17292 8381 17304 8415
rect 17420 8412 17448 8511
rect 17788 8492 17816 8520
rect 18966 8508 18972 8520
rect 19024 8548 19030 8560
rect 19024 8520 19380 8548
rect 19024 8508 19030 8520
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 18138 8480 18144 8492
rect 17880 8452 18144 8480
rect 17880 8421 17908 8452
rect 18138 8440 18144 8452
rect 18196 8480 18202 8492
rect 19242 8480 19248 8492
rect 18196 8452 19248 8480
rect 18196 8440 18202 8452
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 17681 8415 17739 8421
rect 17681 8412 17693 8415
rect 17420 8384 17693 8412
rect 17276 8375 17304 8381
rect 17681 8381 17693 8384
rect 17727 8381 17739 8415
rect 17681 8375 17739 8381
rect 17865 8415 17923 8421
rect 17865 8381 17877 8415
rect 17911 8381 17923 8415
rect 17865 8375 17923 8381
rect 17276 8372 17282 8375
rect 17954 8372 17960 8424
rect 18012 8372 18018 8424
rect 7650 8304 7656 8356
rect 7708 8304 7714 8356
rect 9490 8304 9496 8356
rect 9548 8344 9554 8356
rect 10229 8347 10287 8353
rect 10229 8344 10241 8347
rect 9548 8316 10241 8344
rect 9548 8304 9554 8316
rect 10229 8313 10241 8316
rect 10275 8344 10287 8347
rect 12526 8344 12532 8356
rect 10275 8316 12532 8344
rect 10275 8313 10287 8316
rect 10229 8307 10287 8313
rect 12526 8304 12532 8316
rect 12584 8304 12590 8356
rect 13449 8347 13507 8353
rect 13449 8313 13461 8347
rect 13495 8344 13507 8347
rect 13906 8344 13912 8356
rect 13495 8316 13912 8344
rect 13495 8313 13507 8316
rect 13449 8307 13507 8313
rect 13906 8304 13912 8316
rect 13964 8304 13970 8356
rect 15197 8347 15255 8353
rect 15197 8313 15209 8347
rect 15243 8313 15255 8347
rect 15197 8307 15255 8313
rect 4798 8236 4804 8288
rect 4856 8236 4862 8288
rect 6178 8236 6184 8288
rect 6236 8276 6242 8288
rect 6546 8276 6552 8288
rect 6236 8248 6552 8276
rect 6236 8236 6242 8248
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 9214 8236 9220 8288
rect 9272 8236 9278 8288
rect 14918 8236 14924 8288
rect 14976 8276 14982 8288
rect 15212 8276 15240 8307
rect 16574 8304 16580 8356
rect 16632 8344 16638 8356
rect 16669 8347 16727 8353
rect 16669 8344 16681 8347
rect 16632 8316 16681 8344
rect 16632 8304 16638 8316
rect 16669 8313 16681 8316
rect 16715 8313 16727 8347
rect 16669 8307 16727 8313
rect 17037 8347 17095 8353
rect 17037 8313 17049 8347
rect 17083 8344 17095 8347
rect 19260 8344 19288 8440
rect 19352 8412 19380 8520
rect 19455 8483 19513 8489
rect 19455 8449 19467 8483
rect 19501 8480 19513 8483
rect 20732 8480 20760 8588
rect 21726 8576 21732 8588
rect 21784 8576 21790 8628
rect 22094 8576 22100 8628
rect 22152 8616 22158 8628
rect 22152 8588 22784 8616
rect 22152 8576 22158 8588
rect 20806 8508 20812 8560
rect 20864 8548 20870 8560
rect 22756 8548 22784 8588
rect 22830 8576 22836 8628
rect 22888 8616 22894 8628
rect 23017 8619 23075 8625
rect 23017 8616 23029 8619
rect 22888 8588 23029 8616
rect 22888 8576 22894 8588
rect 23017 8585 23029 8588
rect 23063 8585 23075 8619
rect 23017 8579 23075 8585
rect 23308 8588 23520 8616
rect 23308 8548 23336 8588
rect 20864 8520 21312 8548
rect 22756 8520 23336 8548
rect 20864 8508 20870 8520
rect 21284 8489 21312 8520
rect 23382 8508 23388 8560
rect 23440 8508 23446 8560
rect 23492 8548 23520 8588
rect 23566 8576 23572 8628
rect 23624 8576 23630 8628
rect 24210 8616 24216 8628
rect 23776 8588 24216 8616
rect 23776 8548 23804 8588
rect 24210 8576 24216 8588
rect 24268 8616 24274 8628
rect 24268 8588 25176 8616
rect 24268 8576 24274 8588
rect 23492 8520 23804 8548
rect 25148 8548 25176 8588
rect 25314 8576 25320 8628
rect 25372 8576 25378 8628
rect 25682 8576 25688 8628
rect 25740 8616 25746 8628
rect 26237 8619 26295 8625
rect 26237 8616 26249 8619
rect 25740 8588 26249 8616
rect 25740 8576 25746 8588
rect 26237 8585 26249 8588
rect 26283 8585 26295 8619
rect 26237 8579 26295 8585
rect 26326 8576 26332 8628
rect 26384 8616 26390 8628
rect 27341 8619 27399 8625
rect 26384 8588 27292 8616
rect 26384 8576 26390 8588
rect 25593 8551 25651 8557
rect 25593 8548 25605 8551
rect 25148 8520 25605 8548
rect 25593 8517 25605 8520
rect 25639 8548 25651 8551
rect 26694 8548 26700 8560
rect 25639 8520 26700 8548
rect 25639 8517 25651 8520
rect 25593 8511 25651 8517
rect 26694 8508 26700 8520
rect 26752 8548 26758 8560
rect 26878 8548 26884 8560
rect 26752 8520 26884 8548
rect 26752 8508 26758 8520
rect 26878 8508 26884 8520
rect 26936 8508 26942 8560
rect 27264 8548 27292 8588
rect 27341 8585 27353 8619
rect 27387 8616 27399 8619
rect 27430 8616 27436 8628
rect 27387 8588 27436 8616
rect 27387 8585 27399 8588
rect 27341 8579 27399 8585
rect 27430 8576 27436 8588
rect 27488 8576 27494 8628
rect 28442 8576 28448 8628
rect 28500 8576 28506 8628
rect 28994 8576 29000 8628
rect 29052 8616 29058 8628
rect 29454 8616 29460 8628
rect 29052 8588 29460 8616
rect 29052 8576 29058 8588
rect 29454 8576 29460 8588
rect 29512 8576 29518 8628
rect 29549 8619 29607 8625
rect 29549 8585 29561 8619
rect 29595 8616 29607 8619
rect 29914 8616 29920 8628
rect 29595 8588 29920 8616
rect 29595 8585 29607 8588
rect 29549 8579 29607 8585
rect 29914 8576 29920 8588
rect 29972 8576 29978 8628
rect 32999 8619 33057 8625
rect 32999 8616 33011 8619
rect 30024 8588 33011 8616
rect 28460 8548 28488 8576
rect 30024 8548 30052 8588
rect 32999 8585 33011 8588
rect 33045 8585 33057 8619
rect 32999 8579 33057 8585
rect 33413 8619 33471 8625
rect 33413 8585 33425 8619
rect 33459 8616 33471 8619
rect 33502 8616 33508 8628
rect 33459 8588 33508 8616
rect 33459 8585 33471 8588
rect 33413 8579 33471 8585
rect 33502 8576 33508 8588
rect 33560 8576 33566 8628
rect 27264 8520 28120 8548
rect 28460 8520 30052 8548
rect 19501 8452 20760 8480
rect 21269 8483 21327 8489
rect 19501 8449 19513 8452
rect 19455 8443 19513 8449
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21634 8480 21640 8492
rect 21315 8452 21640 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21634 8440 21640 8452
rect 21692 8440 21698 8492
rect 21726 8440 21732 8492
rect 21784 8440 21790 8492
rect 21818 8440 21824 8492
rect 21876 8480 21882 8492
rect 22143 8483 22201 8489
rect 21876 8452 22048 8480
rect 21876 8440 21882 8452
rect 19613 8415 19671 8421
rect 19613 8412 19625 8415
rect 19352 8384 19625 8412
rect 19613 8381 19625 8384
rect 19659 8381 19671 8415
rect 19613 8375 19671 8381
rect 19794 8372 19800 8424
rect 19852 8372 19858 8424
rect 20530 8372 20536 8424
rect 20588 8372 20594 8424
rect 21082 8372 21088 8424
rect 21140 8372 21146 8424
rect 22020 8421 22048 8452
rect 22143 8449 22155 8483
rect 22189 8480 22201 8483
rect 23106 8480 23112 8492
rect 22189 8452 23112 8480
rect 22189 8449 22201 8452
rect 22143 8443 22201 8449
rect 23106 8440 23112 8452
rect 23164 8440 23170 8492
rect 23400 8480 23428 8508
rect 23400 8452 24992 8480
rect 22005 8415 22063 8421
rect 22005 8381 22017 8415
rect 22051 8381 22063 8415
rect 22005 8375 22063 8381
rect 22278 8372 22284 8424
rect 22336 8372 22342 8424
rect 23676 8421 23704 8452
rect 22925 8415 22983 8421
rect 22925 8381 22937 8415
rect 22971 8412 22983 8415
rect 23201 8415 23259 8421
rect 23201 8412 23213 8415
rect 22971 8384 23213 8412
rect 22971 8381 22983 8384
rect 22925 8375 22983 8381
rect 23201 8381 23213 8384
rect 23247 8381 23259 8415
rect 23201 8375 23259 8381
rect 23293 8415 23351 8421
rect 23293 8381 23305 8415
rect 23339 8381 23351 8415
rect 23293 8375 23351 8381
rect 23661 8415 23719 8421
rect 23661 8381 23673 8415
rect 23707 8381 23719 8415
rect 23661 8375 23719 8381
rect 20073 8347 20131 8353
rect 20073 8344 20085 8347
rect 17083 8316 17724 8344
rect 19260 8316 20085 8344
rect 17083 8313 17095 8316
rect 17037 8307 17095 8313
rect 17696 8288 17724 8316
rect 20073 8313 20085 8316
rect 20119 8313 20131 8347
rect 20548 8344 20576 8372
rect 23308 8344 23336 8375
rect 24854 8372 24860 8424
rect 24912 8372 24918 8424
rect 24964 8412 24992 8452
rect 26896 8452 27752 8480
rect 26896 8424 26924 8452
rect 25222 8412 25228 8424
rect 24964 8384 25228 8412
rect 25222 8372 25228 8384
rect 25280 8372 25286 8424
rect 26326 8372 26332 8424
rect 26384 8412 26390 8424
rect 26510 8412 26516 8424
rect 26384 8384 26516 8412
rect 26384 8372 26390 8384
rect 26510 8372 26516 8384
rect 26568 8372 26574 8424
rect 26878 8372 26884 8424
rect 26936 8372 26942 8424
rect 27062 8372 27068 8424
rect 27120 8412 27126 8424
rect 27430 8412 27436 8424
rect 27120 8384 27436 8412
rect 27120 8372 27126 8384
rect 27430 8372 27436 8384
rect 27488 8372 27494 8424
rect 27522 8372 27528 8424
rect 27580 8372 27586 8424
rect 27617 8415 27675 8421
rect 27617 8381 27629 8415
rect 27663 8381 27675 8415
rect 27724 8412 27752 8452
rect 27890 8440 27896 8492
rect 27948 8480 27954 8492
rect 27985 8483 28043 8489
rect 27985 8480 27997 8483
rect 27948 8452 27997 8480
rect 27948 8440 27954 8452
rect 27985 8449 27997 8452
rect 28031 8449 28043 8483
rect 27985 8443 28043 8449
rect 28092 8421 28120 8520
rect 33778 8508 33784 8560
rect 33836 8508 33842 8560
rect 28166 8440 28172 8492
rect 28224 8480 28230 8492
rect 30561 8483 30619 8489
rect 30561 8480 30573 8483
rect 28224 8452 30573 8480
rect 28224 8440 28230 8452
rect 28077 8415 28135 8421
rect 27724 8384 27844 8412
rect 27617 8375 27675 8381
rect 25682 8344 25688 8356
rect 20548 8316 21312 8344
rect 20073 8307 20131 8313
rect 14976 8248 15240 8276
rect 14976 8236 14982 8248
rect 15378 8236 15384 8288
rect 15436 8285 15442 8288
rect 15436 8279 15455 8285
rect 15443 8245 15455 8279
rect 15436 8239 15455 8245
rect 15436 8236 15442 8239
rect 15562 8236 15568 8288
rect 15620 8236 15626 8288
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17497 8279 17555 8285
rect 17497 8276 17509 8279
rect 17460 8248 17509 8276
rect 17460 8236 17466 8248
rect 17497 8245 17509 8248
rect 17543 8245 17555 8279
rect 17497 8239 17555 8245
rect 17678 8236 17684 8288
rect 17736 8236 17742 8288
rect 19426 8236 19432 8288
rect 19484 8276 19490 8288
rect 20990 8276 20996 8288
rect 19484 8248 20996 8276
rect 19484 8236 19490 8248
rect 20990 8236 20996 8248
rect 21048 8236 21054 8288
rect 21284 8276 21312 8316
rect 23308 8316 25688 8344
rect 23308 8276 23336 8316
rect 25682 8304 25688 8316
rect 25740 8344 25746 8356
rect 27632 8344 27660 8375
rect 27706 8344 27712 8356
rect 25740 8316 27712 8344
rect 25740 8304 25746 8316
rect 27706 8304 27712 8316
rect 27764 8304 27770 8356
rect 27816 8344 27844 8384
rect 28077 8381 28089 8415
rect 28123 8412 28135 8415
rect 28718 8412 28724 8424
rect 28123 8384 28724 8412
rect 28123 8381 28135 8384
rect 28077 8375 28135 8381
rect 28718 8372 28724 8384
rect 28776 8372 28782 8424
rect 28994 8372 29000 8424
rect 29052 8372 29058 8424
rect 29196 8421 29224 8452
rect 30561 8449 30573 8452
rect 30607 8449 30619 8483
rect 30561 8443 30619 8449
rect 31202 8440 31208 8492
rect 31260 8440 31266 8492
rect 29181 8415 29239 8421
rect 29181 8381 29193 8415
rect 29227 8381 29239 8415
rect 29181 8375 29239 8381
rect 29365 8415 29423 8421
rect 29365 8381 29377 8415
rect 29411 8381 29423 8415
rect 29365 8375 29423 8381
rect 28353 8347 28411 8353
rect 28353 8344 28365 8347
rect 27816 8316 28365 8344
rect 28353 8313 28365 8316
rect 28399 8313 28411 8347
rect 28353 8307 28411 8313
rect 28445 8347 28503 8353
rect 28445 8313 28457 8347
rect 28491 8344 28503 8347
rect 29086 8344 29092 8356
rect 28491 8316 29092 8344
rect 28491 8313 28503 8316
rect 28445 8307 28503 8313
rect 21284 8248 23336 8276
rect 24302 8236 24308 8288
rect 24360 8236 24366 8288
rect 24486 8236 24492 8288
rect 24544 8276 24550 8288
rect 26697 8279 26755 8285
rect 26697 8276 26709 8279
rect 24544 8248 26709 8276
rect 24544 8236 24550 8248
rect 26697 8245 26709 8248
rect 26743 8276 26755 8279
rect 26878 8276 26884 8288
rect 26743 8248 26884 8276
rect 26743 8245 26755 8248
rect 26697 8239 26755 8245
rect 26878 8236 26884 8248
rect 26936 8236 26942 8288
rect 26970 8236 26976 8288
rect 27028 8236 27034 8288
rect 27801 8279 27859 8285
rect 27801 8245 27813 8279
rect 27847 8276 27859 8279
rect 28166 8276 28172 8288
rect 27847 8248 28172 8276
rect 27847 8245 27859 8248
rect 27801 8239 27859 8245
rect 28166 8236 28172 8248
rect 28224 8236 28230 8288
rect 28368 8276 28396 8307
rect 29086 8304 29092 8316
rect 29144 8304 29150 8356
rect 29270 8304 29276 8356
rect 29328 8304 29334 8356
rect 29380 8344 29408 8375
rect 29454 8372 29460 8424
rect 29512 8412 29518 8424
rect 30193 8415 30251 8421
rect 30193 8412 30205 8415
rect 29512 8384 30205 8412
rect 29512 8372 29518 8384
rect 30193 8381 30205 8384
rect 30239 8381 30251 8415
rect 30193 8375 30251 8381
rect 31570 8372 31576 8424
rect 31628 8372 31634 8424
rect 33965 8415 34023 8421
rect 33965 8381 33977 8415
rect 34011 8412 34023 8415
rect 34011 8384 34468 8412
rect 34011 8381 34023 8384
rect 33965 8375 34023 8381
rect 34440 8356 34468 8384
rect 29822 8344 29828 8356
rect 29380 8316 29828 8344
rect 29380 8276 29408 8316
rect 29822 8304 29828 8316
rect 29880 8344 29886 8356
rect 29917 8347 29975 8353
rect 29917 8344 29929 8347
rect 29880 8316 29929 8344
rect 29880 8304 29886 8316
rect 29917 8313 29929 8316
rect 29963 8313 29975 8347
rect 29917 8307 29975 8313
rect 31864 8316 31970 8344
rect 31864 8288 31892 8316
rect 34422 8304 34428 8356
rect 34480 8304 34486 8356
rect 28368 8248 29408 8276
rect 31846 8236 31852 8288
rect 31904 8236 31910 8288
rect 2760 8186 34316 8208
rect 2760 8134 7210 8186
rect 7262 8134 7274 8186
rect 7326 8134 7338 8186
rect 7390 8134 7402 8186
rect 7454 8134 7466 8186
rect 7518 8134 15099 8186
rect 15151 8134 15163 8186
rect 15215 8134 15227 8186
rect 15279 8134 15291 8186
rect 15343 8134 15355 8186
rect 15407 8134 22988 8186
rect 23040 8134 23052 8186
rect 23104 8134 23116 8186
rect 23168 8134 23180 8186
rect 23232 8134 23244 8186
rect 23296 8134 30877 8186
rect 30929 8134 30941 8186
rect 30993 8134 31005 8186
rect 31057 8134 31069 8186
rect 31121 8134 31133 8186
rect 31185 8134 34316 8186
rect 2760 8112 34316 8134
rect 3234 8032 3240 8084
rect 3292 8032 3298 8084
rect 3789 8075 3847 8081
rect 3789 8041 3801 8075
rect 3835 8072 3847 8075
rect 4154 8072 4160 8084
rect 3835 8044 4160 8072
rect 3835 8041 3847 8044
rect 3789 8035 3847 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4246 8032 4252 8084
rect 4304 8032 4310 8084
rect 5721 8075 5779 8081
rect 5721 8041 5733 8075
rect 5767 8072 5779 8075
rect 5810 8072 5816 8084
rect 5767 8044 5816 8072
rect 5767 8041 5779 8044
rect 5721 8035 5779 8041
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 6328 8044 6469 8072
rect 6328 8032 6334 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 8113 8075 8171 8081
rect 8113 8072 8125 8075
rect 7708 8044 8125 8072
rect 7708 8032 7714 8044
rect 8113 8041 8125 8044
rect 8159 8041 8171 8075
rect 8113 8035 8171 8041
rect 8478 8032 8484 8084
rect 8536 8032 8542 8084
rect 8573 8075 8631 8081
rect 8573 8041 8585 8075
rect 8619 8072 8631 8075
rect 9214 8072 9220 8084
rect 8619 8044 9220 8072
rect 8619 8041 8631 8044
rect 8573 8035 8631 8041
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 9732 8044 10609 8072
rect 9732 8032 9738 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 11974 8072 11980 8084
rect 11756 8044 11980 8072
rect 11756 8032 11762 8044
rect 11974 8032 11980 8044
rect 12032 8072 12038 8084
rect 12434 8072 12440 8084
rect 12032 8044 12440 8072
rect 12032 8032 12038 8044
rect 12434 8032 12440 8044
rect 12492 8032 12498 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 14277 8075 14335 8081
rect 14277 8072 14289 8075
rect 12584 8044 14289 8072
rect 12584 8032 12590 8044
rect 14277 8041 14289 8044
rect 14323 8041 14335 8075
rect 14277 8035 14335 8041
rect 14645 8075 14703 8081
rect 14645 8041 14657 8075
rect 14691 8072 14703 8075
rect 14918 8072 14924 8084
rect 14691 8044 14924 8072
rect 14691 8041 14703 8044
rect 14645 8035 14703 8041
rect 4264 8004 4292 8032
rect 7469 8007 7527 8013
rect 7469 8004 7481 8007
rect 4172 7976 4292 8004
rect 6104 7976 7481 8004
rect 1302 7896 1308 7948
rect 1360 7936 1366 7948
rect 4172 7945 4200 7976
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 1360 7908 3065 7936
rect 1360 7896 1366 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3053 7899 3111 7905
rect 4157 7939 4215 7945
rect 4157 7905 4169 7939
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 4249 7939 4307 7945
rect 4249 7905 4261 7939
rect 4295 7936 4307 7939
rect 4617 7939 4675 7945
rect 4617 7936 4629 7939
rect 4295 7908 4629 7936
rect 4295 7905 4307 7908
rect 4249 7899 4307 7905
rect 4617 7905 4629 7908
rect 4663 7905 4675 7939
rect 4617 7899 4675 7905
rect 5629 7939 5687 7945
rect 5629 7905 5641 7939
rect 5675 7905 5687 7939
rect 5629 7899 5687 7905
rect 3697 7871 3755 7877
rect 3697 7837 3709 7871
rect 3743 7868 3755 7871
rect 4062 7868 4068 7880
rect 3743 7840 4068 7868
rect 3743 7837 3755 7840
rect 3697 7831 3755 7837
rect 4062 7828 4068 7840
rect 4120 7868 4126 7880
rect 4341 7871 4399 7877
rect 4341 7868 4353 7871
rect 4120 7840 4353 7868
rect 4120 7828 4126 7840
rect 4341 7837 4353 7840
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 4798 7868 4804 7880
rect 4488 7840 4804 7868
rect 4488 7828 4494 7840
rect 4798 7828 4804 7840
rect 4856 7868 4862 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4856 7840 5181 7868
rect 4856 7828 4862 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5644 7868 5672 7899
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6104 7945 6132 7976
rect 7469 7973 7481 7976
rect 7515 8004 7527 8007
rect 14182 8004 14188 8016
rect 7515 7976 14188 8004
rect 7515 7973 7527 7976
rect 7469 7967 7527 7973
rect 14182 7964 14188 7976
rect 14240 7964 14246 8016
rect 14292 8004 14320 8035
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 15746 8072 15752 8084
rect 15396 8044 15752 8072
rect 15286 8004 15292 8016
rect 14292 7976 15292 8004
rect 5905 7939 5963 7945
rect 5905 7936 5917 7939
rect 5776 7908 5917 7936
rect 5776 7896 5782 7908
rect 5905 7905 5917 7908
rect 5951 7905 5963 7939
rect 5905 7899 5963 7905
rect 6089 7939 6147 7945
rect 6089 7905 6101 7939
rect 6135 7905 6147 7939
rect 6089 7899 6147 7905
rect 6270 7896 6276 7948
rect 6328 7896 6334 7948
rect 6365 7939 6423 7945
rect 6365 7905 6377 7939
rect 6411 7905 6423 7939
rect 6365 7899 6423 7905
rect 6380 7868 6408 7899
rect 6454 7896 6460 7948
rect 6512 7936 6518 7948
rect 7009 7939 7067 7945
rect 7009 7936 7021 7939
rect 6512 7908 7021 7936
rect 6512 7896 6518 7908
rect 7009 7905 7021 7908
rect 7055 7905 7067 7939
rect 7009 7899 7067 7905
rect 8662 7896 8668 7948
rect 8720 7936 8726 7948
rect 8720 7908 8800 7936
rect 8720 7896 8726 7908
rect 8772 7877 8800 7908
rect 8846 7896 8852 7948
rect 8904 7936 8910 7948
rect 9033 7939 9091 7945
rect 9033 7936 9045 7939
rect 8904 7908 9045 7936
rect 8904 7896 8910 7908
rect 9033 7905 9045 7908
rect 9079 7905 9091 7939
rect 9033 7899 9091 7905
rect 5408 7840 6408 7868
rect 5408 7828 5414 7840
rect 6380 7800 6408 7840
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7837 8815 7871
rect 9048 7868 9076 7899
rect 9214 7896 9220 7948
rect 9272 7896 9278 7948
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7936 9827 7939
rect 10042 7936 10048 7948
rect 9815 7908 10048 7936
rect 9815 7905 9827 7908
rect 9769 7899 9827 7905
rect 10042 7896 10048 7908
rect 10100 7896 10106 7948
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10502 7936 10508 7948
rect 10183 7908 10508 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10502 7896 10508 7908
rect 10560 7896 10566 7948
rect 10689 7939 10747 7945
rect 10689 7905 10701 7939
rect 10735 7936 10747 7939
rect 10778 7936 10784 7948
rect 10735 7908 10784 7936
rect 10735 7905 10747 7908
rect 10689 7899 10747 7905
rect 10778 7896 10784 7908
rect 10836 7896 10842 7948
rect 11606 7896 11612 7948
rect 11664 7896 11670 7948
rect 11790 7896 11796 7948
rect 11848 7896 11854 7948
rect 11882 7896 11888 7948
rect 11940 7896 11946 7948
rect 11974 7896 11980 7948
rect 12032 7896 12038 7948
rect 14476 7945 14504 7976
rect 15286 7964 15292 7976
rect 15344 8004 15350 8016
rect 15396 8004 15424 8044
rect 15746 8032 15752 8044
rect 15804 8032 15810 8084
rect 16485 8075 16543 8081
rect 16485 8041 16497 8075
rect 16531 8072 16543 8075
rect 16758 8072 16764 8084
rect 16531 8044 16764 8072
rect 16531 8041 16543 8044
rect 16485 8035 16543 8041
rect 16758 8032 16764 8044
rect 16816 8032 16822 8084
rect 17126 8032 17132 8084
rect 17184 8032 17190 8084
rect 17405 8075 17463 8081
rect 17405 8041 17417 8075
rect 17451 8072 17463 8075
rect 17954 8072 17960 8084
rect 17451 8044 17960 8072
rect 17451 8041 17463 8044
rect 17405 8035 17463 8041
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18138 8032 18144 8084
rect 18196 8032 18202 8084
rect 19978 8072 19984 8084
rect 18800 8044 19984 8072
rect 15344 7976 15424 8004
rect 15344 7964 15350 7976
rect 14461 7939 14519 7945
rect 12636 7908 14320 7936
rect 9493 7871 9551 7877
rect 9493 7868 9505 7871
rect 9048 7840 9505 7868
rect 8757 7831 8815 7837
rect 9493 7837 9505 7840
rect 9539 7868 9551 7871
rect 9674 7868 9680 7880
rect 9539 7840 9680 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 9907 7840 10180 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 8202 7800 8208 7812
rect 6380 7772 8208 7800
rect 8202 7760 8208 7772
rect 8260 7760 8266 7812
rect 9306 7760 9312 7812
rect 9364 7800 9370 7812
rect 9876 7800 9904 7831
rect 9364 7772 9904 7800
rect 10152 7800 10180 7840
rect 10226 7828 10232 7880
rect 10284 7868 10290 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 10284 7840 11437 7868
rect 10284 7828 10290 7840
rect 11425 7837 11437 7840
rect 11471 7868 11483 7871
rect 12636 7868 12664 7908
rect 14292 7880 14320 7908
rect 14461 7905 14473 7939
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 11471 7840 12664 7868
rect 12989 7871 13047 7877
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 12989 7837 13001 7871
rect 13035 7868 13047 7871
rect 13035 7840 13584 7868
rect 13035 7837 13047 7840
rect 12989 7831 13047 7837
rect 10152 7772 11100 7800
rect 9364 7760 9370 7772
rect 6086 7692 6092 7744
rect 6144 7692 6150 7744
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 9950 7732 9956 7744
rect 8628 7704 9956 7732
rect 8628 7692 8634 7704
rect 9950 7692 9956 7704
rect 10008 7692 10014 7744
rect 10410 7692 10416 7744
rect 10468 7692 10474 7744
rect 11072 7741 11100 7772
rect 11882 7760 11888 7812
rect 11940 7800 11946 7812
rect 13556 7800 13584 7840
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13688 7840 13737 7868
rect 13688 7828 13694 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14660 7800 14688 7899
rect 14734 7896 14740 7948
rect 14792 7896 14798 7948
rect 16666 7936 16672 7948
rect 16146 7908 16672 7936
rect 16666 7896 16672 7908
rect 16724 7896 16730 7948
rect 17144 7945 17172 8032
rect 17678 7964 17684 8016
rect 17736 7964 17742 8016
rect 17770 7964 17776 8016
rect 17828 7964 17834 8016
rect 16853 7939 16911 7945
rect 16853 7905 16865 7939
rect 16899 7905 16911 7939
rect 16853 7899 16911 7905
rect 17129 7939 17187 7945
rect 17129 7905 17141 7939
rect 17175 7905 17187 7939
rect 17129 7899 17187 7905
rect 15013 7871 15071 7877
rect 15013 7837 15025 7871
rect 15059 7868 15071 7871
rect 15746 7868 15752 7880
rect 15059 7840 15752 7868
rect 15059 7837 15071 7840
rect 15013 7831 15071 7837
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 16868 7868 16896 7899
rect 17218 7868 17224 7880
rect 16868 7840 17224 7868
rect 17218 7828 17224 7840
rect 17276 7828 17282 7880
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 17368 7840 17417 7868
rect 17368 7828 17374 7840
rect 17405 7837 17417 7840
rect 17451 7868 17463 7871
rect 17696 7868 17724 7964
rect 18325 7939 18383 7945
rect 18325 7905 18337 7939
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 17451 7840 17724 7868
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 18340 7800 18368 7899
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 18800 7945 18828 8044
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 21560 8044 22784 8072
rect 19242 7964 19248 8016
rect 19300 7964 19306 8016
rect 19889 8007 19947 8013
rect 19889 7973 19901 8007
rect 19935 8004 19947 8007
rect 21450 8004 21456 8016
rect 19935 7976 21456 8004
rect 19935 7973 19947 7976
rect 19889 7967 19947 7973
rect 21450 7964 21456 7976
rect 21508 8004 21514 8016
rect 21560 8004 21588 8044
rect 21508 7976 21588 8004
rect 21508 7964 21514 7976
rect 21634 7964 21640 8016
rect 21692 8004 21698 8016
rect 21913 8007 21971 8013
rect 21913 8004 21925 8007
rect 21692 7976 21925 8004
rect 21692 7964 21698 7976
rect 21913 7973 21925 7976
rect 21959 7973 21971 8007
rect 21913 7967 21971 7973
rect 18785 7939 18843 7945
rect 18785 7936 18797 7939
rect 18748 7908 18797 7936
rect 18748 7896 18754 7908
rect 18785 7905 18797 7908
rect 18831 7905 18843 7939
rect 18785 7899 18843 7905
rect 19061 7939 19119 7945
rect 19061 7905 19073 7939
rect 19107 7905 19119 7939
rect 19061 7899 19119 7905
rect 11940 7772 13216 7800
rect 13556 7772 14688 7800
rect 11940 7760 11946 7772
rect 11057 7735 11115 7741
rect 11057 7701 11069 7735
rect 11103 7732 11115 7735
rect 11606 7732 11612 7744
rect 11103 7704 11612 7732
rect 11103 7701 11115 7704
rect 11057 7695 11115 7701
rect 11606 7692 11612 7704
rect 11664 7692 11670 7744
rect 12158 7692 12164 7744
rect 12216 7692 12222 7744
rect 13188 7741 13216 7772
rect 13173 7735 13231 7741
rect 13173 7701 13185 7735
rect 13219 7732 13231 7735
rect 13998 7732 14004 7744
rect 13219 7704 14004 7732
rect 13219 7701 13231 7704
rect 13173 7695 13231 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 14660 7732 14688 7772
rect 16776 7772 18368 7800
rect 16776 7744 16804 7772
rect 18598 7760 18604 7812
rect 18656 7800 18662 7812
rect 18785 7803 18843 7809
rect 18785 7800 18797 7803
rect 18656 7772 18797 7800
rect 18656 7760 18662 7772
rect 18785 7769 18797 7772
rect 18831 7769 18843 7803
rect 19076 7800 19104 7899
rect 19150 7896 19156 7948
rect 19208 7896 19214 7948
rect 19260 7936 19288 7964
rect 22756 7948 22784 8044
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 23109 8075 23167 8081
rect 23109 8072 23121 8075
rect 22888 8044 23121 8072
rect 22888 8032 22894 8044
rect 23109 8041 23121 8044
rect 23155 8072 23167 8075
rect 23382 8072 23388 8084
rect 23155 8044 23388 8072
rect 23155 8041 23167 8044
rect 23109 8035 23167 8041
rect 23382 8032 23388 8044
rect 23440 8032 23446 8084
rect 24302 8072 24308 8084
rect 24136 8044 24308 8072
rect 24136 8013 24164 8044
rect 24302 8032 24308 8044
rect 24360 8032 24366 8084
rect 24946 8032 24952 8084
rect 25004 8072 25010 8084
rect 25685 8075 25743 8081
rect 25685 8072 25697 8075
rect 25004 8044 25697 8072
rect 25004 8032 25010 8044
rect 25685 8041 25697 8044
rect 25731 8041 25743 8075
rect 25685 8035 25743 8041
rect 26418 8032 26424 8084
rect 26476 8072 26482 8084
rect 27065 8075 27123 8081
rect 27065 8072 27077 8075
rect 26476 8044 27077 8072
rect 26476 8032 26482 8044
rect 27065 8041 27077 8044
rect 27111 8041 27123 8075
rect 27065 8035 27123 8041
rect 27890 8032 27896 8084
rect 27948 8072 27954 8084
rect 28077 8075 28135 8081
rect 28077 8072 28089 8075
rect 27948 8044 28089 8072
rect 27948 8032 27954 8044
rect 28077 8041 28089 8044
rect 28123 8041 28135 8075
rect 28077 8035 28135 8041
rect 29086 8032 29092 8084
rect 29144 8072 29150 8084
rect 30190 8072 30196 8084
rect 29144 8044 30196 8072
rect 29144 8032 29150 8044
rect 30190 8032 30196 8044
rect 30248 8072 30254 8084
rect 31205 8075 31263 8081
rect 31205 8072 31217 8075
rect 30248 8044 31217 8072
rect 30248 8032 30254 8044
rect 31205 8041 31217 8044
rect 31251 8041 31263 8075
rect 31205 8035 31263 8041
rect 32033 8075 32091 8081
rect 32033 8041 32045 8075
rect 32079 8072 32091 8075
rect 32582 8072 32588 8084
rect 32079 8044 32588 8072
rect 32079 8041 32091 8044
rect 32033 8035 32091 8041
rect 32582 8032 32588 8044
rect 32640 8032 32646 8084
rect 24121 8007 24179 8013
rect 24121 7973 24133 8007
rect 24167 7973 24179 8007
rect 25406 8004 25412 8016
rect 25346 7976 25412 8004
rect 24121 7967 24179 7973
rect 25406 7964 25412 7976
rect 25464 7964 25470 8016
rect 28810 7964 28816 8016
rect 28868 8004 28874 8016
rect 32401 8007 32459 8013
rect 32401 8004 32413 8007
rect 28868 7976 29394 8004
rect 30208 7976 32413 8004
rect 28868 7964 28874 7976
rect 19429 7939 19487 7945
rect 19429 7936 19441 7939
rect 19260 7908 19441 7936
rect 19429 7905 19441 7908
rect 19475 7905 19487 7939
rect 19429 7899 19487 7905
rect 21726 7896 21732 7948
rect 21784 7936 21790 7948
rect 22646 7936 22652 7948
rect 21784 7908 22652 7936
rect 21784 7896 21790 7908
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 22738 7896 22744 7948
rect 22796 7896 22802 7948
rect 25498 7896 25504 7948
rect 25556 7936 25562 7948
rect 27157 7939 27215 7945
rect 27157 7936 27169 7939
rect 25556 7908 27169 7936
rect 25556 7896 25562 7908
rect 27157 7905 27169 7908
rect 27203 7905 27215 7939
rect 27157 7899 27215 7905
rect 19702 7800 19708 7812
rect 19076 7772 19708 7800
rect 18785 7763 18843 7769
rect 19702 7760 19708 7772
rect 19760 7760 19766 7812
rect 21744 7800 21772 7896
rect 23566 7868 23572 7880
rect 22066 7840 23572 7868
rect 22066 7800 22094 7840
rect 23566 7828 23572 7840
rect 23624 7828 23630 7880
rect 23842 7828 23848 7880
rect 23900 7868 23906 7880
rect 24762 7868 24768 7880
rect 23900 7840 24768 7868
rect 23900 7828 23906 7840
rect 24762 7828 24768 7840
rect 24820 7828 24826 7880
rect 25593 7871 25651 7877
rect 25593 7837 25605 7871
rect 25639 7868 25651 7871
rect 26237 7871 26295 7877
rect 26237 7868 26249 7871
rect 25639 7840 26249 7868
rect 25639 7837 25651 7840
rect 25593 7831 25651 7837
rect 26237 7837 26249 7840
rect 26283 7837 26295 7871
rect 26237 7831 26295 7837
rect 26418 7828 26424 7880
rect 26476 7828 26482 7880
rect 27798 7828 27804 7880
rect 27856 7868 27862 7880
rect 28629 7871 28687 7877
rect 28629 7868 28641 7871
rect 27856 7840 28641 7868
rect 27856 7828 27862 7840
rect 28629 7837 28641 7840
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 28902 7828 28908 7880
rect 28960 7828 28966 7880
rect 30208 7868 30236 7976
rect 32401 7973 32413 7976
rect 32447 7973 32459 8007
rect 32401 7967 32459 7973
rect 30558 7896 30564 7948
rect 30616 7936 30622 7948
rect 32582 7936 32588 7948
rect 30616 7908 32588 7936
rect 30616 7896 30622 7908
rect 32582 7896 32588 7908
rect 32640 7936 32646 7948
rect 32861 7939 32919 7945
rect 32861 7936 32873 7939
rect 32640 7908 32873 7936
rect 32640 7896 32646 7908
rect 32861 7905 32873 7908
rect 32907 7905 32919 7939
rect 32861 7899 32919 7905
rect 33410 7896 33416 7948
rect 33468 7896 33474 7948
rect 29932 7840 30236 7868
rect 19812 7772 21772 7800
rect 21836 7772 22094 7800
rect 22296 7772 23980 7800
rect 15194 7732 15200 7744
rect 14660 7704 15200 7732
rect 15194 7692 15200 7704
rect 15252 7692 15258 7744
rect 16758 7692 16764 7744
rect 16816 7692 16822 7744
rect 16945 7735 17003 7741
rect 16945 7701 16957 7735
rect 16991 7732 17003 7735
rect 17221 7735 17279 7741
rect 17221 7732 17233 7735
rect 16991 7704 17233 7732
rect 16991 7701 17003 7704
rect 16945 7695 17003 7701
rect 17221 7701 17233 7704
rect 17267 7701 17279 7735
rect 17221 7695 17279 7701
rect 18414 7692 18420 7744
rect 18472 7692 18478 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19521 7735 19579 7741
rect 19521 7732 19533 7735
rect 19392 7704 19533 7732
rect 19392 7692 19398 7704
rect 19521 7701 19533 7704
rect 19567 7732 19579 7735
rect 19812 7732 19840 7772
rect 19567 7704 19840 7732
rect 19567 7701 19579 7704
rect 19521 7695 19579 7701
rect 21174 7692 21180 7744
rect 21232 7692 21238 7744
rect 21542 7692 21548 7744
rect 21600 7732 21606 7744
rect 21836 7732 21864 7772
rect 21600 7704 21864 7732
rect 21600 7692 21606 7704
rect 22002 7692 22008 7744
rect 22060 7732 22066 7744
rect 22296 7732 22324 7772
rect 22060 7704 22324 7732
rect 22373 7735 22431 7741
rect 22060 7692 22066 7704
rect 22373 7701 22385 7735
rect 22419 7732 22431 7735
rect 22646 7732 22652 7744
rect 22419 7704 22652 7732
rect 22419 7701 22431 7704
rect 22373 7695 22431 7701
rect 22646 7692 22652 7704
rect 22704 7692 22710 7744
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 23750 7732 23756 7744
rect 22796 7704 23756 7732
rect 22796 7692 22802 7704
rect 23750 7692 23756 7704
rect 23808 7692 23814 7744
rect 23952 7732 23980 7772
rect 27801 7735 27859 7741
rect 27801 7732 27813 7735
rect 23952 7704 27813 7732
rect 27801 7701 27813 7704
rect 27847 7732 27859 7735
rect 29932 7732 29960 7840
rect 30742 7828 30748 7880
rect 30800 7868 30806 7880
rect 31021 7871 31079 7877
rect 31021 7868 31033 7871
rect 30800 7840 31033 7868
rect 30800 7828 30806 7840
rect 31021 7837 31033 7840
rect 31067 7837 31079 7871
rect 31021 7831 31079 7837
rect 31757 7871 31815 7877
rect 31757 7837 31769 7871
rect 31803 7837 31815 7871
rect 31757 7831 31815 7837
rect 30377 7803 30435 7809
rect 30377 7769 30389 7803
rect 30423 7800 30435 7803
rect 31772 7800 31800 7831
rect 32306 7828 32312 7880
rect 32364 7868 32370 7880
rect 32493 7871 32551 7877
rect 32493 7868 32505 7871
rect 32364 7840 32505 7868
rect 32364 7828 32370 7840
rect 32493 7837 32505 7840
rect 32539 7837 32551 7871
rect 32493 7831 32551 7837
rect 32674 7828 32680 7880
rect 32732 7868 32738 7880
rect 33502 7868 33508 7880
rect 32732 7840 33508 7868
rect 32732 7828 32738 7840
rect 33502 7828 33508 7840
rect 33560 7828 33566 7880
rect 30423 7772 31800 7800
rect 30423 7769 30435 7772
rect 30377 7763 30435 7769
rect 27847 7704 29960 7732
rect 27847 7701 27859 7704
rect 27801 7695 27859 7701
rect 30006 7692 30012 7744
rect 30064 7732 30070 7744
rect 30469 7735 30527 7741
rect 30469 7732 30481 7735
rect 30064 7704 30481 7732
rect 30064 7692 30070 7704
rect 30469 7701 30481 7704
rect 30515 7701 30527 7735
rect 30469 7695 30527 7701
rect 2760 7642 34316 7664
rect 2760 7590 6550 7642
rect 6602 7590 6614 7642
rect 6666 7590 6678 7642
rect 6730 7590 6742 7642
rect 6794 7590 6806 7642
rect 6858 7590 14439 7642
rect 14491 7590 14503 7642
rect 14555 7590 14567 7642
rect 14619 7590 14631 7642
rect 14683 7590 14695 7642
rect 14747 7590 22328 7642
rect 22380 7590 22392 7642
rect 22444 7590 22456 7642
rect 22508 7590 22520 7642
rect 22572 7590 22584 7642
rect 22636 7590 30217 7642
rect 30269 7590 30281 7642
rect 30333 7590 30345 7642
rect 30397 7590 30409 7642
rect 30461 7590 30473 7642
rect 30525 7590 34316 7642
rect 2760 7568 34316 7590
rect 7469 7531 7527 7537
rect 7469 7528 7481 7531
rect 6012 7500 7481 7528
rect 3510 7352 3516 7404
rect 3568 7352 3574 7404
rect 6012 7392 6040 7500
rect 7469 7497 7481 7500
rect 7515 7528 7527 7531
rect 9030 7528 9036 7540
rect 7515 7500 9036 7528
rect 7515 7497 7527 7500
rect 7469 7491 7527 7497
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 10134 7488 10140 7540
rect 10192 7528 10198 7540
rect 10594 7528 10600 7540
rect 10192 7500 10600 7528
rect 10192 7488 10198 7500
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 12158 7537 12164 7540
rect 12148 7531 12164 7537
rect 12148 7497 12160 7531
rect 12148 7491 12164 7497
rect 12158 7488 12164 7491
rect 12216 7488 12222 7540
rect 13630 7488 13636 7540
rect 13688 7488 13694 7540
rect 14090 7488 14096 7540
rect 14148 7488 14154 7540
rect 15289 7531 15347 7537
rect 15289 7497 15301 7531
rect 15335 7528 15347 7531
rect 15470 7528 15476 7540
rect 15335 7500 15476 7528
rect 15335 7497 15347 7500
rect 15289 7491 15347 7497
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 15746 7488 15752 7540
rect 15804 7488 15810 7540
rect 16666 7488 16672 7540
rect 16724 7488 16730 7540
rect 17310 7528 17316 7540
rect 16868 7500 17316 7528
rect 6086 7420 6092 7472
rect 6144 7460 6150 7472
rect 6144 7432 9444 7460
rect 6144 7420 6150 7432
rect 6012 7364 6224 7392
rect 6196 7336 6224 7364
rect 3142 7284 3148 7336
rect 3200 7284 3206 7336
rect 5261 7327 5319 7333
rect 5261 7293 5273 7327
rect 5307 7324 5319 7327
rect 5442 7324 5448 7336
rect 5307 7296 5448 7324
rect 5307 7293 5319 7296
rect 5261 7287 5319 7293
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 6086 7284 6092 7336
rect 6144 7284 6150 7336
rect 6178 7284 6184 7336
rect 6236 7284 6242 7336
rect 6380 7333 6408 7432
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6512 7364 7021 7392
rect 6512 7352 6518 7364
rect 6564 7333 6592 7364
rect 7009 7361 7021 7364
rect 7055 7392 7067 7395
rect 9306 7392 9312 7404
rect 7055 7364 9312 7392
rect 7055 7361 7067 7364
rect 7009 7355 7067 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 6549 7327 6607 7333
rect 6549 7293 6561 7327
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8665 7327 8723 7333
rect 8665 7324 8677 7327
rect 8352 7296 8677 7324
rect 8352 7284 8358 7296
rect 8665 7293 8677 7296
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 6457 7259 6515 7265
rect 6457 7225 6469 7259
rect 6503 7225 6515 7259
rect 9416 7256 9444 7432
rect 10410 7420 10416 7472
rect 10468 7420 10474 7472
rect 10428 7392 10456 7420
rect 11149 7395 11207 7401
rect 11149 7392 11161 7395
rect 10428 7364 11161 7392
rect 11149 7361 11161 7364
rect 11195 7361 11207 7395
rect 11149 7355 11207 7361
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7392 11943 7395
rect 12250 7392 12256 7404
rect 11931 7364 12256 7392
rect 11931 7361 11943 7364
rect 11885 7355 11943 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 14108 7392 14136 7488
rect 14826 7460 14832 7472
rect 14660 7432 14832 7460
rect 14660 7392 14688 7432
rect 14826 7420 14832 7432
rect 14884 7460 14890 7472
rect 14884 7432 16344 7460
rect 14884 7420 14890 7432
rect 14108 7364 14688 7392
rect 10778 7284 10784 7336
rect 10836 7324 10842 7336
rect 11333 7327 11391 7333
rect 11333 7324 11345 7327
rect 10836 7296 11345 7324
rect 10836 7284 10842 7296
rect 11333 7293 11345 7296
rect 11379 7293 11391 7327
rect 11333 7287 11391 7293
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14660 7333 14688 7364
rect 15562 7352 15568 7404
rect 15620 7392 15626 7404
rect 16209 7395 16267 7401
rect 16209 7392 16221 7395
rect 15620 7364 16221 7392
rect 15620 7352 15626 7364
rect 16209 7361 16221 7364
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 14277 7327 14335 7333
rect 14277 7324 14289 7327
rect 13872 7296 14289 7324
rect 13872 7284 13878 7296
rect 14277 7293 14289 7296
rect 14323 7293 14335 7327
rect 14277 7287 14335 7293
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7324 14979 7327
rect 15286 7324 15292 7336
rect 14967 7296 15292 7324
rect 14967 7293 14979 7296
rect 14921 7287 14979 7293
rect 15286 7284 15292 7296
rect 15344 7324 15350 7336
rect 15470 7324 15476 7336
rect 15344 7296 15476 7324
rect 15344 7284 15350 7296
rect 15470 7284 15476 7296
rect 15528 7284 15534 7336
rect 15930 7284 15936 7336
rect 15988 7324 15994 7336
rect 16117 7327 16175 7333
rect 16117 7324 16129 7327
rect 15988 7296 16129 7324
rect 15988 7284 15994 7296
rect 16117 7293 16129 7296
rect 16163 7293 16175 7327
rect 16316 7324 16344 7432
rect 16393 7395 16451 7401
rect 16393 7361 16405 7395
rect 16439 7392 16451 7395
rect 16868 7392 16896 7500
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 18782 7488 18788 7540
rect 18840 7488 18846 7540
rect 19702 7488 19708 7540
rect 19760 7488 19766 7540
rect 22002 7488 22008 7540
rect 22060 7488 22066 7540
rect 23382 7528 23388 7540
rect 22204 7500 23388 7528
rect 16439 7364 16896 7392
rect 17313 7395 17371 7401
rect 16439 7361 16451 7364
rect 16393 7355 16451 7361
rect 17313 7361 17325 7395
rect 17359 7392 17371 7395
rect 17402 7392 17408 7404
rect 17359 7364 17408 7392
rect 17359 7361 17371 7364
rect 17313 7355 17371 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 19720 7392 19748 7488
rect 21266 7420 21272 7472
rect 21324 7460 21330 7472
rect 21910 7460 21916 7472
rect 21324 7432 21916 7460
rect 21324 7420 21330 7432
rect 21910 7420 21916 7432
rect 21968 7420 21974 7472
rect 19797 7395 19855 7401
rect 19797 7392 19809 7395
rect 19720 7364 19809 7392
rect 19797 7361 19809 7364
rect 19843 7361 19855 7395
rect 21453 7395 21511 7401
rect 21453 7392 21465 7395
rect 19797 7355 19855 7361
rect 20272 7364 21465 7392
rect 20272 7336 20300 7364
rect 21453 7361 21465 7364
rect 21499 7361 21511 7395
rect 21453 7355 21511 7361
rect 21545 7395 21603 7401
rect 21545 7361 21557 7395
rect 21591 7392 21603 7395
rect 22020 7392 22048 7488
rect 21591 7364 22048 7392
rect 21591 7361 21603 7364
rect 21545 7355 21603 7361
rect 16758 7324 16764 7336
rect 16316 7296 16764 7324
rect 16117 7287 16175 7293
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17037 7327 17095 7333
rect 17037 7324 17049 7327
rect 17000 7296 17049 7324
rect 17000 7284 17006 7296
rect 17037 7293 17049 7296
rect 17083 7293 17095 7327
rect 17037 7287 17095 7293
rect 18414 7284 18420 7336
rect 18472 7284 18478 7336
rect 19337 7327 19395 7333
rect 19337 7293 19349 7327
rect 19383 7324 19395 7327
rect 19705 7327 19763 7333
rect 19705 7324 19717 7327
rect 19383 7296 19717 7324
rect 19383 7293 19395 7296
rect 19337 7287 19395 7293
rect 19705 7293 19717 7296
rect 19751 7324 19763 7327
rect 20254 7324 20260 7336
rect 19751 7296 20260 7324
rect 19751 7293 19763 7296
rect 19705 7287 19763 7293
rect 20254 7284 20260 7296
rect 20312 7284 20318 7336
rect 20533 7327 20591 7333
rect 20533 7324 20545 7327
rect 20364 7296 20545 7324
rect 14553 7259 14611 7265
rect 14553 7256 14565 7259
rect 9416 7228 12020 7256
rect 13386 7228 14565 7256
rect 6457 7219 6515 7225
rect 4614 7148 4620 7200
rect 4672 7148 4678 7200
rect 5258 7148 5264 7200
rect 5316 7188 5322 7200
rect 5445 7191 5503 7197
rect 5445 7188 5457 7191
rect 5316 7160 5457 7188
rect 5316 7148 5322 7160
rect 5445 7157 5457 7160
rect 5491 7188 5503 7191
rect 6472 7188 6500 7219
rect 11992 7200 12020 7228
rect 14553 7225 14565 7228
rect 14599 7225 14611 7259
rect 14553 7219 14611 7225
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7256 15163 7259
rect 15194 7256 15200 7268
rect 15151 7228 15200 7256
rect 15151 7225 15163 7228
rect 15105 7219 15163 7225
rect 15194 7216 15200 7228
rect 15252 7256 15258 7268
rect 15948 7256 15976 7284
rect 20364 7268 20392 7296
rect 20533 7293 20545 7296
rect 20579 7293 20591 7327
rect 20533 7287 20591 7293
rect 21085 7327 21143 7333
rect 21085 7293 21097 7327
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 21177 7327 21235 7333
rect 21177 7293 21189 7327
rect 21223 7324 21235 7327
rect 21266 7324 21272 7336
rect 21223 7296 21272 7324
rect 21223 7293 21235 7296
rect 21177 7287 21235 7293
rect 15252 7228 15976 7256
rect 15252 7216 15258 7228
rect 20346 7216 20352 7268
rect 20404 7216 20410 7268
rect 21100 7256 21128 7287
rect 21266 7284 21272 7296
rect 21324 7284 21330 7336
rect 21468 7324 21496 7355
rect 22204 7333 22232 7500
rect 23382 7488 23388 7500
rect 23440 7488 23446 7540
rect 24489 7531 24547 7537
rect 24489 7497 24501 7531
rect 24535 7528 24547 7531
rect 24854 7528 24860 7540
rect 24535 7500 24860 7528
rect 24535 7497 24547 7500
rect 24489 7491 24547 7497
rect 24854 7488 24860 7500
rect 24912 7488 24918 7540
rect 25406 7488 25412 7540
rect 25464 7488 25470 7540
rect 26053 7531 26111 7537
rect 26053 7497 26065 7531
rect 26099 7528 26111 7531
rect 26418 7528 26424 7540
rect 26099 7500 26424 7528
rect 26099 7497 26111 7500
rect 26053 7491 26111 7497
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 28169 7531 28227 7537
rect 28169 7497 28181 7531
rect 28215 7528 28227 7531
rect 28810 7528 28816 7540
rect 28215 7500 28816 7528
rect 28215 7497 28227 7500
rect 28169 7491 28227 7497
rect 28810 7488 28816 7500
rect 28868 7488 28874 7540
rect 28902 7488 28908 7540
rect 28960 7528 28966 7540
rect 28997 7531 29055 7537
rect 28997 7528 29009 7531
rect 28960 7500 29009 7528
rect 28960 7488 28966 7500
rect 28997 7497 29009 7500
rect 29043 7497 29055 7531
rect 28997 7491 29055 7497
rect 29536 7531 29594 7537
rect 29536 7497 29548 7531
rect 29582 7528 29594 7531
rect 30006 7528 30012 7540
rect 29582 7500 30012 7528
rect 29582 7497 29594 7500
rect 29536 7491 29594 7497
rect 30006 7488 30012 7500
rect 30064 7488 30070 7540
rect 30650 7488 30656 7540
rect 30708 7488 30714 7540
rect 31573 7531 31631 7537
rect 31573 7497 31585 7531
rect 31619 7528 31631 7531
rect 31846 7528 31852 7540
rect 31619 7500 31852 7528
rect 31619 7497 31631 7500
rect 31573 7491 31631 7497
rect 31846 7488 31852 7500
rect 31904 7488 31910 7540
rect 24118 7420 24124 7472
rect 24176 7460 24182 7472
rect 24176 7432 25084 7460
rect 24176 7420 24182 7432
rect 22557 7395 22615 7401
rect 22557 7361 22569 7395
rect 22603 7392 22615 7395
rect 23842 7392 23848 7404
rect 22603 7364 23848 7392
rect 22603 7361 22615 7364
rect 22557 7355 22615 7361
rect 23842 7352 23848 7364
rect 23900 7352 23906 7404
rect 24946 7352 24952 7404
rect 25004 7352 25010 7404
rect 25056 7401 25084 7432
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7361 25099 7395
rect 25041 7355 25099 7361
rect 27798 7352 27804 7404
rect 27856 7392 27862 7404
rect 29273 7395 29331 7401
rect 29273 7392 29285 7395
rect 27856 7364 29285 7392
rect 27856 7352 27862 7364
rect 29273 7361 29285 7364
rect 29319 7392 29331 7395
rect 30190 7392 30196 7404
rect 29319 7364 30196 7392
rect 29319 7361 29331 7364
rect 29273 7355 29331 7361
rect 30190 7352 30196 7364
rect 30248 7352 30254 7404
rect 30668 7392 30696 7488
rect 30668 7364 30788 7392
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21468 7296 21833 7324
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 21913 7327 21971 7333
rect 21913 7293 21925 7327
rect 21959 7324 21971 7327
rect 22189 7327 22247 7333
rect 21959 7296 22140 7324
rect 21959 7293 21971 7296
rect 21913 7287 21971 7293
rect 20456 7228 21128 7256
rect 5491 7160 6500 7188
rect 5491 7157 5503 7160
rect 5445 7151 5503 7157
rect 6546 7148 6552 7200
rect 6604 7188 6610 7200
rect 6733 7191 6791 7197
rect 6733 7188 6745 7191
rect 6604 7160 6745 7188
rect 6604 7148 6610 7160
rect 6733 7157 6745 7160
rect 6779 7157 6791 7191
rect 6733 7151 6791 7157
rect 8573 7191 8631 7197
rect 8573 7157 8585 7191
rect 8619 7188 8631 7191
rect 8662 7188 8668 7200
rect 8619 7160 8668 7188
rect 8619 7157 8631 7160
rect 8573 7151 8631 7157
rect 8662 7148 8668 7160
rect 8720 7188 8726 7200
rect 9030 7188 9036 7200
rect 8720 7160 9036 7188
rect 8720 7148 8726 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9674 7148 9680 7200
rect 9732 7188 9738 7200
rect 10226 7188 10232 7200
rect 9732 7160 10232 7188
rect 9732 7148 9738 7160
rect 10226 7148 10232 7160
rect 10284 7148 10290 7200
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 10560 7160 10609 7188
rect 10560 7148 10566 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 10597 7151 10655 7157
rect 11422 7148 11428 7200
rect 11480 7148 11486 7200
rect 11974 7148 11980 7200
rect 12032 7148 12038 7200
rect 13538 7148 13544 7200
rect 13596 7188 13602 7200
rect 13725 7191 13783 7197
rect 13725 7188 13737 7191
rect 13596 7160 13737 7188
rect 13596 7148 13602 7160
rect 13725 7157 13737 7160
rect 13771 7157 13783 7191
rect 13725 7151 13783 7157
rect 14274 7148 14280 7200
rect 14332 7188 14338 7200
rect 19426 7188 19432 7200
rect 14332 7160 19432 7188
rect 14332 7148 14338 7160
rect 19426 7148 19432 7160
rect 19484 7148 19490 7200
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 20456 7197 20484 7228
rect 21726 7216 21732 7268
rect 21784 7256 21790 7268
rect 22005 7259 22063 7265
rect 22005 7256 22017 7259
rect 21784 7228 22017 7256
rect 21784 7216 21790 7228
rect 22005 7225 22017 7228
rect 22051 7225 22063 7259
rect 22112 7256 22140 7296
rect 22189 7293 22201 7327
rect 22235 7293 22247 7327
rect 22189 7287 22247 7293
rect 22462 7284 22468 7336
rect 22520 7284 22526 7336
rect 25317 7327 25375 7333
rect 25317 7293 25329 7327
rect 25363 7293 25375 7327
rect 25317 7287 25375 7293
rect 28077 7327 28135 7333
rect 28077 7293 28089 7327
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 22480 7256 22508 7284
rect 22112 7228 22508 7256
rect 22833 7259 22891 7265
rect 22005 7219 22063 7225
rect 22833 7225 22845 7259
rect 22879 7225 22891 7259
rect 25130 7256 25136 7268
rect 24058 7228 25136 7256
rect 22833 7219 22891 7225
rect 20441 7191 20499 7197
rect 20441 7188 20453 7191
rect 19944 7160 20453 7188
rect 19944 7148 19950 7160
rect 20441 7157 20453 7160
rect 20487 7157 20499 7191
rect 20441 7151 20499 7157
rect 20625 7191 20683 7197
rect 20625 7157 20637 7191
rect 20671 7188 20683 7191
rect 20714 7188 20720 7200
rect 20671 7160 20720 7188
rect 20671 7157 20683 7160
rect 20625 7151 20683 7157
rect 20714 7148 20720 7160
rect 20772 7148 20778 7200
rect 20901 7191 20959 7197
rect 20901 7157 20913 7191
rect 20947 7188 20959 7191
rect 20990 7188 20996 7200
rect 20947 7160 20996 7188
rect 20947 7157 20959 7160
rect 20901 7151 20959 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21637 7191 21695 7197
rect 21637 7157 21649 7191
rect 21683 7188 21695 7191
rect 22094 7188 22100 7200
rect 21683 7160 22100 7188
rect 21683 7157 21695 7160
rect 21637 7151 21695 7157
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 22848 7188 22876 7219
rect 25130 7216 25136 7228
rect 25188 7216 25194 7268
rect 25222 7216 25228 7268
rect 25280 7256 25286 7268
rect 25332 7256 25360 7287
rect 25280 7228 25360 7256
rect 25280 7216 25286 7228
rect 26970 7216 26976 7268
rect 27028 7216 27034 7268
rect 27525 7259 27583 7265
rect 27525 7225 27537 7259
rect 27571 7256 27583 7259
rect 27614 7256 27620 7268
rect 27571 7228 27620 7256
rect 27571 7225 27583 7228
rect 27525 7219 27583 7225
rect 27614 7216 27620 7228
rect 27672 7216 27678 7268
rect 23474 7188 23480 7200
rect 22848 7160 23480 7188
rect 23474 7148 23480 7160
rect 23532 7148 23538 7200
rect 24302 7148 24308 7200
rect 24360 7148 24366 7200
rect 24854 7148 24860 7200
rect 24912 7148 24918 7200
rect 25774 7148 25780 7200
rect 25832 7148 25838 7200
rect 27430 7148 27436 7200
rect 27488 7188 27494 7200
rect 28092 7188 28120 7287
rect 28166 7284 28172 7336
rect 28224 7324 28230 7336
rect 28353 7327 28411 7333
rect 28353 7324 28365 7327
rect 28224 7296 28365 7324
rect 28224 7284 28230 7296
rect 28353 7293 28365 7296
rect 28399 7293 28411 7327
rect 30760 7324 30788 7364
rect 31202 7352 31208 7404
rect 31260 7392 31266 7404
rect 31757 7395 31815 7401
rect 31757 7392 31769 7395
rect 31260 7364 31769 7392
rect 31260 7352 31266 7364
rect 31757 7361 31769 7364
rect 31803 7361 31815 7395
rect 31757 7355 31815 7361
rect 32030 7352 32036 7404
rect 32088 7352 32094 7404
rect 31389 7327 31447 7333
rect 31389 7324 31401 7327
rect 30760 7296 31401 7324
rect 28353 7287 28411 7293
rect 31389 7293 31401 7296
rect 31435 7324 31447 7327
rect 31481 7327 31539 7333
rect 31481 7324 31493 7327
rect 31435 7296 31493 7324
rect 31435 7293 31447 7296
rect 31389 7287 31447 7293
rect 31481 7293 31493 7296
rect 31527 7293 31539 7327
rect 31481 7287 31539 7293
rect 31297 7259 31355 7265
rect 31297 7256 31309 7259
rect 30774 7228 31309 7256
rect 31297 7225 31309 7228
rect 31343 7225 31355 7259
rect 31297 7219 31355 7225
rect 32306 7216 32312 7268
rect 32364 7216 32370 7268
rect 33686 7256 33692 7268
rect 33258 7228 33692 7256
rect 33686 7216 33692 7228
rect 33744 7216 33750 7268
rect 27488 7160 28120 7188
rect 31021 7191 31079 7197
rect 27488 7148 27494 7160
rect 31021 7157 31033 7191
rect 31067 7188 31079 7191
rect 31202 7188 31208 7200
rect 31067 7160 31208 7188
rect 31067 7157 31079 7160
rect 31021 7151 31079 7157
rect 31202 7148 31208 7160
rect 31260 7148 31266 7200
rect 32324 7188 32352 7216
rect 33505 7191 33563 7197
rect 33505 7188 33517 7191
rect 32324 7160 33517 7188
rect 33505 7157 33517 7160
rect 33551 7157 33563 7191
rect 33505 7151 33563 7157
rect 2760 7098 34316 7120
rect 2760 7046 7210 7098
rect 7262 7046 7274 7098
rect 7326 7046 7338 7098
rect 7390 7046 7402 7098
rect 7454 7046 7466 7098
rect 7518 7046 15099 7098
rect 15151 7046 15163 7098
rect 15215 7046 15227 7098
rect 15279 7046 15291 7098
rect 15343 7046 15355 7098
rect 15407 7046 22988 7098
rect 23040 7046 23052 7098
rect 23104 7046 23116 7098
rect 23168 7046 23180 7098
rect 23232 7046 23244 7098
rect 23296 7046 30877 7098
rect 30929 7046 30941 7098
rect 30993 7046 31005 7098
rect 31057 7046 31069 7098
rect 31121 7046 31133 7098
rect 31185 7046 34316 7098
rect 2760 7024 34316 7046
rect 3789 6987 3847 6993
rect 3789 6953 3801 6987
rect 3835 6984 3847 6987
rect 5258 6984 5264 6996
rect 3835 6956 5264 6984
rect 3835 6953 3847 6956
rect 3789 6947 3847 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 6086 6944 6092 6996
rect 6144 6944 6150 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12894 6984 12900 6996
rect 12492 6956 12900 6984
rect 12492 6944 12498 6956
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 14182 6944 14188 6996
rect 14240 6984 14246 6996
rect 18690 6984 18696 6996
rect 14240 6956 18696 6984
rect 14240 6944 14246 6956
rect 18690 6944 18696 6956
rect 18748 6984 18754 6996
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 18748 6956 18797 6984
rect 18748 6944 18754 6956
rect 18785 6953 18797 6956
rect 18831 6953 18843 6987
rect 18785 6947 18843 6953
rect 19334 6944 19340 6996
rect 19392 6944 19398 6996
rect 20346 6944 20352 6996
rect 20404 6984 20410 6996
rect 20404 6956 22094 6984
rect 20404 6944 20410 6956
rect 3142 6876 3148 6928
rect 3200 6916 3206 6928
rect 3697 6919 3755 6925
rect 3697 6916 3709 6919
rect 3200 6888 3709 6916
rect 3200 6876 3206 6888
rect 3697 6885 3709 6888
rect 3743 6885 3755 6919
rect 3697 6879 3755 6885
rect 4525 6919 4583 6925
rect 4525 6885 4537 6919
rect 4571 6916 4583 6919
rect 4614 6916 4620 6928
rect 4571 6888 4620 6916
rect 4571 6885 4583 6888
rect 4525 6879 4583 6885
rect 4614 6876 4620 6888
rect 4672 6876 4678 6928
rect 6270 6916 6276 6928
rect 5750 6888 6276 6916
rect 6270 6876 6276 6888
rect 6328 6876 6334 6928
rect 7098 6876 7104 6928
rect 7156 6876 7162 6928
rect 15930 6876 15936 6928
rect 15988 6916 15994 6928
rect 16945 6919 17003 6925
rect 16945 6916 16957 6919
rect 15988 6888 16957 6916
rect 15988 6876 15994 6888
rect 16945 6885 16957 6888
rect 16991 6885 17003 6919
rect 16945 6879 17003 6885
rect 18141 6919 18199 6925
rect 18141 6885 18153 6919
rect 18187 6916 18199 6919
rect 19352 6916 19380 6944
rect 18187 6888 19380 6916
rect 18187 6885 18199 6888
rect 18141 6879 18199 6885
rect 20714 6876 20720 6928
rect 20772 6876 20778 6928
rect 22066 6916 22094 6956
rect 23566 6944 23572 6996
rect 23624 6984 23630 6996
rect 23624 6956 24808 6984
rect 23624 6944 23630 6956
rect 24780 6916 24808 6956
rect 24854 6944 24860 6996
rect 24912 6984 24918 6996
rect 25317 6987 25375 6993
rect 25317 6984 25329 6987
rect 24912 6956 25329 6984
rect 24912 6944 24918 6956
rect 25317 6953 25329 6956
rect 25363 6953 25375 6987
rect 25317 6947 25375 6953
rect 26510 6944 26516 6996
rect 26568 6944 26574 6996
rect 27614 6944 27620 6996
rect 27672 6984 27678 6996
rect 27709 6987 27767 6993
rect 27709 6984 27721 6987
rect 27672 6956 27721 6984
rect 27672 6944 27678 6956
rect 27709 6953 27721 6956
rect 27755 6953 27767 6987
rect 27709 6947 27767 6953
rect 30098 6944 30104 6996
rect 30156 6944 30162 6996
rect 30469 6987 30527 6993
rect 30469 6953 30481 6987
rect 30515 6984 30527 6987
rect 30742 6984 30748 6996
rect 30515 6956 30748 6984
rect 30515 6953 30527 6956
rect 30469 6947 30527 6953
rect 30742 6944 30748 6956
rect 30800 6944 30806 6996
rect 32125 6987 32183 6993
rect 32125 6984 32137 6987
rect 32083 6956 32137 6984
rect 32125 6953 32137 6956
rect 32171 6984 32183 6987
rect 32674 6984 32680 6996
rect 32171 6956 32680 6984
rect 32171 6953 32183 6956
rect 32125 6947 32183 6953
rect 25774 6916 25780 6928
rect 22066 6888 22232 6916
rect 22204 6860 22232 6888
rect 23400 6888 24348 6916
rect 24780 6888 25780 6916
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 3375 6820 4200 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3878 6780 3884 6792
rect 3651 6752 3884 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4172 6780 4200 6820
rect 4246 6808 4252 6860
rect 4304 6808 4310 6860
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6848 8355 6851
rect 8386 6848 8392 6860
rect 8343 6820 8392 6848
rect 8343 6817 8355 6820
rect 8297 6811 8355 6817
rect 8386 6808 8392 6820
rect 8444 6808 8450 6860
rect 10502 6808 10508 6860
rect 10560 6808 10566 6860
rect 11422 6848 11428 6860
rect 10626 6820 11428 6848
rect 11422 6808 11428 6820
rect 11480 6808 11486 6860
rect 13722 6808 13728 6860
rect 13780 6848 13786 6860
rect 13817 6851 13875 6857
rect 13817 6848 13829 6851
rect 13780 6820 13829 6848
rect 13780 6808 13786 6820
rect 13817 6817 13829 6820
rect 13863 6817 13875 6851
rect 13817 6811 13875 6817
rect 16025 6851 16083 6857
rect 16025 6817 16037 6851
rect 16071 6848 16083 6851
rect 16574 6848 16580 6860
rect 16071 6820 16580 6848
rect 16071 6817 16083 6820
rect 16025 6811 16083 6817
rect 16574 6808 16580 6820
rect 16632 6848 16638 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 16632 6820 17417 6848
rect 16632 6808 16638 6820
rect 17405 6817 17417 6820
rect 17451 6848 17463 6851
rect 18046 6848 18052 6860
rect 17451 6820 18052 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 20990 6808 20996 6860
rect 21048 6808 21054 6860
rect 22094 6808 22100 6860
rect 22152 6808 22158 6860
rect 22186 6808 22192 6860
rect 22244 6808 22250 6860
rect 23400 6848 23428 6888
rect 22940 6820 23428 6848
rect 23477 6851 23535 6857
rect 5258 6780 5264 6792
rect 4172 6752 5264 6780
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 7466 6740 7472 6792
rect 7524 6780 7530 6792
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 7524 6752 7573 6780
rect 7524 6740 7530 6752
rect 7561 6749 7573 6752
rect 7607 6749 7619 6783
rect 7561 6743 7619 6749
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 7892 6752 9229 6780
rect 7892 6740 7898 6752
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 10520 6780 10548 6808
rect 9539 6752 10548 6780
rect 10965 6783 11023 6789
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 10965 6749 10977 6783
rect 11011 6780 11023 6783
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 11011 6752 11069 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 11057 6743 11115 6749
rect 3234 6604 3240 6656
rect 3292 6604 3298 6656
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6644 4215 6647
rect 5258 6644 5264 6656
rect 4203 6616 5264 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 5258 6604 5264 6616
rect 5316 6604 5322 6656
rect 5994 6604 6000 6656
rect 6052 6604 6058 6656
rect 9232 6644 9260 6743
rect 12434 6740 12440 6792
rect 12492 6740 12498 6792
rect 16298 6740 16304 6792
rect 16356 6740 16362 6792
rect 16942 6740 16948 6792
rect 17000 6740 17006 6792
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18840 6752 18981 6780
rect 18840 6740 18846 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 19058 6740 19064 6792
rect 19116 6780 19122 6792
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19116 6752 19717 6780
rect 19116 6740 19122 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 19981 6783 20039 6789
rect 19981 6749 19993 6783
rect 20027 6780 20039 6783
rect 21008 6780 21036 6808
rect 20027 6752 21036 6780
rect 21453 6783 21511 6789
rect 20027 6749 20039 6752
rect 19981 6743 20039 6749
rect 21453 6749 21465 6783
rect 21499 6780 21511 6783
rect 22940 6780 22968 6820
rect 23477 6817 23489 6851
rect 23523 6848 23535 6851
rect 23750 6848 23756 6860
rect 23523 6820 23756 6848
rect 23523 6817 23535 6820
rect 23477 6811 23535 6817
rect 23750 6808 23756 6820
rect 23808 6848 23814 6860
rect 24118 6848 24124 6860
rect 23808 6820 24124 6848
rect 23808 6808 23814 6820
rect 24118 6808 24124 6820
rect 24176 6808 24182 6860
rect 24320 6848 24348 6888
rect 25774 6876 25780 6888
rect 25832 6876 25838 6928
rect 27801 6919 27859 6925
rect 27801 6916 27813 6919
rect 26620 6888 27813 6916
rect 25406 6848 25412 6860
rect 24320 6820 25412 6848
rect 25406 6808 25412 6820
rect 25464 6808 25470 6860
rect 25498 6808 25504 6860
rect 25556 6808 25562 6860
rect 26620 6857 26648 6888
rect 27801 6885 27813 6888
rect 27847 6885 27859 6919
rect 30116 6916 30144 6944
rect 30837 6919 30895 6925
rect 30837 6916 30849 6919
rect 30116 6888 30849 6916
rect 27801 6879 27859 6885
rect 30837 6885 30849 6888
rect 30883 6885 30895 6919
rect 30837 6879 30895 6885
rect 26605 6851 26663 6857
rect 26605 6817 26617 6851
rect 26651 6817 26663 6851
rect 27065 6851 27123 6857
rect 27065 6848 27077 6851
rect 26605 6811 26663 6817
rect 26988 6820 27077 6848
rect 21499 6752 22968 6780
rect 21499 6749 21511 6752
rect 21453 6743 21511 6749
rect 15105 6715 15163 6721
rect 11624 6684 12434 6712
rect 10134 6644 10140 6656
rect 9232 6616 10140 6644
rect 10134 6604 10140 6616
rect 10192 6604 10198 6656
rect 10226 6604 10232 6656
rect 10284 6644 10290 6656
rect 11624 6644 11652 6684
rect 10284 6616 11652 6644
rect 10284 6604 10290 6616
rect 11698 6604 11704 6656
rect 11756 6604 11762 6656
rect 11882 6604 11888 6656
rect 11940 6604 11946 6656
rect 12406 6644 12434 6684
rect 15105 6681 15117 6715
rect 15151 6712 15163 6715
rect 16960 6712 16988 6740
rect 15151 6684 16988 6712
rect 15151 6681 15163 6684
rect 15105 6675 15163 6681
rect 19334 6644 19340 6656
rect 12406 6616 19340 6644
rect 19334 6604 19340 6616
rect 19392 6604 19398 6656
rect 19610 6604 19616 6656
rect 19668 6604 19674 6656
rect 19720 6644 19748 6743
rect 23014 6740 23020 6792
rect 23072 6740 23078 6792
rect 25682 6740 25688 6792
rect 25740 6740 25746 6792
rect 26326 6740 26332 6792
rect 26384 6740 26390 6792
rect 26988 6721 27016 6820
rect 27065 6817 27077 6820
rect 27111 6817 27123 6851
rect 27065 6811 27123 6817
rect 27706 6808 27712 6860
rect 27764 6808 27770 6860
rect 27982 6808 27988 6860
rect 28040 6808 28046 6860
rect 28626 6808 28632 6860
rect 28684 6848 28690 6860
rect 30558 6848 30564 6860
rect 28684 6820 30564 6848
rect 28684 6808 28690 6820
rect 30558 6808 30564 6820
rect 30616 6808 30622 6860
rect 30929 6851 30987 6857
rect 30929 6817 30941 6851
rect 30975 6848 30987 6851
rect 32140 6848 32168 6947
rect 32674 6944 32680 6956
rect 32732 6944 32738 6996
rect 30975 6820 31248 6848
rect 30975 6817 30987 6820
rect 30929 6811 30987 6817
rect 27724 6780 27752 6808
rect 31220 6792 31248 6820
rect 32048 6820 32168 6848
rect 28169 6783 28227 6789
rect 28169 6780 28181 6783
rect 27724 6752 28181 6780
rect 28169 6749 28181 6752
rect 28215 6749 28227 6783
rect 28169 6743 28227 6749
rect 31113 6783 31171 6789
rect 31113 6749 31125 6783
rect 31159 6749 31171 6783
rect 31113 6743 31171 6749
rect 26973 6715 27031 6721
rect 26973 6681 26985 6715
rect 27019 6681 27031 6715
rect 26973 6675 27031 6681
rect 28442 6672 28448 6724
rect 28500 6712 28506 6724
rect 29454 6712 29460 6724
rect 28500 6684 29460 6712
rect 28500 6672 28506 6684
rect 29454 6672 29460 6684
rect 29512 6672 29518 6724
rect 21174 6644 21180 6656
rect 19720 6616 21180 6644
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 21542 6604 21548 6656
rect 21600 6604 21606 6656
rect 22462 6604 22468 6656
rect 22520 6644 22526 6656
rect 22830 6644 22836 6656
rect 22520 6616 22836 6644
rect 22520 6604 22526 6616
rect 22830 6604 22836 6616
rect 22888 6604 22894 6656
rect 24762 6604 24768 6656
rect 24820 6604 24826 6656
rect 24854 6604 24860 6656
rect 24912 6644 24918 6656
rect 25961 6647 26019 6653
rect 25961 6644 25973 6647
rect 24912 6616 25973 6644
rect 24912 6604 24918 6616
rect 25961 6613 25973 6616
rect 26007 6613 26019 6647
rect 25961 6607 26019 6613
rect 26234 6604 26240 6656
rect 26292 6644 26298 6656
rect 30006 6644 30012 6656
rect 26292 6616 30012 6644
rect 26292 6604 26298 6616
rect 30006 6604 30012 6616
rect 30064 6604 30070 6656
rect 30101 6647 30159 6653
rect 30101 6613 30113 6647
rect 30147 6644 30159 6647
rect 30190 6644 30196 6656
rect 30147 6616 30196 6644
rect 30147 6613 30159 6616
rect 30101 6607 30159 6613
rect 30190 6604 30196 6616
rect 30248 6644 30254 6656
rect 30742 6644 30748 6656
rect 30248 6616 30748 6644
rect 30248 6604 30254 6616
rect 30742 6604 30748 6616
rect 30800 6604 30806 6656
rect 31128 6644 31156 6743
rect 31202 6740 31208 6792
rect 31260 6740 31266 6792
rect 32048 6724 32076 6820
rect 32306 6808 32312 6860
rect 32364 6808 32370 6860
rect 33413 6851 33471 6857
rect 33413 6817 33425 6851
rect 33459 6848 33471 6851
rect 34698 6848 34704 6860
rect 33459 6820 34704 6848
rect 33459 6817 33471 6820
rect 33413 6811 33471 6817
rect 34698 6808 34704 6820
rect 34756 6808 34762 6860
rect 32030 6712 32036 6724
rect 31726 6684 32036 6712
rect 31478 6644 31484 6656
rect 31128 6616 31484 6644
rect 31478 6604 31484 6616
rect 31536 6644 31542 6656
rect 31726 6644 31754 6684
rect 32030 6672 32036 6684
rect 32088 6672 32094 6724
rect 31536 6616 31754 6644
rect 31536 6604 31542 6616
rect 2760 6554 34316 6576
rect 2760 6502 6550 6554
rect 6602 6502 6614 6554
rect 6666 6502 6678 6554
rect 6730 6502 6742 6554
rect 6794 6502 6806 6554
rect 6858 6502 14439 6554
rect 14491 6502 14503 6554
rect 14555 6502 14567 6554
rect 14619 6502 14631 6554
rect 14683 6502 14695 6554
rect 14747 6502 22328 6554
rect 22380 6502 22392 6554
rect 22444 6502 22456 6554
rect 22508 6502 22520 6554
rect 22572 6502 22584 6554
rect 22636 6502 30217 6554
rect 30269 6502 30281 6554
rect 30333 6502 30345 6554
rect 30397 6502 30409 6554
rect 30461 6502 30473 6554
rect 30525 6502 34316 6554
rect 2760 6480 34316 6502
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4246 6440 4252 6452
rect 4019 6412 4252 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 5721 6443 5779 6449
rect 5721 6409 5733 6443
rect 5767 6440 5779 6443
rect 8294 6440 8300 6452
rect 5767 6412 8300 6440
rect 5767 6409 5779 6412
rect 5721 6403 5779 6409
rect 3050 6196 3056 6248
rect 3108 6196 3114 6248
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5736 6236 5764 6403
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 12345 6443 12403 6449
rect 12345 6409 12357 6443
rect 12391 6440 12403 6443
rect 12434 6440 12440 6452
rect 12391 6412 12440 6440
rect 12391 6409 12403 6412
rect 12345 6403 12403 6409
rect 12434 6400 12440 6412
rect 12492 6400 12498 6452
rect 13081 6443 13139 6449
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 13814 6440 13820 6452
rect 13127 6412 13820 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 13814 6400 13820 6412
rect 13872 6400 13878 6452
rect 15470 6400 15476 6452
rect 15528 6400 15534 6452
rect 19610 6400 19616 6452
rect 19668 6400 19674 6452
rect 21440 6443 21498 6449
rect 21440 6409 21452 6443
rect 21486 6440 21498 6443
rect 21542 6440 21548 6452
rect 21486 6412 21548 6440
rect 21486 6409 21498 6412
rect 21440 6403 21498 6409
rect 21542 6400 21548 6412
rect 21600 6400 21606 6452
rect 22925 6443 22983 6449
rect 22925 6409 22937 6443
rect 22971 6440 22983 6443
rect 23014 6440 23020 6452
rect 22971 6412 23020 6440
rect 22971 6409 22983 6412
rect 22925 6403 22983 6409
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 23474 6400 23480 6452
rect 23532 6400 23538 6452
rect 25130 6400 25136 6452
rect 25188 6400 25194 6452
rect 25314 6400 25320 6452
rect 25372 6440 25378 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 25372 6412 25513 6440
rect 25372 6400 25378 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 30006 6400 30012 6452
rect 30064 6400 30070 6452
rect 30558 6400 30564 6452
rect 30616 6440 30622 6452
rect 30837 6443 30895 6449
rect 30837 6440 30849 6443
rect 30616 6412 30849 6440
rect 30616 6400 30622 6412
rect 30837 6409 30849 6412
rect 30883 6440 30895 6443
rect 31386 6440 31392 6452
rect 30883 6412 31392 6440
rect 30883 6409 30895 6412
rect 30837 6403 30895 6409
rect 31386 6400 31392 6412
rect 31444 6400 31450 6452
rect 33686 6400 33692 6452
rect 33744 6400 33750 6452
rect 5994 6332 6000 6384
rect 6052 6332 6058 6384
rect 6454 6332 6460 6384
rect 6512 6332 6518 6384
rect 7466 6332 7472 6384
rect 7524 6332 7530 6384
rect 18785 6375 18843 6381
rect 18785 6341 18797 6375
rect 18831 6341 18843 6375
rect 19628 6372 19656 6400
rect 18785 6335 18843 6341
rect 19260 6344 19656 6372
rect 26973 6375 27031 6381
rect 5307 6208 5764 6236
rect 6012 6236 6040 6332
rect 6472 6304 6500 6332
rect 6825 6307 6883 6313
rect 6825 6304 6837 6307
rect 6472 6276 6837 6304
rect 6825 6273 6837 6276
rect 6871 6273 6883 6307
rect 6825 6267 6883 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7834 6304 7840 6316
rect 7607 6276 7840 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 10321 6307 10379 6313
rect 10321 6304 10333 6307
rect 9088 6276 10333 6304
rect 9088 6264 9094 6276
rect 10321 6273 10333 6276
rect 10367 6304 10379 6307
rect 10410 6304 10416 6316
rect 10367 6276 10416 6304
rect 10367 6273 10379 6276
rect 10321 6267 10379 6273
rect 10410 6264 10416 6276
rect 10468 6264 10474 6316
rect 10597 6307 10655 6313
rect 10597 6273 10609 6307
rect 10643 6304 10655 6307
rect 11514 6304 11520 6316
rect 10643 6276 11520 6304
rect 10643 6273 10655 6276
rect 10597 6267 10655 6273
rect 11514 6264 11520 6276
rect 11572 6304 11578 6316
rect 12250 6304 12256 6316
rect 11572 6276 12256 6304
rect 11572 6264 11578 6276
rect 12250 6264 12256 6276
rect 12308 6304 12314 6316
rect 13449 6307 13507 6313
rect 12308 6276 13216 6304
rect 12308 6264 12314 6276
rect 6457 6239 6515 6245
rect 6457 6236 6469 6239
rect 6012 6208 6469 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 6457 6205 6469 6208
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 9582 6196 9588 6248
rect 9640 6236 9646 6248
rect 9861 6239 9919 6245
rect 9861 6236 9873 6239
rect 9640 6208 9873 6236
rect 9640 6196 9646 6208
rect 9861 6205 9873 6208
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 12526 6196 12532 6248
rect 12584 6196 12590 6248
rect 12894 6196 12900 6248
rect 12952 6196 12958 6248
rect 13188 6245 13216 6276
rect 13449 6273 13461 6307
rect 13495 6304 13507 6307
rect 13538 6304 13544 6316
rect 13495 6276 13544 6304
rect 13495 6273 13507 6276
rect 13449 6267 13507 6273
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 16850 6304 16856 6316
rect 16632 6276 16856 6304
rect 16632 6264 16638 6276
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17221 6307 17279 6313
rect 17221 6273 17233 6307
rect 17267 6304 17279 6307
rect 18800 6304 18828 6335
rect 19260 6313 19288 6344
rect 26973 6341 26985 6375
rect 27019 6341 27031 6375
rect 26973 6335 27031 6341
rect 28997 6375 29055 6381
rect 28997 6341 29009 6375
rect 29043 6341 29055 6375
rect 28997 6335 29055 6341
rect 29089 6375 29147 6381
rect 29089 6341 29101 6375
rect 29135 6372 29147 6375
rect 29178 6372 29184 6384
rect 29135 6344 29184 6372
rect 29135 6341 29147 6344
rect 29089 6335 29147 6341
rect 17267 6276 18828 6304
rect 19245 6307 19303 6313
rect 17267 6273 17279 6276
rect 17221 6267 17279 6273
rect 19245 6273 19257 6307
rect 19291 6273 19303 6307
rect 19245 6267 19303 6273
rect 19337 6307 19395 6313
rect 19337 6273 19349 6307
rect 19383 6273 19395 6307
rect 19337 6267 19395 6273
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6205 13231 6239
rect 13173 6199 13231 6205
rect 7837 6171 7895 6177
rect 7837 6137 7849 6171
rect 7883 6168 7895 6171
rect 7926 6168 7932 6180
rect 7883 6140 7932 6168
rect 7883 6137 7895 6140
rect 7837 6131 7895 6137
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 9493 6171 9551 6177
rect 9493 6168 9505 6171
rect 9062 6140 9505 6168
rect 9493 6137 9505 6140
rect 9539 6137 9551 6171
rect 9493 6131 9551 6137
rect 10870 6128 10876 6180
rect 10928 6128 10934 6180
rect 12158 6168 12164 6180
rect 12098 6140 12164 6168
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 12713 6171 12771 6177
rect 12713 6168 12725 6171
rect 12406 6140 12725 6168
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 4062 6100 4068 6112
rect 3283 6072 4068 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 5902 6060 5908 6112
rect 5960 6060 5966 6112
rect 9309 6103 9367 6109
rect 9309 6069 9321 6103
rect 9355 6100 9367 6103
rect 9766 6100 9772 6112
rect 9355 6072 9772 6100
rect 9355 6069 9367 6072
rect 9309 6063 9367 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 11790 6060 11796 6112
rect 11848 6100 11854 6112
rect 12406 6100 12434 6140
rect 12713 6137 12725 6140
rect 12759 6137 12771 6171
rect 12713 6131 12771 6137
rect 12802 6128 12808 6180
rect 12860 6128 12866 6180
rect 13188 6168 13216 6199
rect 15654 6196 15660 6248
rect 15712 6236 15718 6248
rect 16025 6239 16083 6245
rect 16025 6236 16037 6239
rect 15712 6208 16037 6236
rect 15712 6196 15718 6208
rect 16025 6205 16037 6208
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16942 6196 16948 6248
rect 17000 6196 17006 6248
rect 18690 6196 18696 6248
rect 18748 6196 18754 6248
rect 18966 6196 18972 6248
rect 19024 6236 19030 6248
rect 19153 6239 19211 6245
rect 19153 6236 19165 6239
rect 19024 6208 19165 6236
rect 19024 6196 19030 6208
rect 19153 6205 19165 6208
rect 19199 6205 19211 6239
rect 19352 6236 19380 6267
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 19794 6304 19800 6316
rect 19484 6276 19800 6304
rect 19484 6264 19490 6276
rect 19794 6264 19800 6276
rect 19852 6264 19858 6316
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6304 20223 6307
rect 20254 6304 20260 6316
rect 20211 6276 20260 6304
rect 20211 6273 20223 6276
rect 20165 6267 20223 6273
rect 20254 6264 20260 6276
rect 20312 6304 20318 6316
rect 20533 6307 20591 6313
rect 20533 6304 20545 6307
rect 20312 6276 20545 6304
rect 20312 6264 20318 6276
rect 20533 6273 20545 6276
rect 20579 6273 20591 6307
rect 20533 6267 20591 6273
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 23842 6304 23848 6316
rect 21223 6276 23848 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 23842 6264 23848 6276
rect 23900 6264 23906 6316
rect 26988 6304 27016 6335
rect 27065 6307 27123 6313
rect 27065 6304 27077 6307
rect 26988 6276 27077 6304
rect 27065 6273 27077 6276
rect 27111 6273 27123 6307
rect 27065 6267 27123 6273
rect 28810 6264 28816 6316
rect 28868 6304 28874 6316
rect 29012 6304 29040 6335
rect 29178 6332 29184 6344
rect 29236 6332 29242 6384
rect 29454 6332 29460 6384
rect 29512 6372 29518 6384
rect 30377 6375 30435 6381
rect 30377 6372 30389 6375
rect 29512 6344 30389 6372
rect 29512 6332 29518 6344
rect 30377 6341 30389 6344
rect 30423 6341 30435 6375
rect 30377 6335 30435 6341
rect 32769 6375 32827 6381
rect 32769 6341 32781 6375
rect 32815 6372 32827 6375
rect 32815 6344 33456 6372
rect 32815 6341 32827 6344
rect 32769 6335 32827 6341
rect 29641 6307 29699 6313
rect 29641 6304 29653 6307
rect 28868 6276 28912 6304
rect 29012 6276 29653 6304
rect 28868 6264 28874 6276
rect 29641 6273 29653 6276
rect 29687 6273 29699 6307
rect 29641 6267 29699 6273
rect 30558 6264 30564 6316
rect 30616 6304 30622 6316
rect 31757 6307 31815 6313
rect 31757 6304 31769 6307
rect 30616 6276 31769 6304
rect 30616 6264 30622 6276
rect 31757 6273 31769 6276
rect 31803 6273 31815 6307
rect 31757 6267 31815 6273
rect 32030 6264 32036 6316
rect 32088 6304 32094 6316
rect 33428 6313 33456 6344
rect 32125 6307 32183 6313
rect 32125 6304 32137 6307
rect 32088 6276 32137 6304
rect 32088 6264 32094 6276
rect 32125 6273 32137 6276
rect 32171 6273 32183 6307
rect 32125 6267 32183 6273
rect 33413 6307 33471 6313
rect 33413 6273 33425 6307
rect 33459 6273 33471 6307
rect 33413 6267 33471 6273
rect 19153 6199 19211 6205
rect 19306 6208 19380 6236
rect 13188 6140 13400 6168
rect 13372 6112 13400 6140
rect 14182 6128 14188 6180
rect 14240 6128 14246 6180
rect 17954 6128 17960 6180
rect 18012 6128 18018 6180
rect 18708 6168 18736 6196
rect 19306 6168 19334 6208
rect 19886 6196 19892 6248
rect 19944 6196 19950 6248
rect 23201 6239 23259 6245
rect 23201 6205 23213 6239
rect 23247 6205 23259 6239
rect 23201 6199 23259 6205
rect 18708 6140 19334 6168
rect 20257 6171 20315 6177
rect 20257 6137 20269 6171
rect 20303 6168 20315 6171
rect 21726 6168 21732 6180
rect 20303 6140 21732 6168
rect 20303 6137 20315 6140
rect 20257 6131 20315 6137
rect 21726 6128 21732 6140
rect 21784 6128 21790 6180
rect 23109 6171 23167 6177
rect 23109 6168 23121 6171
rect 22678 6140 23121 6168
rect 23109 6137 23121 6140
rect 23155 6137 23167 6171
rect 23109 6131 23167 6137
rect 11848 6072 12434 6100
rect 11848 6060 11854 6072
rect 13354 6060 13360 6112
rect 13412 6060 13418 6112
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 14921 6103 14979 6109
rect 14921 6100 14933 6103
rect 14516 6072 14933 6100
rect 14516 6060 14522 6072
rect 14921 6069 14933 6072
rect 14967 6069 14979 6103
rect 14921 6063 14979 6069
rect 18693 6103 18751 6109
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 18782 6100 18788 6112
rect 18739 6072 18788 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 18782 6060 18788 6072
rect 18840 6060 18846 6112
rect 19610 6060 19616 6112
rect 19668 6060 19674 6112
rect 22186 6060 22192 6112
rect 22244 6100 22250 6112
rect 23216 6100 23244 6199
rect 23566 6196 23572 6248
rect 23624 6196 23630 6248
rect 23658 6196 23664 6248
rect 23716 6196 23722 6248
rect 23750 6196 23756 6248
rect 23808 6196 23814 6248
rect 24026 6196 24032 6248
rect 24084 6196 24090 6248
rect 24302 6196 24308 6248
rect 24360 6196 24366 6248
rect 25222 6196 25228 6248
rect 25280 6196 25286 6248
rect 26418 6196 26424 6248
rect 26476 6196 26482 6248
rect 26789 6239 26847 6245
rect 26789 6205 26801 6239
rect 26835 6236 26847 6239
rect 26878 6236 26884 6248
rect 26835 6208 26884 6236
rect 26835 6205 26847 6208
rect 26789 6199 26847 6205
rect 26878 6196 26884 6208
rect 26936 6236 26942 6248
rect 28077 6239 28135 6245
rect 28077 6236 28089 6239
rect 26936 6208 28089 6236
rect 26936 6196 26942 6208
rect 28077 6205 28089 6208
rect 28123 6236 28135 6239
rect 28442 6236 28448 6248
rect 28123 6208 28448 6236
rect 28123 6205 28135 6208
rect 28077 6199 28135 6205
rect 28442 6196 28448 6208
rect 28500 6196 28506 6248
rect 28718 6236 28724 6248
rect 28679 6208 28724 6236
rect 28718 6196 28724 6208
rect 28776 6196 28782 6248
rect 32401 6239 32459 6245
rect 32401 6205 32413 6239
rect 32447 6236 32459 6239
rect 32582 6236 32588 6248
rect 32447 6208 32588 6236
rect 32447 6205 32459 6208
rect 32401 6199 32459 6205
rect 32582 6196 32588 6208
rect 32640 6196 32646 6248
rect 33781 6239 33839 6245
rect 33781 6205 33793 6239
rect 33827 6205 33839 6239
rect 33781 6199 33839 6205
rect 23584 6168 23612 6196
rect 23845 6171 23903 6177
rect 23845 6168 23857 6171
rect 23584 6140 23857 6168
rect 23845 6137 23857 6140
rect 23891 6137 23903 6171
rect 23845 6131 23903 6137
rect 25774 6128 25780 6180
rect 25832 6168 25838 6180
rect 26605 6171 26663 6177
rect 25832 6140 26372 6168
rect 25832 6128 25838 6140
rect 23382 6100 23388 6112
rect 22244 6072 23388 6100
rect 22244 6060 22250 6072
rect 23382 6060 23388 6072
rect 23440 6060 23446 6112
rect 23658 6060 23664 6112
rect 23716 6100 23722 6112
rect 24486 6100 24492 6112
rect 23716 6072 24492 6100
rect 23716 6060 23722 6072
rect 24486 6060 24492 6072
rect 24544 6060 24550 6112
rect 24946 6060 24952 6112
rect 25004 6060 25010 6112
rect 25682 6060 25688 6112
rect 25740 6100 25746 6112
rect 26237 6103 26295 6109
rect 26237 6100 26249 6103
rect 25740 6072 26249 6100
rect 25740 6060 25746 6072
rect 26237 6069 26249 6072
rect 26283 6069 26295 6103
rect 26344 6100 26372 6140
rect 26605 6137 26617 6171
rect 26651 6137 26663 6171
rect 26605 6131 26663 6137
rect 26697 6171 26755 6177
rect 26697 6137 26709 6171
rect 26743 6137 26755 6171
rect 26697 6131 26755 6137
rect 26620 6100 26648 6131
rect 26344 6072 26648 6100
rect 26712 6100 26740 6131
rect 26970 6128 26976 6180
rect 27028 6168 27034 6180
rect 28353 6171 28411 6177
rect 27028 6140 27844 6168
rect 27028 6128 27034 6140
rect 27246 6100 27252 6112
rect 26712 6072 27252 6100
rect 26237 6063 26295 6069
rect 27246 6060 27252 6072
rect 27304 6060 27310 6112
rect 27706 6060 27712 6112
rect 27764 6060 27770 6112
rect 27816 6100 27844 6140
rect 28353 6137 28365 6171
rect 28399 6168 28411 6171
rect 30650 6168 30656 6180
rect 28399 6140 30656 6168
rect 28399 6137 28411 6140
rect 28353 6131 28411 6137
rect 30650 6128 30656 6140
rect 30708 6128 30714 6180
rect 28902 6100 28908 6112
rect 27816 6072 28908 6100
rect 28902 6060 28908 6072
rect 28960 6060 28966 6112
rect 30668 6100 30696 6128
rect 33796 6112 33824 6199
rect 31205 6103 31263 6109
rect 31205 6100 31217 6103
rect 30668 6072 31217 6100
rect 31205 6069 31217 6072
rect 31251 6069 31263 6103
rect 31205 6063 31263 6069
rect 32306 6060 32312 6112
rect 32364 6060 32370 6112
rect 32858 6060 32864 6112
rect 32916 6060 32922 6112
rect 33778 6060 33784 6112
rect 33836 6060 33842 6112
rect 2760 6010 34316 6032
rect 2760 5958 7210 6010
rect 7262 5958 7274 6010
rect 7326 5958 7338 6010
rect 7390 5958 7402 6010
rect 7454 5958 7466 6010
rect 7518 5958 15099 6010
rect 15151 5958 15163 6010
rect 15215 5958 15227 6010
rect 15279 5958 15291 6010
rect 15343 5958 15355 6010
rect 15407 5958 22988 6010
rect 23040 5958 23052 6010
rect 23104 5958 23116 6010
rect 23168 5958 23180 6010
rect 23232 5958 23244 6010
rect 23296 5958 30877 6010
rect 30929 5958 30941 6010
rect 30993 5958 31005 6010
rect 31057 5958 31069 6010
rect 31121 5958 31133 6010
rect 31185 5958 34316 6010
rect 2760 5936 34316 5958
rect 3053 5899 3111 5905
rect 3053 5865 3065 5899
rect 3099 5896 3111 5899
rect 3142 5896 3148 5908
rect 3099 5868 3148 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 4246 5856 4252 5908
rect 4304 5856 4310 5908
rect 5258 5856 5264 5908
rect 5316 5856 5322 5908
rect 7098 5856 7104 5908
rect 7156 5896 7162 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 7156 5868 7481 5896
rect 7156 5856 7162 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 7469 5859 7527 5865
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 8021 5899 8079 5905
rect 8021 5896 8033 5899
rect 7984 5868 8033 5896
rect 7984 5856 7990 5868
rect 8021 5865 8033 5868
rect 8067 5865 8079 5899
rect 8021 5859 8079 5865
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8444 5868 9045 5896
rect 8444 5856 8450 5868
rect 9033 5865 9045 5868
rect 9079 5896 9091 5899
rect 9306 5896 9312 5908
rect 9079 5868 9312 5896
rect 9079 5865 9091 5868
rect 9033 5859 9091 5865
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 10229 5899 10287 5905
rect 10229 5896 10241 5899
rect 10100 5868 10241 5896
rect 10100 5856 10106 5868
rect 10229 5865 10241 5868
rect 10275 5896 10287 5899
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10275 5868 10701 5896
rect 10275 5865 10287 5868
rect 10229 5859 10287 5865
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 10689 5859 10747 5865
rect 10870 5856 10876 5908
rect 10928 5896 10934 5908
rect 11425 5899 11483 5905
rect 11425 5896 11437 5899
rect 10928 5868 11437 5896
rect 10928 5856 10934 5868
rect 11425 5865 11437 5868
rect 11471 5865 11483 5899
rect 11425 5859 11483 5865
rect 11698 5856 11704 5908
rect 11756 5856 11762 5908
rect 12158 5856 12164 5908
rect 12216 5856 12222 5908
rect 12802 5856 12808 5908
rect 12860 5896 12866 5908
rect 13541 5899 13599 5905
rect 13541 5896 13553 5899
rect 12860 5868 13553 5896
rect 12860 5856 12866 5868
rect 13541 5865 13553 5868
rect 13587 5896 13599 5899
rect 14001 5899 14059 5905
rect 14001 5896 14013 5899
rect 13587 5868 14013 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 14001 5865 14013 5868
rect 14047 5865 14059 5899
rect 16942 5896 16948 5908
rect 14001 5859 14059 5865
rect 14752 5868 16948 5896
rect 3234 5788 3240 5840
rect 3292 5828 3298 5840
rect 4264 5828 4292 5856
rect 3292 5800 3358 5828
rect 4264 5800 4844 5828
rect 3292 5788 3298 5800
rect 4816 5769 4844 5800
rect 4801 5763 4859 5769
rect 4801 5729 4813 5763
rect 4847 5760 4859 5763
rect 5074 5760 5080 5772
rect 4847 5732 5080 5760
rect 4847 5729 4859 5732
rect 4801 5723 4859 5729
rect 5074 5720 5080 5732
rect 5132 5720 5138 5772
rect 5276 5760 5304 5856
rect 6454 5788 6460 5840
rect 6512 5828 6518 5840
rect 7745 5831 7803 5837
rect 7745 5828 7757 5831
rect 6512 5800 7757 5828
rect 6512 5788 6518 5800
rect 7745 5797 7757 5800
rect 7791 5797 7803 5831
rect 8202 5828 8208 5840
rect 7745 5791 7803 5797
rect 7852 5800 8208 5828
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 5276 5732 6377 5760
rect 6365 5729 6377 5732
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 7561 5763 7619 5769
rect 7561 5729 7573 5763
rect 7607 5760 7619 5763
rect 7650 5760 7656 5772
rect 7607 5732 7656 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 7650 5720 7656 5732
rect 7708 5760 7714 5772
rect 7852 5769 7880 5800
rect 8202 5788 8208 5800
rect 8260 5828 8266 5840
rect 11716 5828 11744 5856
rect 8260 5800 10824 5828
rect 8260 5788 8266 5800
rect 10796 5772 10824 5800
rect 11348 5800 11744 5828
rect 7837 5763 7895 5769
rect 7837 5760 7849 5763
rect 7708 5732 7849 5760
rect 7708 5720 7714 5732
rect 7837 5729 7849 5732
rect 7883 5729 7895 5763
rect 10321 5763 10379 5769
rect 10321 5760 10333 5763
rect 7837 5723 7895 5729
rect 8680 5732 10333 5760
rect 8680 5704 8708 5732
rect 10321 5729 10333 5732
rect 10367 5729 10379 5763
rect 10321 5723 10379 5729
rect 10778 5720 10784 5772
rect 10836 5720 10842 5772
rect 11348 5769 11376 5800
rect 11790 5788 11796 5840
rect 11848 5788 11854 5840
rect 13354 5788 13360 5840
rect 13412 5828 13418 5840
rect 14752 5828 14780 5868
rect 16942 5856 16948 5868
rect 17000 5856 17006 5908
rect 17954 5856 17960 5908
rect 18012 5856 18018 5908
rect 20254 5856 20260 5908
rect 20312 5896 20318 5908
rect 21729 5899 21787 5905
rect 20312 5868 21680 5896
rect 20312 5856 20318 5868
rect 17405 5831 17463 5837
rect 17405 5828 17417 5831
rect 13412 5800 14780 5828
rect 16238 5800 17417 5828
rect 13412 5788 13418 5800
rect 11333 5763 11391 5769
rect 11333 5729 11345 5763
rect 11379 5729 11391 5763
rect 11333 5723 11391 5729
rect 11606 5720 11612 5772
rect 11664 5720 11670 5772
rect 11701 5763 11759 5769
rect 11701 5729 11713 5763
rect 11747 5729 11759 5763
rect 11701 5723 11759 5729
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4571 5664 4752 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4724 5624 4752 5664
rect 4890 5652 4896 5704
rect 4948 5692 4954 5704
rect 5629 5695 5687 5701
rect 5629 5692 5641 5695
rect 4948 5664 5641 5692
rect 4948 5652 4954 5664
rect 5629 5661 5641 5664
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 6733 5695 6791 5701
rect 6733 5661 6745 5695
rect 6779 5692 6791 5695
rect 6914 5692 6920 5704
rect 6779 5664 6920 5692
rect 6779 5661 6791 5664
rect 6733 5655 6791 5661
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 8570 5652 8576 5704
rect 8628 5652 8634 5704
rect 8662 5652 8668 5704
rect 8720 5652 8726 5704
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5692 9275 5695
rect 9263 5664 9904 5692
rect 9263 5661 9275 5664
rect 9217 5655 9275 5661
rect 9876 5633 9904 5664
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 5813 5627 5871 5633
rect 5813 5624 5825 5627
rect 4724 5596 5825 5624
rect 5813 5593 5825 5596
rect 5859 5593 5871 5627
rect 5813 5587 5871 5593
rect 9861 5627 9919 5633
rect 9861 5593 9873 5627
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 4982 5516 4988 5568
rect 5040 5556 5046 5568
rect 5077 5559 5135 5565
rect 5077 5556 5089 5559
rect 5040 5528 5089 5556
rect 5040 5516 5046 5528
rect 5077 5525 5089 5528
rect 5123 5525 5135 5559
rect 5077 5519 5135 5525
rect 7282 5516 7288 5568
rect 7340 5516 7346 5568
rect 9769 5559 9827 5565
rect 9769 5525 9781 5559
rect 9815 5556 9827 5559
rect 10042 5556 10048 5568
rect 9815 5528 10048 5556
rect 9815 5525 9827 5528
rect 9769 5519 9827 5525
rect 10042 5516 10048 5528
rect 10100 5516 10106 5568
rect 10428 5556 10456 5652
rect 11624 5624 11652 5720
rect 11716 5692 11744 5723
rect 11974 5720 11980 5772
rect 12032 5720 12038 5772
rect 12066 5720 12072 5772
rect 12124 5760 12130 5772
rect 12253 5763 12311 5769
rect 12253 5760 12265 5763
rect 12124 5732 12265 5760
rect 12124 5720 12130 5732
rect 12253 5729 12265 5732
rect 12299 5729 12311 5763
rect 12253 5723 12311 5729
rect 13633 5763 13691 5769
rect 13633 5729 13645 5763
rect 13679 5760 13691 5763
rect 14090 5760 14096 5772
rect 13679 5732 14096 5760
rect 13679 5729 13691 5732
rect 13633 5723 13691 5729
rect 14090 5720 14096 5732
rect 14148 5720 14154 5772
rect 14458 5720 14464 5772
rect 14516 5760 14522 5772
rect 14752 5769 14780 5800
rect 17405 5797 17417 5800
rect 17451 5797 17463 5831
rect 20993 5831 21051 5837
rect 20993 5828 21005 5831
rect 20562 5800 21005 5828
rect 17405 5791 17463 5797
rect 20993 5797 21005 5800
rect 21039 5797 21051 5831
rect 21652 5828 21680 5868
rect 21729 5865 21741 5899
rect 21775 5896 21787 5899
rect 21910 5896 21916 5908
rect 21775 5868 21916 5896
rect 21775 5865 21787 5868
rect 21729 5859 21787 5865
rect 21910 5856 21916 5868
rect 21968 5856 21974 5908
rect 23569 5899 23627 5905
rect 23569 5865 23581 5899
rect 23615 5896 23627 5899
rect 25498 5896 25504 5908
rect 23615 5868 25504 5896
rect 23615 5865 23627 5868
rect 23569 5859 23627 5865
rect 25498 5856 25504 5868
rect 25556 5856 25562 5908
rect 27246 5856 27252 5908
rect 27304 5856 27310 5908
rect 27341 5899 27399 5905
rect 27341 5865 27353 5899
rect 27387 5896 27399 5899
rect 27982 5896 27988 5908
rect 27387 5868 27988 5896
rect 27387 5865 27399 5868
rect 27341 5859 27399 5865
rect 27982 5856 27988 5868
rect 28040 5856 28046 5908
rect 29270 5896 29276 5908
rect 28368 5868 29276 5896
rect 23109 5831 23167 5837
rect 23109 5828 23121 5831
rect 21652 5800 23121 5828
rect 20993 5791 21051 5797
rect 23109 5797 23121 5800
rect 23155 5828 23167 5831
rect 23658 5828 23664 5840
rect 23155 5800 23664 5828
rect 23155 5797 23167 5800
rect 23109 5791 23167 5797
rect 23658 5788 23664 5800
rect 23716 5788 23722 5840
rect 25314 5788 25320 5840
rect 25372 5828 25378 5840
rect 27264 5828 27292 5856
rect 28368 5837 28396 5868
rect 29270 5856 29276 5868
rect 29328 5856 29334 5908
rect 30377 5899 30435 5905
rect 30377 5865 30389 5899
rect 30423 5896 30435 5899
rect 30558 5896 30564 5908
rect 30423 5868 30564 5896
rect 30423 5865 30435 5868
rect 30377 5859 30435 5865
rect 30558 5856 30564 5868
rect 30616 5856 30622 5908
rect 30650 5856 30656 5908
rect 30708 5896 30714 5908
rect 30837 5899 30895 5905
rect 30837 5896 30849 5899
rect 30708 5868 30849 5896
rect 30708 5856 30714 5868
rect 30837 5865 30849 5868
rect 30883 5865 30895 5899
rect 30837 5859 30895 5865
rect 31205 5899 31263 5905
rect 31205 5865 31217 5899
rect 31251 5896 31263 5899
rect 31754 5896 31760 5908
rect 31251 5868 31760 5896
rect 31251 5865 31263 5868
rect 31205 5859 31263 5865
rect 31754 5856 31760 5868
rect 31812 5856 31818 5908
rect 32858 5896 32864 5908
rect 32048 5868 32864 5896
rect 28353 5831 28411 5837
rect 28353 5828 28365 5831
rect 25372 5800 25728 5828
rect 27264 5800 28365 5828
rect 25372 5788 25378 5800
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 14516 5732 14565 5760
rect 14516 5720 14522 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 16758 5720 16764 5772
rect 16816 5760 16822 5772
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 16816 5732 17509 5760
rect 16816 5720 16822 5732
rect 17497 5729 17509 5732
rect 17543 5760 17555 5763
rect 17862 5760 17868 5772
rect 17543 5732 17868 5760
rect 17543 5729 17555 5732
rect 17497 5723 17555 5729
rect 17862 5720 17868 5732
rect 17920 5720 17926 5772
rect 21085 5763 21143 5769
rect 21085 5729 21097 5763
rect 21131 5760 21143 5763
rect 22186 5760 22192 5772
rect 21131 5732 22192 5760
rect 21131 5729 21143 5732
rect 21085 5723 21143 5729
rect 22186 5720 22192 5732
rect 22244 5720 22250 5772
rect 24210 5720 24216 5772
rect 24268 5720 24274 5772
rect 25501 5763 25559 5769
rect 25501 5760 25513 5763
rect 25056 5732 25513 5760
rect 11882 5692 11888 5704
rect 11716 5664 11888 5692
rect 11882 5652 11888 5664
rect 11940 5692 11946 5704
rect 12158 5692 12164 5704
rect 11940 5664 12164 5692
rect 11940 5652 11946 5664
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12342 5652 12348 5704
rect 12400 5652 12406 5704
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5661 13047 5695
rect 12989 5655 13047 5661
rect 12250 5624 12256 5636
rect 11624 5596 12256 5624
rect 12250 5584 12256 5596
rect 12308 5584 12314 5636
rect 13004 5624 13032 5655
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 15010 5652 15016 5704
rect 15068 5652 15074 5704
rect 17129 5695 17187 5701
rect 17129 5692 17141 5695
rect 16500 5664 17141 5692
rect 13173 5627 13231 5633
rect 13173 5624 13185 5627
rect 13004 5596 13185 5624
rect 13173 5593 13185 5596
rect 13219 5593 13231 5627
rect 13173 5587 13231 5593
rect 13722 5556 13728 5568
rect 10428 5528 13728 5556
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 16390 5516 16396 5568
rect 16448 5556 16454 5568
rect 16500 5565 16528 5664
rect 17129 5661 17141 5664
rect 17175 5661 17187 5695
rect 17129 5655 17187 5661
rect 18322 5652 18328 5704
rect 18380 5692 18386 5704
rect 19058 5692 19064 5704
rect 18380 5664 19064 5692
rect 18380 5652 18386 5664
rect 19058 5652 19064 5664
rect 19116 5652 19122 5704
rect 19334 5652 19340 5704
rect 19392 5652 19398 5704
rect 24302 5652 24308 5704
rect 24360 5701 24366 5704
rect 24360 5695 24409 5701
rect 24360 5661 24363 5695
rect 24397 5661 24409 5695
rect 24360 5655 24409 5661
rect 24360 5652 24366 5655
rect 24486 5652 24492 5704
rect 24544 5652 24550 5704
rect 24854 5652 24860 5704
rect 24912 5692 24918 5704
rect 25056 5692 25084 5732
rect 25501 5729 25513 5732
rect 25547 5729 25559 5763
rect 25700 5760 25728 5800
rect 28353 5797 28365 5800
rect 28399 5797 28411 5831
rect 29178 5828 29184 5840
rect 28353 5791 28411 5797
rect 28644 5800 29184 5828
rect 25700 5732 25820 5760
rect 25501 5723 25559 5729
rect 24912 5664 25084 5692
rect 24912 5652 24918 5664
rect 25222 5652 25228 5704
rect 25280 5652 25286 5704
rect 25406 5652 25412 5704
rect 25464 5652 25470 5704
rect 25682 5652 25688 5704
rect 25740 5652 25746 5704
rect 25792 5692 25820 5732
rect 26694 5720 26700 5772
rect 26752 5720 26758 5772
rect 27430 5720 27436 5772
rect 27488 5760 27494 5772
rect 28644 5769 28672 5800
rect 29178 5788 29184 5800
rect 29236 5788 29242 5840
rect 30745 5831 30803 5837
rect 30745 5797 30757 5831
rect 30791 5828 30803 5831
rect 31938 5828 31944 5840
rect 30791 5800 31944 5828
rect 30791 5797 30803 5800
rect 30745 5791 30803 5797
rect 31938 5788 31944 5800
rect 31996 5788 32002 5840
rect 32048 5837 32076 5868
rect 32858 5856 32864 5868
rect 32916 5856 32922 5908
rect 32033 5831 32091 5837
rect 32033 5797 32045 5831
rect 32079 5797 32091 5831
rect 33873 5831 33931 5837
rect 33873 5828 33885 5831
rect 33258 5800 33885 5828
rect 32033 5791 32091 5797
rect 33873 5797 33885 5800
rect 33919 5797 33931 5831
rect 33873 5791 33931 5797
rect 27617 5763 27675 5769
rect 27617 5760 27629 5763
rect 27488 5732 27629 5760
rect 27488 5720 27494 5732
rect 27617 5729 27629 5732
rect 27663 5729 27675 5763
rect 27617 5723 27675 5729
rect 28629 5763 28687 5769
rect 28629 5729 28641 5763
rect 28675 5729 28687 5763
rect 28629 5723 28687 5729
rect 30006 5720 30012 5772
rect 30064 5720 30070 5772
rect 30834 5720 30840 5772
rect 30892 5760 30898 5772
rect 31757 5763 31815 5769
rect 31757 5760 31769 5763
rect 30892 5732 31769 5760
rect 30892 5720 30898 5732
rect 31757 5729 31769 5732
rect 31803 5729 31815 5763
rect 31757 5723 31815 5729
rect 33778 5720 33784 5772
rect 33836 5720 33842 5772
rect 26145 5695 26203 5701
rect 26145 5692 26157 5695
rect 25792 5664 26157 5692
rect 22646 5584 22652 5636
rect 22704 5624 22710 5636
rect 22833 5627 22891 5633
rect 22833 5624 22845 5627
rect 22704 5596 22845 5624
rect 22704 5584 22710 5596
rect 22833 5593 22845 5596
rect 22879 5624 22891 5627
rect 24765 5627 24823 5633
rect 22879 5596 23888 5624
rect 22879 5593 22891 5596
rect 22833 5587 22891 5593
rect 16485 5559 16543 5565
rect 16485 5556 16497 5559
rect 16448 5528 16497 5556
rect 16448 5516 16454 5528
rect 16485 5525 16497 5528
rect 16531 5525 16543 5559
rect 16485 5519 16543 5525
rect 16574 5516 16580 5568
rect 16632 5516 16638 5568
rect 18690 5516 18696 5568
rect 18748 5516 18754 5568
rect 20806 5516 20812 5568
rect 20864 5516 20870 5568
rect 23860 5556 23888 5596
rect 24765 5593 24777 5627
rect 24811 5624 24823 5627
rect 25792 5624 25820 5664
rect 26145 5661 26157 5664
rect 26191 5661 26203 5695
rect 26421 5695 26479 5701
rect 26421 5692 26433 5695
rect 26145 5655 26203 5661
rect 26252 5664 26433 5692
rect 24811 5596 25820 5624
rect 24811 5593 24823 5596
rect 24765 5587 24823 5593
rect 24780 5556 24808 5587
rect 23860 5528 24808 5556
rect 26252 5556 26280 5664
rect 26421 5661 26433 5664
rect 26467 5661 26479 5695
rect 26421 5655 26479 5661
rect 26559 5695 26617 5701
rect 26559 5661 26571 5695
rect 26605 5692 26617 5695
rect 26605 5664 27752 5692
rect 26605 5661 26617 5664
rect 26559 5655 26617 5661
rect 27614 5624 27620 5636
rect 27448 5596 27620 5624
rect 27448 5556 27476 5596
rect 27614 5584 27620 5596
rect 27672 5584 27678 5636
rect 27724 5624 27752 5664
rect 27798 5652 27804 5704
rect 27856 5652 27862 5704
rect 28166 5652 28172 5704
rect 28224 5652 28230 5704
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5692 28963 5695
rect 29362 5692 29368 5704
rect 28951 5664 29368 5692
rect 28951 5661 28963 5664
rect 28905 5655 28963 5661
rect 29362 5652 29368 5664
rect 29420 5652 29426 5704
rect 29546 5652 29552 5704
rect 29604 5692 29610 5704
rect 30561 5695 30619 5701
rect 30561 5692 30573 5695
rect 29604 5664 30573 5692
rect 29604 5652 29610 5664
rect 30561 5661 30573 5664
rect 30607 5692 30619 5695
rect 31478 5692 31484 5704
rect 30607 5664 31484 5692
rect 30607 5661 30619 5664
rect 30561 5655 30619 5661
rect 31478 5652 31484 5664
rect 31536 5652 31542 5704
rect 33796 5692 33824 5720
rect 33152 5664 33824 5692
rect 28184 5624 28212 5652
rect 33152 5636 33180 5664
rect 27724 5596 28212 5624
rect 33134 5584 33140 5636
rect 33192 5584 33198 5636
rect 26252 5528 27476 5556
rect 27522 5516 27528 5568
rect 27580 5516 27586 5568
rect 32398 5516 32404 5568
rect 32456 5556 32462 5568
rect 33505 5559 33563 5565
rect 33505 5556 33517 5559
rect 32456 5528 33517 5556
rect 32456 5516 32462 5528
rect 33505 5525 33517 5528
rect 33551 5525 33563 5559
rect 33505 5519 33563 5525
rect 2760 5466 34316 5488
rect 2760 5414 6550 5466
rect 6602 5414 6614 5466
rect 6666 5414 6678 5466
rect 6730 5414 6742 5466
rect 6794 5414 6806 5466
rect 6858 5414 14439 5466
rect 14491 5414 14503 5466
rect 14555 5414 14567 5466
rect 14619 5414 14631 5466
rect 14683 5414 14695 5466
rect 14747 5414 22328 5466
rect 22380 5414 22392 5466
rect 22444 5414 22456 5466
rect 22508 5414 22520 5466
rect 22572 5414 22584 5466
rect 22636 5414 30217 5466
rect 30269 5414 30281 5466
rect 30333 5414 30345 5466
rect 30397 5414 30409 5466
rect 30461 5414 30473 5466
rect 30525 5414 34316 5466
rect 2760 5392 34316 5414
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8570 5352 8576 5364
rect 7975 5324 8576 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 9824 5324 10548 5352
rect 9824 5312 9830 5324
rect 4172 5256 5120 5284
rect 4172 5228 4200 5256
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4982 5176 4988 5228
rect 5040 5176 5046 5228
rect 5092 5225 5120 5256
rect 7116 5256 7972 5284
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5534 5216 5540 5228
rect 5123 5188 5540 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 7116 5216 7144 5256
rect 7944 5228 7972 5256
rect 5736 5188 7144 5216
rect 7193 5219 7251 5225
rect 4433 5151 4491 5157
rect 4433 5117 4445 5151
rect 4479 5148 4491 5151
rect 5736 5148 5764 5188
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7834 5216 7840 5228
rect 7239 5188 7840 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7834 5176 7840 5188
rect 7892 5176 7898 5228
rect 7926 5176 7932 5228
rect 7984 5176 7990 5228
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5216 8171 5219
rect 8294 5216 8300 5228
rect 8159 5188 8300 5216
rect 8159 5185 8171 5188
rect 8113 5179 8171 5185
rect 8294 5176 8300 5188
rect 8352 5216 8358 5228
rect 8478 5216 8484 5228
rect 8352 5188 8484 5216
rect 8352 5176 8358 5188
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 10134 5176 10140 5228
rect 10192 5216 10198 5228
rect 10413 5219 10471 5225
rect 10413 5216 10425 5219
rect 10192 5188 10425 5216
rect 10192 5176 10198 5188
rect 10413 5185 10425 5188
rect 10459 5185 10471 5219
rect 10520 5216 10548 5324
rect 11514 5312 11520 5364
rect 11572 5312 11578 5364
rect 11882 5312 11888 5364
rect 11940 5352 11946 5364
rect 11940 5324 14044 5352
rect 11940 5312 11946 5324
rect 11532 5225 11560 5312
rect 14016 5284 14044 5324
rect 14090 5312 14096 5364
rect 14148 5312 14154 5364
rect 14182 5312 14188 5364
rect 14240 5352 14246 5364
rect 14277 5355 14335 5361
rect 14277 5352 14289 5355
rect 14240 5324 14289 5352
rect 14240 5312 14246 5324
rect 14277 5321 14289 5324
rect 14323 5321 14335 5355
rect 14277 5315 14335 5321
rect 14829 5355 14887 5361
rect 14829 5321 14841 5355
rect 14875 5352 14887 5355
rect 15010 5352 15016 5364
rect 14875 5324 15016 5352
rect 14875 5321 14887 5324
rect 14829 5315 14887 5321
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 15654 5312 15660 5364
rect 15712 5352 15718 5364
rect 15933 5355 15991 5361
rect 15933 5352 15945 5355
rect 15712 5324 15945 5352
rect 15712 5312 15718 5324
rect 15933 5321 15945 5324
rect 15979 5321 15991 5355
rect 15933 5315 15991 5321
rect 16022 5312 16028 5364
rect 16080 5352 16086 5364
rect 18598 5352 18604 5364
rect 16080 5324 18604 5352
rect 16080 5312 16086 5324
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 19334 5312 19340 5364
rect 19392 5352 19398 5364
rect 19521 5355 19579 5361
rect 19521 5352 19533 5355
rect 19392 5324 19533 5352
rect 19392 5312 19398 5324
rect 19521 5321 19533 5324
rect 19567 5321 19579 5355
rect 19521 5315 19579 5321
rect 19794 5312 19800 5364
rect 19852 5352 19858 5364
rect 20441 5355 20499 5361
rect 20441 5352 20453 5355
rect 19852 5324 20453 5352
rect 19852 5312 19858 5324
rect 20441 5321 20453 5324
rect 20487 5321 20499 5355
rect 20441 5315 20499 5321
rect 21726 5312 21732 5364
rect 21784 5312 21790 5364
rect 23293 5355 23351 5361
rect 23293 5321 23305 5355
rect 23339 5352 23351 5355
rect 23566 5352 23572 5364
rect 23339 5324 23572 5352
rect 23339 5321 23351 5324
rect 23293 5315 23351 5321
rect 23566 5312 23572 5324
rect 23624 5312 23630 5364
rect 23750 5312 23756 5364
rect 23808 5352 23814 5364
rect 24121 5355 24179 5361
rect 24121 5352 24133 5355
rect 23808 5324 24133 5352
rect 23808 5312 23814 5324
rect 24121 5321 24133 5324
rect 24167 5321 24179 5355
rect 24121 5315 24179 5321
rect 24210 5312 24216 5364
rect 24268 5312 24274 5364
rect 26697 5355 26755 5361
rect 26697 5321 26709 5355
rect 26743 5352 26755 5355
rect 27798 5352 27804 5364
rect 26743 5324 27804 5352
rect 26743 5321 26755 5324
rect 26697 5315 26755 5321
rect 27798 5312 27804 5324
rect 27856 5312 27862 5364
rect 30006 5312 30012 5364
rect 30064 5352 30070 5364
rect 30101 5355 30159 5361
rect 30101 5352 30113 5355
rect 30064 5324 30113 5352
rect 30064 5312 30070 5324
rect 30101 5321 30113 5324
rect 30147 5321 30159 5355
rect 30101 5315 30159 5321
rect 23017 5287 23075 5293
rect 14016 5256 19564 5284
rect 19536 5228 19564 5256
rect 23017 5253 23029 5287
rect 23063 5284 23075 5287
rect 24228 5284 24256 5312
rect 23063 5256 24256 5284
rect 25869 5287 25927 5293
rect 23063 5253 23075 5256
rect 23017 5247 23075 5253
rect 25869 5253 25881 5287
rect 25915 5284 25927 5287
rect 26602 5284 26608 5296
rect 25915 5256 26608 5284
rect 25915 5253 25927 5256
rect 25869 5247 25927 5253
rect 26602 5244 26608 5256
rect 26660 5244 26666 5296
rect 28902 5244 28908 5296
rect 28960 5284 28966 5296
rect 30469 5287 30527 5293
rect 30469 5284 30481 5287
rect 28960 5256 30481 5284
rect 28960 5244 28966 5256
rect 30469 5253 30481 5256
rect 30515 5253 30527 5287
rect 30469 5247 30527 5253
rect 31202 5244 31208 5296
rect 31260 5284 31266 5296
rect 31260 5256 32628 5284
rect 31260 5244 31266 5256
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 10520 5188 11161 5216
rect 10413 5179 10471 5185
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 12342 5216 12348 5228
rect 11839 5188 12348 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 13780 5188 15393 5216
rect 13780 5176 13786 5188
rect 15381 5185 15393 5188
rect 15427 5216 15439 5219
rect 16298 5216 16304 5228
rect 15427 5188 16304 5216
rect 15427 5185 15439 5188
rect 15381 5179 15439 5185
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 16574 5176 16580 5228
rect 16632 5176 16638 5228
rect 16850 5176 16856 5228
rect 16908 5176 16914 5228
rect 19150 5216 19156 5228
rect 17880 5188 19156 5216
rect 4479 5120 5764 5148
rect 4479 5117 4491 5120
rect 4433 5111 4491 5117
rect 7282 5108 7288 5160
rect 7340 5108 7346 5160
rect 7650 5108 7656 5160
rect 7708 5108 7714 5160
rect 8205 5151 8263 5157
rect 8205 5117 8217 5151
rect 8251 5148 8263 5151
rect 8846 5148 8852 5160
rect 8251 5120 8852 5148
rect 8251 5117 8263 5120
rect 8205 5111 8263 5117
rect 3234 5040 3240 5092
rect 3292 5040 3298 5092
rect 4893 5083 4951 5089
rect 4893 5049 4905 5083
rect 4939 5080 4951 5083
rect 4939 5052 5580 5080
rect 4939 5049 4951 5052
rect 4893 5043 4951 5049
rect 4522 4972 4528 5024
rect 4580 4972 4586 5024
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 5445 5015 5503 5021
rect 5445 5012 5457 5015
rect 5316 4984 5457 5012
rect 5316 4972 5322 4984
rect 5445 4981 5457 4984
rect 5491 4981 5503 5015
rect 5552 5012 5580 5052
rect 6454 5040 6460 5092
rect 6512 5040 6518 5092
rect 6917 5083 6975 5089
rect 6917 5049 6929 5083
rect 6963 5080 6975 5083
rect 7300 5080 7328 5108
rect 6963 5052 7328 5080
rect 7561 5083 7619 5089
rect 6963 5049 6975 5052
rect 6917 5043 6975 5049
rect 7561 5049 7573 5083
rect 7607 5080 7619 5083
rect 8220 5080 8248 5111
rect 8846 5108 8852 5120
rect 8904 5108 8910 5160
rect 13262 5108 13268 5160
rect 13320 5148 13326 5160
rect 13449 5151 13507 5157
rect 13449 5148 13461 5151
rect 13320 5120 13461 5148
rect 13320 5108 13326 5120
rect 13449 5117 13461 5120
rect 13495 5117 13507 5151
rect 13449 5111 13507 5117
rect 14185 5151 14243 5157
rect 14185 5117 14197 5151
rect 14231 5148 14243 5151
rect 14645 5151 14703 5157
rect 14645 5148 14657 5151
rect 14231 5120 14657 5148
rect 14231 5117 14243 5120
rect 14185 5111 14243 5117
rect 14645 5117 14657 5120
rect 14691 5148 14703 5151
rect 14826 5148 14832 5160
rect 14691 5120 14832 5148
rect 14691 5117 14703 5120
rect 14645 5111 14703 5117
rect 14826 5108 14832 5120
rect 14884 5108 14890 5160
rect 15289 5151 15347 5157
rect 15289 5117 15301 5151
rect 15335 5148 15347 5151
rect 16592 5148 16620 5176
rect 15335 5120 16620 5148
rect 15335 5117 15347 5120
rect 15289 5111 15347 5117
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 7607 5052 8248 5080
rect 7607 5049 7619 5052
rect 7561 5043 7619 5049
rect 8386 5040 8392 5092
rect 8444 5080 8450 5092
rect 8481 5083 8539 5089
rect 8481 5080 8493 5083
rect 8444 5052 8493 5080
rect 8444 5040 8450 5052
rect 8481 5049 8493 5052
rect 8527 5049 8539 5083
rect 8481 5043 8539 5049
rect 8570 5040 8576 5092
rect 8628 5080 8634 5092
rect 8628 5052 8892 5080
rect 8628 5040 8634 5052
rect 5902 5012 5908 5024
rect 5552 4984 5908 5012
rect 5445 4975 5503 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 7742 4972 7748 5024
rect 7800 4972 7806 5024
rect 8662 4972 8668 5024
rect 8720 4972 8726 5024
rect 8864 5012 8892 5052
rect 9674 5040 9680 5092
rect 9732 5040 9738 5092
rect 10042 5040 10048 5092
rect 10100 5080 10106 5092
rect 10137 5083 10195 5089
rect 10137 5080 10149 5083
rect 10100 5052 10149 5080
rect 10100 5040 10106 5052
rect 10137 5049 10149 5052
rect 10183 5049 10195 5083
rect 14553 5083 14611 5089
rect 14553 5080 14565 5083
rect 13018 5052 14565 5080
rect 10137 5043 10195 5049
rect 14553 5049 14565 5052
rect 14599 5049 14611 5083
rect 14553 5043 14611 5049
rect 15197 5083 15255 5089
rect 15197 5049 15209 5083
rect 15243 5080 15255 5083
rect 17880 5080 17908 5188
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 19518 5176 19524 5228
rect 19576 5176 19582 5228
rect 19610 5176 19616 5228
rect 19668 5216 19674 5228
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 19668 5188 20085 5216
rect 19668 5176 19674 5188
rect 20073 5185 20085 5188
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 20806 5176 20812 5228
rect 20864 5216 20870 5228
rect 21085 5219 21143 5225
rect 21085 5216 21097 5219
rect 20864 5188 21097 5216
rect 20864 5176 20870 5188
rect 21085 5185 21097 5188
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 22830 5176 22836 5228
rect 22888 5216 22894 5228
rect 24765 5219 24823 5225
rect 22888 5188 23796 5216
rect 22888 5176 22894 5188
rect 17957 5151 18015 5157
rect 17957 5117 17969 5151
rect 18003 5117 18015 5151
rect 17957 5111 18015 5117
rect 18509 5151 18567 5157
rect 18509 5117 18521 5151
rect 18555 5148 18567 5151
rect 18966 5148 18972 5160
rect 18555 5120 18972 5148
rect 18555 5117 18567 5120
rect 18509 5111 18567 5117
rect 15243 5052 17908 5080
rect 15243 5049 15255 5052
rect 15197 5043 15255 5049
rect 17972 5024 18000 5111
rect 18966 5108 18972 5120
rect 19024 5108 19030 5160
rect 19061 5151 19119 5157
rect 19061 5117 19073 5151
rect 19107 5148 19119 5151
rect 20346 5148 20352 5160
rect 19107 5120 20352 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 20346 5108 20352 5120
rect 20404 5108 20410 5160
rect 23382 5108 23388 5160
rect 23440 5148 23446 5160
rect 23661 5151 23719 5157
rect 23661 5148 23673 5151
rect 23440 5120 23673 5148
rect 23440 5108 23446 5120
rect 23661 5117 23673 5120
rect 23707 5117 23719 5151
rect 23768 5148 23796 5188
rect 24765 5185 24777 5219
rect 24811 5216 24823 5219
rect 24946 5216 24952 5228
rect 24811 5188 24952 5216
rect 24811 5185 24823 5188
rect 24765 5179 24823 5185
rect 24946 5176 24952 5188
rect 25004 5176 25010 5228
rect 25317 5219 25375 5225
rect 25317 5185 25329 5219
rect 25363 5216 25375 5219
rect 25958 5216 25964 5228
rect 25363 5188 25964 5216
rect 25363 5185 25375 5188
rect 25317 5179 25375 5185
rect 25958 5176 25964 5188
rect 26016 5176 26022 5228
rect 26329 5219 26387 5225
rect 26329 5185 26341 5219
rect 26375 5216 26387 5219
rect 26694 5216 26700 5228
rect 26375 5188 26700 5216
rect 26375 5185 26387 5188
rect 26329 5179 26387 5185
rect 26694 5176 26700 5188
rect 26752 5176 26758 5228
rect 27706 5176 27712 5228
rect 27764 5216 27770 5228
rect 28169 5219 28227 5225
rect 28169 5216 28181 5219
rect 27764 5188 28181 5216
rect 27764 5176 27770 5188
rect 28169 5185 28181 5188
rect 28215 5185 28227 5219
rect 28169 5179 28227 5185
rect 28442 5176 28448 5228
rect 28500 5216 28506 5228
rect 29178 5216 29184 5228
rect 28500 5188 29184 5216
rect 28500 5176 28506 5188
rect 29178 5176 29184 5188
rect 29236 5216 29242 5228
rect 30742 5216 30748 5228
rect 29236 5188 30748 5216
rect 29236 5176 29242 5188
rect 30742 5176 30748 5188
rect 30800 5176 30806 5228
rect 31754 5176 31760 5228
rect 31812 5176 31818 5228
rect 25501 5151 25559 5157
rect 25501 5148 25513 5151
rect 23768 5120 25513 5148
rect 23661 5111 23719 5117
rect 25501 5117 25513 5120
rect 25547 5117 25559 5151
rect 25501 5111 25559 5117
rect 28626 5108 28632 5160
rect 28684 5148 28690 5160
rect 29089 5151 29147 5157
rect 29089 5148 29101 5151
rect 28684 5120 29101 5148
rect 28684 5108 28690 5120
rect 29089 5117 29101 5120
rect 29135 5117 29147 5151
rect 29089 5111 29147 5117
rect 29822 5108 29828 5160
rect 29880 5108 29886 5160
rect 30006 5108 30012 5160
rect 30064 5148 30070 5160
rect 32600 5157 32628 5256
rect 33781 5219 33839 5225
rect 33781 5185 33793 5219
rect 33827 5216 33839 5219
rect 34882 5216 34888 5228
rect 33827 5188 34888 5216
rect 33827 5185 33839 5188
rect 33781 5179 33839 5185
rect 34882 5176 34888 5188
rect 34940 5176 34946 5228
rect 30193 5151 30251 5157
rect 30193 5148 30205 5151
rect 30064 5120 30205 5148
rect 30064 5108 30070 5120
rect 30193 5117 30205 5120
rect 30239 5148 30251 5151
rect 32125 5151 32183 5157
rect 32125 5148 32137 5151
rect 30239 5120 32137 5148
rect 30239 5117 30251 5120
rect 30193 5111 30251 5117
rect 32125 5117 32137 5120
rect 32171 5148 32183 5151
rect 32585 5151 32643 5157
rect 32171 5120 32536 5148
rect 32171 5117 32183 5120
rect 32125 5111 32183 5117
rect 20070 5040 20076 5092
rect 20128 5080 20134 5092
rect 20128 5052 26924 5080
rect 20128 5040 20134 5052
rect 10597 5015 10655 5021
rect 10597 5012 10609 5015
rect 8864 4984 10609 5012
rect 10597 4981 10609 4984
rect 10643 4981 10655 5015
rect 10597 4975 10655 4981
rect 13262 4972 13268 5024
rect 13320 4972 13326 5024
rect 16298 4972 16304 5024
rect 16356 4972 16362 5024
rect 16761 5015 16819 5021
rect 16761 4981 16773 5015
rect 16807 5012 16819 5015
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 16807 4984 17325 5012
rect 16807 4981 16819 4984
rect 16761 4975 16819 4981
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 17313 4975 17371 4981
rect 17954 4972 17960 5024
rect 18012 4972 18018 5024
rect 19150 4972 19156 5024
rect 19208 4972 19214 5024
rect 23753 5015 23811 5021
rect 23753 4981 23765 5015
rect 23799 5012 23811 5015
rect 23842 5012 23848 5024
rect 23799 4984 23848 5012
rect 23799 4981 23811 4984
rect 23753 4975 23811 4981
rect 23842 4972 23848 4984
rect 23900 4972 23906 5024
rect 25406 4972 25412 5024
rect 25464 4972 25470 5024
rect 26896 5012 26924 5052
rect 27522 5040 27528 5092
rect 27580 5040 27586 5092
rect 32508 5080 32536 5120
rect 32585 5117 32597 5151
rect 32631 5117 32643 5151
rect 32585 5111 32643 5117
rect 33134 5080 33140 5092
rect 28276 5052 32260 5080
rect 32508 5052 33140 5080
rect 28276 5012 28304 5052
rect 32232 5024 32260 5052
rect 33134 5040 33140 5052
rect 33192 5040 33198 5092
rect 26896 4984 28304 5012
rect 28534 4972 28540 5024
rect 28592 4972 28598 5024
rect 29086 4972 29092 5024
rect 29144 5012 29150 5024
rect 29273 5015 29331 5021
rect 29273 5012 29285 5015
rect 29144 4984 29285 5012
rect 29144 4972 29150 4984
rect 29273 4981 29285 4984
rect 29319 4981 29331 5015
rect 29273 4975 29331 4981
rect 31202 4972 31208 5024
rect 31260 4972 31266 5024
rect 32030 4972 32036 5024
rect 32088 4972 32094 5024
rect 32214 4972 32220 5024
rect 32272 4972 32278 5024
rect 2760 4922 34316 4944
rect 2760 4870 7210 4922
rect 7262 4870 7274 4922
rect 7326 4870 7338 4922
rect 7390 4870 7402 4922
rect 7454 4870 7466 4922
rect 7518 4870 15099 4922
rect 15151 4870 15163 4922
rect 15215 4870 15227 4922
rect 15279 4870 15291 4922
rect 15343 4870 15355 4922
rect 15407 4870 22988 4922
rect 23040 4870 23052 4922
rect 23104 4870 23116 4922
rect 23168 4870 23180 4922
rect 23232 4870 23244 4922
rect 23296 4870 30877 4922
rect 30929 4870 30941 4922
rect 30993 4870 31005 4922
rect 31057 4870 31069 4922
rect 31121 4870 31133 4922
rect 31185 4870 34316 4922
rect 2760 4848 34316 4870
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 4890 4808 4896 4820
rect 3375 4780 4896 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 5350 4768 5356 4820
rect 5408 4768 5414 4820
rect 5442 4768 5448 4820
rect 5500 4768 5506 4820
rect 6270 4808 6276 4820
rect 6012 4780 6276 4808
rect 5261 4743 5319 4749
rect 5261 4740 5273 4743
rect 4370 4712 5273 4740
rect 5261 4709 5273 4712
rect 5307 4709 5319 4743
rect 5261 4703 5319 4709
rect 1302 4632 1308 4684
rect 1360 4672 1366 4684
rect 5368 4681 5396 4768
rect 5721 4743 5779 4749
rect 5721 4709 5733 4743
rect 5767 4740 5779 4743
rect 5902 4740 5908 4752
rect 5767 4712 5908 4740
rect 5767 4709 5779 4712
rect 5721 4703 5779 4709
rect 5902 4700 5908 4712
rect 5960 4700 5966 4752
rect 3053 4675 3111 4681
rect 3053 4672 3065 4675
rect 1360 4644 3065 4672
rect 1360 4632 1366 4644
rect 3053 4641 3065 4644
rect 3099 4641 3111 4675
rect 3053 4635 3111 4641
rect 5353 4675 5411 4681
rect 5353 4641 5365 4675
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 5626 4632 5632 4684
rect 5684 4632 5690 4684
rect 5810 4632 5816 4684
rect 5868 4632 5874 4684
rect 6012 4681 6040 4780
rect 6270 4768 6276 4780
rect 6328 4768 6334 4820
rect 6362 4768 6368 4820
rect 6420 4808 6426 4820
rect 6549 4811 6607 4817
rect 6549 4808 6561 4811
rect 6420 4780 6561 4808
rect 6420 4768 6426 4780
rect 6549 4777 6561 4780
rect 6595 4777 6607 4811
rect 6549 4771 6607 4777
rect 6914 4768 6920 4820
rect 6972 4768 6978 4820
rect 7668 4780 9168 4808
rect 6086 4700 6092 4752
rect 6144 4740 6150 4752
rect 7668 4740 7696 4780
rect 6144 4712 7696 4740
rect 6144 4700 6150 4712
rect 7742 4700 7748 4752
rect 7800 4740 7806 4752
rect 9140 4740 9168 4780
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 10689 4811 10747 4817
rect 10689 4808 10701 4811
rect 9732 4780 10701 4808
rect 9732 4768 9738 4780
rect 10689 4777 10701 4780
rect 10735 4777 10747 4811
rect 10689 4771 10747 4777
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 11885 4811 11943 4817
rect 11885 4808 11897 4811
rect 11848 4780 11897 4808
rect 11848 4768 11854 4780
rect 11885 4777 11897 4780
rect 11931 4777 11943 4811
rect 11885 4771 11943 4777
rect 12250 4768 12256 4820
rect 12308 4768 12314 4820
rect 15930 4808 15936 4820
rect 12406 4780 15936 4808
rect 12406 4740 12434 4780
rect 15930 4768 15936 4780
rect 15988 4768 15994 4820
rect 16942 4808 16948 4820
rect 16040 4780 16948 4808
rect 15286 4740 15292 4752
rect 7800 4712 8326 4740
rect 9140 4712 12434 4740
rect 14858 4712 15292 4740
rect 7800 4700 7806 4712
rect 15286 4700 15292 4712
rect 15344 4700 15350 4752
rect 5997 4675 6055 4681
rect 5997 4641 6009 4675
rect 6043 4641 6055 4675
rect 6457 4675 6515 4681
rect 6457 4672 6469 4675
rect 5997 4635 6055 4641
rect 6104 4644 6469 4672
rect 4798 4564 4804 4616
rect 4856 4564 4862 4616
rect 5074 4564 5080 4616
rect 5132 4564 5138 4616
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 6104 4604 6132 4644
rect 6457 4641 6469 4644
rect 6503 4641 6515 4675
rect 7193 4675 7251 4681
rect 7193 4672 7205 4675
rect 6457 4635 6515 4641
rect 6656 4644 7205 4672
rect 5316 4576 6132 4604
rect 5316 4564 5322 4576
rect 6362 4564 6368 4616
rect 6420 4604 6426 4616
rect 6656 4604 6684 4644
rect 7193 4641 7205 4644
rect 7239 4641 7251 4675
rect 7193 4635 7251 4641
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 10134 4672 10140 4684
rect 9815 4644 10140 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 10134 4632 10140 4644
rect 10192 4632 10198 4684
rect 10778 4632 10784 4684
rect 10836 4632 10842 4684
rect 11790 4632 11796 4684
rect 11848 4672 11854 4684
rect 16040 4681 16068 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 17862 4768 17868 4820
rect 17920 4808 17926 4820
rect 17920 4780 18092 4808
rect 17920 4768 17926 4780
rect 16298 4700 16304 4752
rect 16356 4700 16362 4752
rect 17957 4743 18015 4749
rect 17957 4740 17969 4743
rect 17526 4712 17969 4740
rect 17957 4709 17969 4712
rect 18003 4709 18015 4743
rect 17957 4703 18015 4709
rect 18064 4681 18092 4780
rect 20070 4768 20076 4820
rect 20128 4768 20134 4820
rect 23382 4768 23388 4820
rect 23440 4768 23446 4820
rect 24762 4808 24768 4820
rect 23676 4780 24768 4808
rect 19150 4700 19156 4752
rect 19208 4700 19214 4752
rect 23109 4743 23167 4749
rect 23109 4740 23121 4743
rect 21482 4712 23121 4740
rect 23109 4709 23121 4712
rect 23155 4709 23167 4743
rect 23109 4703 23167 4709
rect 12897 4675 12955 4681
rect 12897 4672 12909 4675
rect 11848 4644 12909 4672
rect 11848 4632 11854 4644
rect 12897 4641 12909 4644
rect 12943 4641 12955 4675
rect 12897 4635 12955 4641
rect 16025 4675 16083 4681
rect 16025 4641 16037 4675
rect 16071 4641 16083 4675
rect 16025 4635 16083 4641
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4641 18107 4675
rect 18049 4635 18107 4641
rect 18322 4632 18328 4684
rect 18380 4632 18386 4684
rect 22189 4675 22247 4681
rect 22189 4641 22201 4675
rect 22235 4672 22247 4675
rect 23201 4675 23259 4681
rect 22235 4644 23152 4672
rect 22235 4641 22247 4644
rect 22189 4635 22247 4641
rect 6420 4576 6684 4604
rect 7668 4576 8524 4604
rect 6420 4564 6426 4576
rect 3237 4471 3295 4477
rect 3237 4437 3249 4471
rect 3283 4468 3295 4471
rect 7668 4468 7696 4576
rect 7926 4496 7932 4548
rect 7984 4536 7990 4548
rect 8021 4539 8079 4545
rect 8021 4536 8033 4539
rect 7984 4508 8033 4536
rect 7984 4496 7990 4508
rect 8021 4505 8033 4508
rect 8067 4536 8079 4539
rect 8386 4536 8392 4548
rect 8067 4508 8392 4536
rect 8067 4505 8079 4508
rect 8021 4499 8079 4505
rect 8386 4496 8392 4508
rect 8444 4496 8450 4548
rect 3283 4440 7696 4468
rect 7837 4471 7895 4477
rect 3283 4437 3295 4440
rect 3237 4431 3295 4437
rect 7837 4437 7849 4471
rect 7883 4468 7895 4471
rect 8294 4468 8300 4480
rect 7883 4440 8300 4468
rect 7883 4437 7895 4440
rect 7837 4431 7895 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 8496 4468 8524 4576
rect 9490 4564 9496 4616
rect 9548 4564 9554 4616
rect 11882 4564 11888 4616
rect 11940 4564 11946 4616
rect 13354 4564 13360 4616
rect 13412 4564 13418 4616
rect 13630 4564 13636 4616
rect 13688 4564 13694 4616
rect 15105 4607 15163 4613
rect 15105 4573 15117 4607
rect 15151 4604 15163 4607
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15151 4576 15853 4604
rect 15151 4573 15163 4576
rect 15105 4567 15163 4573
rect 15841 4573 15853 4576
rect 15887 4604 15899 4607
rect 16758 4604 16764 4616
rect 15887 4576 16764 4604
rect 15887 4573 15899 4576
rect 15841 4567 15899 4573
rect 16758 4564 16764 4576
rect 16816 4564 16822 4616
rect 18598 4564 18604 4616
rect 18656 4564 18662 4616
rect 21913 4607 21971 4613
rect 21913 4573 21925 4607
rect 21959 4604 21971 4607
rect 22281 4607 22339 4613
rect 22281 4604 22293 4607
rect 21959 4576 22293 4604
rect 21959 4573 21971 4576
rect 21913 4567 21971 4573
rect 22281 4573 22293 4576
rect 22327 4573 22339 4607
rect 22281 4567 22339 4573
rect 22830 4564 22836 4616
rect 22888 4564 22894 4616
rect 23124 4604 23152 4644
rect 23201 4641 23213 4675
rect 23247 4672 23259 4675
rect 23400 4672 23428 4768
rect 23247 4644 23428 4672
rect 23247 4641 23259 4644
rect 23201 4635 23259 4641
rect 23676 4604 23704 4780
rect 24762 4768 24768 4780
rect 24820 4808 24826 4820
rect 24820 4780 25268 4808
rect 24820 4768 24826 4780
rect 23842 4632 23848 4684
rect 23900 4632 23906 4684
rect 25240 4681 25268 4780
rect 25406 4768 25412 4820
rect 25464 4808 25470 4820
rect 27157 4811 27215 4817
rect 27157 4808 27169 4811
rect 25464 4780 27169 4808
rect 25464 4768 25470 4780
rect 27157 4777 27169 4780
rect 27203 4777 27215 4811
rect 27157 4771 27215 4777
rect 28166 4768 28172 4820
rect 28224 4768 28230 4820
rect 28626 4768 28632 4820
rect 28684 4768 28690 4820
rect 28994 4768 29000 4820
rect 29052 4768 29058 4820
rect 29086 4768 29092 4820
rect 29144 4768 29150 4820
rect 31202 4808 31208 4820
rect 30392 4780 31208 4808
rect 26878 4740 26884 4752
rect 26818 4712 26884 4740
rect 26878 4700 26884 4712
rect 26936 4700 26942 4752
rect 29546 4740 29552 4752
rect 26988 4712 29552 4740
rect 25225 4675 25283 4681
rect 25225 4641 25237 4675
rect 25271 4672 25283 4675
rect 25317 4675 25375 4681
rect 25317 4672 25329 4675
rect 25271 4644 25329 4672
rect 25271 4641 25283 4644
rect 25225 4635 25283 4641
rect 25317 4641 25329 4644
rect 25363 4641 25375 4675
rect 25317 4635 25375 4641
rect 23124 4576 23704 4604
rect 24946 4564 24952 4616
rect 25004 4564 25010 4616
rect 25590 4564 25596 4616
rect 25648 4564 25654 4616
rect 25958 4564 25964 4616
rect 26016 4604 26022 4616
rect 26988 4604 27016 4712
rect 29546 4700 29552 4712
rect 29604 4700 29610 4752
rect 30392 4749 30420 4780
rect 31202 4768 31208 4780
rect 31260 4768 31266 4820
rect 31849 4811 31907 4817
rect 31849 4777 31861 4811
rect 31895 4808 31907 4811
rect 31938 4808 31944 4820
rect 31895 4780 31944 4808
rect 31895 4777 31907 4780
rect 31849 4771 31907 4777
rect 31938 4768 31944 4780
rect 31996 4768 32002 4820
rect 30377 4743 30435 4749
rect 30377 4709 30389 4743
rect 30423 4709 30435 4743
rect 32030 4740 32036 4752
rect 31602 4712 32036 4740
rect 30377 4703 30435 4709
rect 32030 4700 32036 4712
rect 32088 4700 32094 4752
rect 27430 4632 27436 4684
rect 27488 4672 27494 4684
rect 29641 4675 29699 4681
rect 29641 4672 29653 4675
rect 27488 4644 29653 4672
rect 27488 4632 27494 4644
rect 29641 4641 29653 4644
rect 29687 4672 29699 4675
rect 30006 4672 30012 4684
rect 29687 4644 30012 4672
rect 29687 4641 29699 4644
rect 29641 4635 29699 4641
rect 30006 4632 30012 4644
rect 30064 4632 30070 4684
rect 32214 4632 32220 4684
rect 32272 4632 32278 4684
rect 27709 4607 27767 4613
rect 27709 4604 27721 4607
rect 26016 4576 27016 4604
rect 27080 4576 27721 4604
rect 26016 4564 26022 4576
rect 11900 4468 11928 4564
rect 27080 4480 27108 4576
rect 27709 4573 27721 4576
rect 27755 4573 27767 4607
rect 27709 4567 27767 4573
rect 28902 4564 28908 4616
rect 28960 4604 28966 4616
rect 29181 4607 29239 4613
rect 29181 4604 29193 4607
rect 28960 4576 29193 4604
rect 28960 4564 28966 4576
rect 29181 4573 29193 4576
rect 29227 4573 29239 4607
rect 29181 4567 29239 4573
rect 30101 4607 30159 4613
rect 30101 4573 30113 4607
rect 30147 4604 30159 4607
rect 30742 4604 30748 4616
rect 30147 4576 30748 4604
rect 30147 4573 30159 4576
rect 30101 4567 30159 4573
rect 30742 4564 30748 4576
rect 30800 4564 30806 4616
rect 33413 4607 33471 4613
rect 33413 4573 33425 4607
rect 33459 4604 33471 4607
rect 34698 4604 34704 4616
rect 33459 4576 34704 4604
rect 33459 4573 33471 4576
rect 33413 4567 33471 4573
rect 34698 4564 34704 4576
rect 34756 4564 34762 4616
rect 28718 4496 28724 4548
rect 28776 4536 28782 4548
rect 29917 4539 29975 4545
rect 29917 4536 29929 4539
rect 28776 4508 29929 4536
rect 28776 4496 28782 4508
rect 29917 4505 29929 4508
rect 29963 4505 29975 4539
rect 29917 4499 29975 4505
rect 8496 4440 11928 4468
rect 15194 4428 15200 4480
rect 15252 4428 15258 4480
rect 17773 4471 17831 4477
rect 17773 4437 17785 4471
rect 17819 4468 17831 4471
rect 17954 4468 17960 4480
rect 17819 4440 17960 4468
rect 17819 4437 17831 4440
rect 17773 4431 17831 4437
rect 17954 4428 17960 4440
rect 18012 4468 18018 4480
rect 19334 4468 19340 4480
rect 18012 4440 19340 4468
rect 18012 4428 18018 4440
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 20441 4471 20499 4477
rect 20441 4437 20453 4471
rect 20487 4468 20499 4471
rect 21174 4468 21180 4480
rect 20487 4440 21180 4468
rect 20487 4437 20499 4440
rect 20441 4431 20499 4437
rect 21174 4428 21180 4440
rect 21232 4428 21238 4480
rect 23477 4471 23535 4477
rect 23477 4437 23489 4471
rect 23523 4468 23535 4471
rect 23658 4468 23664 4480
rect 23523 4440 23664 4468
rect 23523 4437 23535 4440
rect 23477 4431 23535 4437
rect 23658 4428 23664 4440
rect 23716 4428 23722 4480
rect 27062 4428 27068 4480
rect 27120 4428 27126 4480
rect 29546 4428 29552 4480
rect 29604 4428 29610 4480
rect 2760 4378 34316 4400
rect 2760 4326 6550 4378
rect 6602 4326 6614 4378
rect 6666 4326 6678 4378
rect 6730 4326 6742 4378
rect 6794 4326 6806 4378
rect 6858 4326 14439 4378
rect 14491 4326 14503 4378
rect 14555 4326 14567 4378
rect 14619 4326 14631 4378
rect 14683 4326 14695 4378
rect 14747 4326 22328 4378
rect 22380 4326 22392 4378
rect 22444 4326 22456 4378
rect 22508 4326 22520 4378
rect 22572 4326 22584 4378
rect 22636 4326 30217 4378
rect 30269 4326 30281 4378
rect 30333 4326 30345 4378
rect 30397 4326 30409 4378
rect 30461 4326 30473 4378
rect 30525 4326 34316 4378
rect 2760 4304 34316 4326
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 5169 4267 5227 4273
rect 5169 4264 5181 4267
rect 4856 4236 5181 4264
rect 4856 4224 4862 4236
rect 5169 4233 5181 4236
rect 5215 4233 5227 4267
rect 5169 4227 5227 4233
rect 5534 4224 5540 4276
rect 5592 4264 5598 4276
rect 5721 4267 5779 4273
rect 5721 4264 5733 4267
rect 5592 4236 5733 4264
rect 5592 4224 5598 4236
rect 5721 4233 5733 4236
rect 5767 4233 5779 4267
rect 5721 4227 5779 4233
rect 6086 4224 6092 4276
rect 6144 4224 6150 4276
rect 6270 4224 6276 4276
rect 6328 4264 6334 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6328 4236 6837 4264
rect 6328 4224 6334 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 6825 4227 6883 4233
rect 8478 4224 8484 4276
rect 8536 4224 8542 4276
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 9548 4236 9597 4264
rect 9548 4224 9554 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 9585 4227 9643 4233
rect 13630 4224 13636 4276
rect 13688 4264 13694 4276
rect 13725 4267 13783 4273
rect 13725 4264 13737 4267
rect 13688 4236 13737 4264
rect 13688 4224 13694 4236
rect 13725 4233 13737 4236
rect 13771 4233 13783 4267
rect 13725 4227 13783 4233
rect 15286 4224 15292 4276
rect 15344 4224 15350 4276
rect 16209 4267 16267 4273
rect 16209 4233 16221 4267
rect 16255 4264 16267 4267
rect 16850 4264 16856 4276
rect 16255 4236 16856 4264
rect 16255 4233 16267 4236
rect 16209 4227 16267 4233
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 18417 4267 18475 4273
rect 18417 4233 18429 4267
rect 18463 4264 18475 4267
rect 18598 4264 18604 4276
rect 18463 4236 18604 4264
rect 18463 4233 18475 4236
rect 18417 4227 18475 4233
rect 18598 4224 18604 4236
rect 18656 4224 18662 4276
rect 24857 4267 24915 4273
rect 24857 4233 24869 4267
rect 24903 4264 24915 4267
rect 24946 4264 24952 4276
rect 24903 4236 24952 4264
rect 24903 4233 24915 4236
rect 24857 4227 24915 4233
rect 24946 4224 24952 4236
rect 25004 4224 25010 4276
rect 25590 4224 25596 4276
rect 25648 4264 25654 4276
rect 26053 4267 26111 4273
rect 26053 4264 26065 4267
rect 25648 4236 26065 4264
rect 25648 4224 25654 4236
rect 26053 4233 26065 4236
rect 26099 4233 26111 4267
rect 26053 4227 26111 4233
rect 26878 4224 26884 4276
rect 26936 4224 26942 4276
rect 28442 4264 28448 4276
rect 27724 4236 28448 4264
rect 4522 4088 4528 4140
rect 4580 4088 4586 4140
rect 5552 4128 5580 4224
rect 5626 4156 5632 4208
rect 5684 4196 5690 4208
rect 6549 4199 6607 4205
rect 6549 4196 6561 4199
rect 5684 4168 6561 4196
rect 5684 4156 5690 4168
rect 6549 4165 6561 4168
rect 6595 4196 6607 4199
rect 8496 4196 8524 4224
rect 16485 4199 16543 4205
rect 16485 4196 16497 4199
rect 6595 4168 8524 4196
rect 14752 4168 16497 4196
rect 6595 4165 6607 4168
rect 6549 4159 6607 4165
rect 6362 4128 6368 4140
rect 5552 4100 6368 4128
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 8297 4131 8355 4137
rect 8297 4097 8309 4131
rect 8343 4097 8355 4131
rect 8297 4091 8355 4097
rect 4430 4020 4436 4072
rect 4488 4020 4494 4072
rect 8312 4060 8340 4091
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 9030 4128 9036 4140
rect 8680 4100 9036 4128
rect 8481 4063 8539 4069
rect 8312 4032 8432 4060
rect 14 3952 20 4004
rect 72 3992 78 4004
rect 3237 3995 3295 4001
rect 3237 3992 3249 3995
rect 72 3964 3249 3992
rect 72 3952 78 3964
rect 3237 3961 3249 3964
rect 3283 3961 3295 3995
rect 8404 3992 8432 4032
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8570 4060 8576 4072
rect 8527 4032 8576 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 8680 3992 8708 4100
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 12584 4100 13185 4128
rect 12584 4088 12590 4100
rect 13173 4097 13185 4100
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 13722 4088 13728 4140
rect 13780 4128 13786 4140
rect 14277 4131 14335 4137
rect 14277 4128 14289 4131
rect 13780 4100 14289 4128
rect 13780 4088 13786 4100
rect 14277 4097 14289 4100
rect 14323 4128 14335 4131
rect 14642 4128 14648 4140
rect 14323 4100 14648 4128
rect 14323 4097 14335 4100
rect 14277 4091 14335 4097
rect 14642 4088 14648 4100
rect 14700 4128 14706 4140
rect 14752 4137 14780 4168
rect 16485 4165 16497 4168
rect 16531 4196 16543 4199
rect 18233 4199 18291 4205
rect 18233 4196 18245 4199
rect 16531 4168 18245 4196
rect 16531 4165 16543 4168
rect 16485 4159 16543 4165
rect 18233 4165 18245 4168
rect 18279 4165 18291 4199
rect 18233 4159 18291 4165
rect 19306 4168 20760 4196
rect 14737 4131 14795 4137
rect 14737 4128 14749 4131
rect 14700 4100 14749 4128
rect 14700 4088 14706 4100
rect 14737 4097 14749 4100
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 18248 4128 18276 4159
rect 18690 4128 18696 4140
rect 18248 4100 18696 4128
rect 18690 4088 18696 4100
rect 18748 4128 18754 4140
rect 18969 4131 19027 4137
rect 18969 4128 18981 4131
rect 18748 4100 18981 4128
rect 18748 4088 18754 4100
rect 18969 4097 18981 4100
rect 19015 4128 19027 4131
rect 19306 4128 19334 4168
rect 19015 4100 19334 4128
rect 19015 4097 19027 4100
rect 18969 4091 19027 4097
rect 20070 4088 20076 4140
rect 20128 4088 20134 4140
rect 20732 4137 20760 4168
rect 21100 4168 23336 4196
rect 21100 4137 21128 4168
rect 20717 4131 20775 4137
rect 20717 4097 20729 4131
rect 20763 4128 20775 4131
rect 21085 4131 21143 4137
rect 21085 4128 21097 4131
rect 20763 4100 21097 4128
rect 20763 4097 20775 4100
rect 20717 4091 20775 4097
rect 21085 4097 21097 4100
rect 21131 4097 21143 4131
rect 21085 4091 21143 4097
rect 21174 4088 21180 4140
rect 21232 4088 21238 4140
rect 23308 4137 23336 4168
rect 23293 4131 23351 4137
rect 23293 4097 23305 4131
rect 23339 4128 23351 4131
rect 23569 4131 23627 4137
rect 23569 4128 23581 4131
rect 23339 4100 23581 4128
rect 23339 4097 23351 4100
rect 23293 4091 23351 4097
rect 23569 4097 23581 4100
rect 23615 4128 23627 4131
rect 23615 4100 24348 4128
rect 23615 4097 23627 4100
rect 23569 4091 23627 4097
rect 8941 4063 8999 4069
rect 8941 4060 8953 4063
rect 8404 3964 8708 3992
rect 8864 4032 8953 4060
rect 3237 3955 3295 3961
rect 8864 3933 8892 4032
rect 8941 4029 8953 4032
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14093 4063 14151 4069
rect 14093 4060 14105 4063
rect 14056 4032 14105 4060
rect 14056 4020 14062 4032
rect 14093 4029 14105 4032
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 14185 4063 14243 4069
rect 14185 4029 14197 4063
rect 14231 4060 14243 4063
rect 15212 4060 15240 4088
rect 14231 4032 15240 4060
rect 15381 4063 15439 4069
rect 14231 4029 14243 4032
rect 14185 4023 14243 4029
rect 15381 4029 15393 4063
rect 15427 4029 15439 4063
rect 15381 4023 15439 4029
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 15396 3992 15424 4023
rect 18230 4020 18236 4072
rect 18288 4060 18294 4072
rect 18785 4063 18843 4069
rect 18785 4060 18797 4063
rect 18288 4032 18797 4060
rect 18288 4020 18294 4032
rect 18785 4029 18797 4032
rect 18831 4029 18843 4063
rect 18785 4023 18843 4029
rect 21269 4063 21327 4069
rect 21269 4029 21281 4063
rect 21315 4060 21327 4063
rect 21726 4060 21732 4072
rect 21315 4032 21732 4060
rect 21315 4029 21327 4032
rect 21269 4023 21327 4029
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 23750 4020 23756 4072
rect 23808 4020 23814 4072
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 24136 4032 24225 4060
rect 14884 3964 15424 3992
rect 14884 3952 14890 3964
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3893 8907 3927
rect 8849 3887 8907 3893
rect 18877 3927 18935 3933
rect 18877 3893 18889 3927
rect 18923 3924 18935 3927
rect 19521 3927 19579 3933
rect 19521 3924 19533 3927
rect 18923 3896 19533 3924
rect 18923 3893 18935 3896
rect 18877 3887 18935 3893
rect 19521 3893 19533 3896
rect 19567 3893 19579 3927
rect 19521 3887 19579 3893
rect 21637 3927 21695 3933
rect 21637 3893 21649 3927
rect 21683 3924 21695 3927
rect 22830 3924 22836 3936
rect 21683 3896 22836 3924
rect 21683 3893 21695 3896
rect 21637 3887 21695 3893
rect 22830 3884 22836 3896
rect 22888 3884 22894 3936
rect 23658 3884 23664 3936
rect 23716 3884 23722 3936
rect 24136 3933 24164 4032
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 24121 3927 24179 3933
rect 24121 3893 24133 3927
rect 24167 3893 24179 3927
rect 24320 3924 24348 4100
rect 25498 4088 25504 4140
rect 25556 4088 25562 4140
rect 26602 4088 26608 4140
rect 26660 4088 26666 4140
rect 27724 4137 27752 4236
rect 28442 4224 28448 4236
rect 28500 4224 28506 4276
rect 29457 4267 29515 4273
rect 29457 4233 29469 4267
rect 29503 4264 29515 4267
rect 29822 4264 29828 4276
rect 29503 4236 29828 4264
rect 29503 4233 29515 4236
rect 29457 4227 29515 4233
rect 29822 4224 29828 4236
rect 29880 4224 29886 4276
rect 27709 4131 27767 4137
rect 27709 4097 27721 4131
rect 27755 4097 27767 4131
rect 27709 4091 27767 4097
rect 27985 4131 28043 4137
rect 27985 4097 27997 4131
rect 28031 4128 28043 4131
rect 28534 4128 28540 4140
rect 28031 4100 28540 4128
rect 28031 4097 28043 4100
rect 27985 4091 28043 4097
rect 28534 4088 28540 4100
rect 28592 4088 28598 4140
rect 28718 4088 28724 4140
rect 28776 4128 28782 4140
rect 28776 4100 33640 4128
rect 28776 4088 28782 4100
rect 26973 4063 27031 4069
rect 26973 4029 26985 4063
rect 27019 4060 27031 4063
rect 27430 4060 27436 4072
rect 27019 4032 27436 4060
rect 27019 4029 27031 4032
rect 26973 4023 27031 4029
rect 27430 4020 27436 4032
rect 27488 4020 27494 4072
rect 29546 4060 29552 4072
rect 29118 4032 29552 4060
rect 29546 4020 29552 4032
rect 29604 4020 29610 4072
rect 31726 3964 33548 3992
rect 28902 3924 28908 3936
rect 24320 3896 28908 3924
rect 24121 3887 24179 3893
rect 28902 3884 28908 3896
rect 28960 3884 28966 3936
rect 28994 3884 29000 3936
rect 29052 3924 29058 3936
rect 31726 3924 31754 3964
rect 33520 3933 33548 3964
rect 29052 3896 31754 3924
rect 33505 3927 33563 3933
rect 29052 3884 29058 3896
rect 33505 3893 33517 3927
rect 33551 3893 33563 3927
rect 33612 3924 33640 4100
rect 33704 4100 34468 4128
rect 33704 4069 33732 4100
rect 34440 4072 34468 4100
rect 33689 4063 33747 4069
rect 33689 4029 33701 4063
rect 33735 4029 33747 4063
rect 33689 4023 33747 4029
rect 33962 4020 33968 4072
rect 34020 4020 34026 4072
rect 34422 4020 34428 4072
rect 34480 4020 34486 4072
rect 33781 3927 33839 3933
rect 33781 3924 33793 3927
rect 33612 3896 33793 3924
rect 33505 3887 33563 3893
rect 33781 3893 33793 3896
rect 33827 3893 33839 3927
rect 33781 3887 33839 3893
rect 2760 3834 34316 3856
rect 2760 3782 7210 3834
rect 7262 3782 7274 3834
rect 7326 3782 7338 3834
rect 7390 3782 7402 3834
rect 7454 3782 7466 3834
rect 7518 3782 15099 3834
rect 15151 3782 15163 3834
rect 15215 3782 15227 3834
rect 15279 3782 15291 3834
rect 15343 3782 15355 3834
rect 15407 3782 22988 3834
rect 23040 3782 23052 3834
rect 23104 3782 23116 3834
rect 23168 3782 23180 3834
rect 23232 3782 23244 3834
rect 23296 3782 30877 3834
rect 30929 3782 30941 3834
rect 30993 3782 31005 3834
rect 31057 3782 31069 3834
rect 31121 3782 31133 3834
rect 31185 3782 34316 3834
rect 2760 3760 34316 3782
rect 9030 3680 9036 3732
rect 9088 3680 9094 3732
rect 14642 3680 14648 3732
rect 14700 3680 14706 3732
rect 25866 3680 25872 3732
rect 25924 3680 25930 3732
rect 25958 3680 25964 3732
rect 26016 3680 26022 3732
rect 26786 3680 26792 3732
rect 26844 3720 26850 3732
rect 28718 3720 28724 3732
rect 26844 3692 28724 3720
rect 26844 3680 26850 3692
rect 28718 3680 28724 3692
rect 28776 3680 28782 3732
rect 28902 3680 28908 3732
rect 28960 3680 28966 3732
rect 1302 3612 1308 3664
rect 1360 3652 1366 3664
rect 3234 3652 3240 3664
rect 1360 3624 3240 3652
rect 1360 3612 1366 3624
rect 3234 3612 3240 3624
rect 3292 3612 3298 3664
rect 25884 3652 25912 3680
rect 28994 3652 29000 3664
rect 25884 3624 29000 3652
rect 28994 3612 29000 3624
rect 29052 3612 29058 3664
rect 4433 3587 4491 3593
rect 4433 3553 4445 3587
rect 4479 3584 4491 3587
rect 4890 3584 4896 3596
rect 4479 3556 4896 3584
rect 4479 3553 4491 3556
rect 4433 3547 4491 3553
rect 4890 3544 4896 3556
rect 4948 3544 4954 3596
rect 6641 3587 6699 3593
rect 6641 3553 6653 3587
rect 6687 3584 6699 3587
rect 8662 3584 8668 3596
rect 6687 3556 8668 3584
rect 6687 3553 6699 3556
rect 6641 3547 6699 3553
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 16390 3544 16396 3596
rect 16448 3544 16454 3596
rect 19334 3544 19340 3596
rect 19392 3584 19398 3596
rect 20717 3587 20775 3593
rect 20717 3584 20729 3587
rect 19392 3556 20729 3584
rect 19392 3544 19398 3556
rect 20717 3553 20729 3556
rect 20763 3553 20775 3587
rect 20717 3547 20775 3553
rect 32306 3544 32312 3596
rect 32364 3544 32370 3596
rect 33965 3587 34023 3593
rect 33965 3553 33977 3587
rect 34011 3584 34023 3587
rect 35434 3584 35440 3596
rect 34011 3556 35440 3584
rect 34011 3553 34023 3556
rect 33965 3547 34023 3553
rect 35434 3544 35440 3556
rect 35492 3544 35498 3596
rect 1302 3476 1308 3528
rect 1360 3516 1366 3528
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 1360 3488 3249 3516
rect 1360 3476 1366 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3237 3479 3295 3485
rect 5166 3476 5172 3528
rect 5224 3516 5230 3528
rect 5445 3519 5503 3525
rect 5445 3516 5457 3519
rect 5224 3488 5457 3516
rect 5224 3476 5230 3488
rect 5445 3485 5457 3488
rect 5491 3485 5503 3519
rect 5445 3479 5503 3485
rect 16114 3476 16120 3528
rect 16172 3516 16178 3528
rect 16669 3519 16727 3525
rect 16669 3516 16681 3519
rect 16172 3488 16681 3516
rect 16172 3476 16178 3488
rect 16669 3485 16681 3488
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 20622 3476 20628 3528
rect 20680 3516 20686 3528
rect 21177 3519 21235 3525
rect 21177 3516 21189 3519
rect 20680 3488 21189 3516
rect 20680 3476 20686 3488
rect 21177 3485 21189 3488
rect 21223 3485 21235 3519
rect 21177 3479 21235 3485
rect 21818 3476 21824 3528
rect 21876 3476 21882 3528
rect 33042 3476 33048 3528
rect 33100 3476 33106 3528
rect 13630 3408 13636 3460
rect 13688 3448 13694 3460
rect 21836 3448 21864 3476
rect 13688 3420 21864 3448
rect 13688 3408 13694 3420
rect 24394 3408 24400 3460
rect 24452 3448 24458 3460
rect 33781 3451 33839 3457
rect 33781 3448 33793 3451
rect 24452 3420 33793 3448
rect 24452 3408 24458 3420
rect 33781 3417 33793 3420
rect 33827 3417 33839 3451
rect 33781 3411 33839 3417
rect 9674 3340 9680 3392
rect 9732 3380 9738 3392
rect 18506 3380 18512 3392
rect 9732 3352 18512 3380
rect 9732 3340 9738 3352
rect 18506 3340 18512 3352
rect 18564 3340 18570 3392
rect 2760 3290 34316 3312
rect 2760 3238 6550 3290
rect 6602 3238 6614 3290
rect 6666 3238 6678 3290
rect 6730 3238 6742 3290
rect 6794 3238 6806 3290
rect 6858 3238 14439 3290
rect 14491 3238 14503 3290
rect 14555 3238 14567 3290
rect 14619 3238 14631 3290
rect 14683 3238 14695 3290
rect 14747 3238 22328 3290
rect 22380 3238 22392 3290
rect 22444 3238 22456 3290
rect 22508 3238 22520 3290
rect 22572 3238 22584 3290
rect 22636 3238 30217 3290
rect 30269 3238 30281 3290
rect 30333 3238 30345 3290
rect 30397 3238 30409 3290
rect 30461 3238 30473 3290
rect 30525 3238 34316 3290
rect 2760 3216 34316 3238
rect 9674 3136 9680 3188
rect 9732 3136 9738 3188
rect 11241 3179 11299 3185
rect 11241 3145 11253 3179
rect 11287 3176 11299 3179
rect 13630 3176 13636 3188
rect 11287 3148 13636 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 23661 3179 23719 3185
rect 23661 3145 23673 3179
rect 23707 3176 23719 3179
rect 24486 3176 24492 3188
rect 23707 3148 24492 3176
rect 23707 3145 23719 3148
rect 23661 3139 23719 3145
rect 24486 3136 24492 3148
rect 24544 3136 24550 3188
rect 25222 3136 25228 3188
rect 25280 3176 25286 3188
rect 26053 3179 26111 3185
rect 26053 3176 26065 3179
rect 25280 3148 26065 3176
rect 25280 3136 25286 3148
rect 26053 3145 26065 3148
rect 26099 3145 26111 3179
rect 26053 3139 26111 3145
rect 27614 3136 27620 3188
rect 27672 3176 27678 3188
rect 28629 3179 28687 3185
rect 28629 3176 28641 3179
rect 27672 3148 28641 3176
rect 27672 3136 27678 3148
rect 28629 3145 28641 3148
rect 28675 3145 28687 3179
rect 28629 3139 28687 3145
rect 31570 3136 31576 3188
rect 31628 3176 31634 3188
rect 31665 3179 31723 3185
rect 31665 3176 31677 3179
rect 31628 3148 31677 3176
rect 31628 3136 31634 3148
rect 31665 3145 31677 3148
rect 31711 3145 31723 3179
rect 31665 3139 31723 3145
rect 3237 3111 3295 3117
rect 3237 3077 3249 3111
rect 3283 3108 3295 3111
rect 13817 3111 13875 3117
rect 3283 3080 9674 3108
rect 3283 3077 3295 3080
rect 3237 3071 3295 3077
rect 2590 3000 2596 3052
rect 2648 3040 2654 3052
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 2648 3012 5457 3040
rect 2648 3000 2654 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 7800 3012 8493 3040
rect 7800 3000 7806 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 3050 2932 3056 2984
rect 3108 2932 3114 2984
rect 5258 2932 5264 2984
rect 5316 2932 5322 2984
rect 7837 2975 7895 2981
rect 7837 2941 7849 2975
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 4062 2864 4068 2916
rect 4120 2864 4126 2916
rect 6638 2864 6644 2916
rect 6696 2864 6702 2916
rect 7852 2904 7880 2935
rect 8018 2932 8024 2984
rect 8076 2932 8082 2984
rect 9030 2932 9036 2984
rect 9088 2972 9094 2984
rect 9493 2975 9551 2981
rect 9493 2972 9505 2975
rect 9088 2944 9505 2972
rect 9088 2932 9094 2944
rect 9493 2941 9505 2944
rect 9539 2941 9551 2975
rect 9493 2935 9551 2941
rect 9122 2904 9128 2916
rect 7852 2876 9128 2904
rect 9122 2864 9128 2876
rect 9180 2864 9186 2916
rect 9646 2836 9674 3080
rect 13817 3077 13829 3111
rect 13863 3108 13875 3111
rect 24302 3108 24308 3120
rect 13863 3080 24308 3108
rect 13863 3077 13875 3080
rect 13817 3071 13875 3077
rect 24302 3068 24308 3080
rect 24360 3068 24366 3120
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 17402 3000 17408 3052
rect 17460 3000 17466 3052
rect 18690 3000 18696 3052
rect 18748 3040 18754 3052
rect 19245 3043 19303 3049
rect 19245 3040 19257 3043
rect 18748 3012 19257 3040
rect 18748 3000 18754 3012
rect 19245 3009 19257 3012
rect 19291 3009 19303 3043
rect 19245 3003 19303 3009
rect 22002 3000 22008 3052
rect 22060 3040 22066 3052
rect 22373 3043 22431 3049
rect 22373 3040 22385 3043
rect 22060 3012 22385 3040
rect 22060 3000 22066 3012
rect 22373 3009 22385 3012
rect 22419 3009 22431 3043
rect 22373 3003 22431 3009
rect 24578 3000 24584 3052
rect 24636 3040 24642 3052
rect 24949 3043 25007 3049
rect 24949 3040 24961 3043
rect 24636 3012 24961 3040
rect 24636 3000 24642 3012
rect 24949 3009 24961 3012
rect 24995 3009 25007 3043
rect 24949 3003 25007 3009
rect 27154 3000 27160 3052
rect 27212 3040 27218 3052
rect 27525 3043 27583 3049
rect 27525 3040 27537 3043
rect 27212 3012 27537 3040
rect 27212 3000 27218 3012
rect 27525 3009 27537 3012
rect 27571 3009 27583 3043
rect 27525 3003 27583 3009
rect 29730 3000 29736 3052
rect 29788 3040 29794 3052
rect 30101 3043 30159 3049
rect 30101 3040 30113 3043
rect 29788 3012 30113 3040
rect 29788 3000 29794 3012
rect 30101 3009 30113 3012
rect 30147 3009 30159 3043
rect 30101 3003 30159 3009
rect 32858 3000 32864 3052
rect 32916 3000 32922 3052
rect 10962 2932 10968 2984
rect 11020 2972 11026 2984
rect 11057 2975 11115 2981
rect 11057 2972 11069 2975
rect 11020 2944 11069 2972
rect 11020 2932 11026 2944
rect 11057 2941 11069 2944
rect 11103 2941 11115 2975
rect 11057 2935 11115 2941
rect 12989 2975 13047 2981
rect 12989 2941 13001 2975
rect 13035 2972 13047 2975
rect 13262 2972 13268 2984
rect 13035 2944 13268 2972
rect 13035 2941 13047 2944
rect 12989 2935 13047 2941
rect 13262 2932 13268 2944
rect 13320 2932 13326 2984
rect 13630 2932 13636 2984
rect 13688 2932 13694 2984
rect 13906 2932 13912 2984
rect 13964 2972 13970 2984
rect 14185 2975 14243 2981
rect 14185 2972 14197 2975
rect 13964 2944 14197 2972
rect 13964 2932 13970 2944
rect 14185 2941 14197 2944
rect 14231 2941 14243 2975
rect 14185 2935 14243 2941
rect 16758 2932 16764 2984
rect 16816 2932 16822 2984
rect 18782 2932 18788 2984
rect 18840 2932 18846 2984
rect 21174 2932 21180 2984
rect 21232 2972 21238 2984
rect 21913 2975 21971 2981
rect 21913 2972 21925 2975
rect 21232 2944 21925 2972
rect 21232 2932 21238 2944
rect 21913 2941 21925 2944
rect 21959 2941 21971 2975
rect 21913 2935 21971 2941
rect 23382 2932 23388 2984
rect 23440 2972 23446 2984
rect 23477 2975 23535 2981
rect 23477 2972 23489 2975
rect 23440 2944 23489 2972
rect 23440 2932 23446 2944
rect 23477 2941 23489 2944
rect 23523 2941 23535 2975
rect 23477 2935 23535 2941
rect 23658 2932 23664 2984
rect 23716 2972 23722 2984
rect 24489 2975 24547 2981
rect 24489 2972 24501 2975
rect 23716 2944 24501 2972
rect 23716 2932 23722 2944
rect 24489 2941 24501 2944
rect 24535 2941 24547 2975
rect 24489 2935 24547 2941
rect 25774 2932 25780 2984
rect 25832 2972 25838 2984
rect 26237 2975 26295 2981
rect 26237 2972 26249 2975
rect 25832 2944 26249 2972
rect 25832 2932 25838 2944
rect 26237 2941 26249 2944
rect 26283 2941 26295 2975
rect 26237 2935 26295 2941
rect 27062 2932 27068 2984
rect 27120 2932 27126 2984
rect 28350 2932 28356 2984
rect 28408 2972 28414 2984
rect 28813 2975 28871 2981
rect 28813 2972 28825 2975
rect 28408 2944 28825 2972
rect 28408 2932 28414 2944
rect 28813 2941 28825 2944
rect 28859 2941 28871 2975
rect 28813 2935 28871 2941
rect 29822 2932 29828 2984
rect 29880 2932 29886 2984
rect 31570 2932 31576 2984
rect 31628 2972 31634 2984
rect 31849 2975 31907 2981
rect 31849 2972 31861 2975
rect 31628 2944 31861 2972
rect 31628 2932 31634 2944
rect 31849 2941 31861 2944
rect 31895 2941 31907 2975
rect 31849 2935 31907 2941
rect 31938 2932 31944 2984
rect 31996 2972 32002 2984
rect 32217 2975 32275 2981
rect 32217 2972 32229 2975
rect 31996 2944 32229 2972
rect 31996 2932 32002 2944
rect 32217 2941 32229 2944
rect 32263 2941 32275 2975
rect 32217 2935 32275 2941
rect 33965 2975 34023 2981
rect 33965 2941 33977 2975
rect 34011 2972 34023 2975
rect 36722 2972 36728 2984
rect 34011 2944 36728 2972
rect 34011 2941 34023 2944
rect 33965 2935 34023 2941
rect 36722 2932 36728 2944
rect 36780 2932 36786 2984
rect 21082 2864 21088 2916
rect 21140 2904 21146 2916
rect 21140 2876 33824 2904
rect 21140 2864 21146 2876
rect 25682 2836 25688 2848
rect 9646 2808 25688 2836
rect 25682 2796 25688 2808
rect 25740 2796 25746 2848
rect 33796 2845 33824 2876
rect 33781 2839 33839 2845
rect 33781 2805 33793 2839
rect 33827 2805 33839 2839
rect 33781 2799 33839 2805
rect 2760 2746 34316 2768
rect 2760 2694 7210 2746
rect 7262 2694 7274 2746
rect 7326 2694 7338 2746
rect 7390 2694 7402 2746
rect 7454 2694 7466 2746
rect 7518 2694 15099 2746
rect 15151 2694 15163 2746
rect 15215 2694 15227 2746
rect 15279 2694 15291 2746
rect 15343 2694 15355 2746
rect 15407 2694 22988 2746
rect 23040 2694 23052 2746
rect 23104 2694 23116 2746
rect 23168 2694 23180 2746
rect 23232 2694 23244 2746
rect 23296 2694 30877 2746
rect 30929 2694 30941 2746
rect 30993 2694 31005 2746
rect 31057 2694 31069 2746
rect 31121 2694 31133 2746
rect 31185 2694 34316 2746
rect 2760 2672 34316 2694
<< via1 >>
rect 7210 34246 7262 34298
rect 7274 34246 7326 34298
rect 7338 34246 7390 34298
rect 7402 34246 7454 34298
rect 7466 34246 7518 34298
rect 15099 34246 15151 34298
rect 15163 34246 15215 34298
rect 15227 34246 15279 34298
rect 15291 34246 15343 34298
rect 15355 34246 15407 34298
rect 22988 34246 23040 34298
rect 23052 34246 23104 34298
rect 23116 34246 23168 34298
rect 23180 34246 23232 34298
rect 23244 34246 23296 34298
rect 30877 34246 30929 34298
rect 30941 34246 30993 34298
rect 31005 34246 31057 34298
rect 31069 34246 31121 34298
rect 31133 34246 31185 34298
rect 7748 34144 7800 34196
rect 15476 34144 15528 34196
rect 22560 34144 22612 34196
rect 4528 34076 4580 34128
rect 5816 34076 5868 34128
rect 3056 34051 3108 34060
rect 3056 34017 3065 34051
rect 3065 34017 3099 34051
rect 3099 34017 3108 34051
rect 3056 34008 3108 34017
rect 4712 34008 4764 34060
rect 6000 34051 6052 34060
rect 6000 34017 6009 34051
rect 6009 34017 6043 34051
rect 6043 34017 6052 34051
rect 6000 34008 6052 34017
rect 12900 34076 12952 34128
rect 9128 34008 9180 34060
rect 9220 33940 9272 33992
rect 10324 34008 10376 34060
rect 10876 33983 10928 33992
rect 10876 33949 10885 33983
rect 10885 33949 10919 33983
rect 10919 33949 10928 33983
rect 10876 33940 10928 33949
rect 11704 33983 11756 33992
rect 11704 33949 11713 33983
rect 11713 33949 11747 33983
rect 11747 33949 11756 33983
rect 11704 33940 11756 33949
rect 10600 33872 10652 33924
rect 12624 34008 12676 34060
rect 13360 34051 13412 34060
rect 13360 34017 13369 34051
rect 13369 34017 13403 34051
rect 13403 34017 13412 34051
rect 13360 34008 13412 34017
rect 14188 34008 14240 34060
rect 19984 34076 20036 34128
rect 18420 34051 18472 34060
rect 18420 34017 18429 34051
rect 18429 34017 18463 34051
rect 18463 34017 18472 34051
rect 18420 34008 18472 34017
rect 22100 34051 22152 34060
rect 22100 34017 22109 34051
rect 22109 34017 22143 34051
rect 22143 34017 22152 34051
rect 22100 34008 22152 34017
rect 23848 34076 23900 34128
rect 28356 34076 28408 34128
rect 15200 33983 15252 33992
rect 15200 33949 15209 33983
rect 15209 33949 15243 33983
rect 15243 33949 15252 33983
rect 15200 33940 15252 33949
rect 17408 33940 17460 33992
rect 24124 34051 24176 34060
rect 24124 34017 24133 34051
rect 24133 34017 24167 34051
rect 24167 34017 24176 34051
rect 24124 34008 24176 34017
rect 26056 34051 26108 34060
rect 26056 34017 26065 34051
rect 26065 34017 26099 34051
rect 26099 34017 26108 34051
rect 26056 34008 26108 34017
rect 30012 34051 30064 34060
rect 30012 34017 30021 34051
rect 30021 34017 30055 34051
rect 30055 34017 30064 34051
rect 30012 34008 30064 34017
rect 31208 34051 31260 34060
rect 31208 34017 31217 34051
rect 31217 34017 31251 34051
rect 31251 34017 31260 34051
rect 31208 34008 31260 34017
rect 25136 33940 25188 33992
rect 29644 33940 29696 33992
rect 5540 33804 5592 33856
rect 8208 33847 8260 33856
rect 8208 33813 8217 33847
rect 8217 33813 8251 33847
rect 8251 33813 8260 33847
rect 8208 33804 8260 33813
rect 12256 33847 12308 33856
rect 12256 33813 12265 33847
rect 12265 33813 12299 33847
rect 12299 33813 12308 33847
rect 12256 33804 12308 33813
rect 12440 33847 12492 33856
rect 12440 33813 12449 33847
rect 12449 33813 12483 33847
rect 12483 33813 12492 33847
rect 12440 33804 12492 33813
rect 14188 33804 14240 33856
rect 15752 33804 15804 33856
rect 16948 33804 17000 33856
rect 22836 33847 22888 33856
rect 22836 33813 22845 33847
rect 22845 33813 22879 33847
rect 22879 33813 22888 33847
rect 22836 33804 22888 33813
rect 6550 33702 6602 33754
rect 6614 33702 6666 33754
rect 6678 33702 6730 33754
rect 6742 33702 6794 33754
rect 6806 33702 6858 33754
rect 14439 33702 14491 33754
rect 14503 33702 14555 33754
rect 14567 33702 14619 33754
rect 14631 33702 14683 33754
rect 14695 33702 14747 33754
rect 22328 33702 22380 33754
rect 22392 33702 22444 33754
rect 22456 33702 22508 33754
rect 22520 33702 22572 33754
rect 22584 33702 22636 33754
rect 30217 33702 30269 33754
rect 30281 33702 30333 33754
rect 30345 33702 30397 33754
rect 30409 33702 30461 33754
rect 30473 33702 30525 33754
rect 12624 33600 12676 33652
rect 3240 33464 3292 33516
rect 5908 33507 5960 33516
rect 5908 33473 5917 33507
rect 5917 33473 5951 33507
rect 5951 33473 5960 33507
rect 5908 33464 5960 33473
rect 12256 33464 12308 33516
rect 14188 33464 14240 33516
rect 5448 33439 5500 33448
rect 5448 33405 5457 33439
rect 5457 33405 5491 33439
rect 5491 33405 5500 33439
rect 5448 33396 5500 33405
rect 7932 33396 7984 33448
rect 10784 33439 10836 33448
rect 10784 33405 10793 33439
rect 10793 33405 10827 33439
rect 10827 33405 10836 33439
rect 10784 33396 10836 33405
rect 8944 33371 8996 33380
rect 8944 33337 8953 33371
rect 8953 33337 8987 33371
rect 8987 33337 8996 33371
rect 8944 33328 8996 33337
rect 12440 33328 12492 33380
rect 13084 33371 13136 33380
rect 13084 33337 13093 33371
rect 13093 33337 13127 33371
rect 13127 33337 13136 33371
rect 13084 33328 13136 33337
rect 13360 33328 13412 33380
rect 18696 33396 18748 33448
rect 19708 33464 19760 33516
rect 26424 33464 26476 33516
rect 33048 33600 33100 33652
rect 31300 33464 31352 33516
rect 14096 33328 14148 33380
rect 21272 33396 21324 33448
rect 26516 33439 26568 33448
rect 26516 33405 26525 33439
rect 26525 33405 26559 33439
rect 26559 33405 26568 33439
rect 26516 33396 26568 33405
rect 31392 33439 31444 33448
rect 31392 33405 31401 33439
rect 31401 33405 31435 33439
rect 31435 33405 31444 33439
rect 31392 33396 31444 33405
rect 32680 33328 32732 33380
rect 5172 33260 5224 33312
rect 11060 33260 11112 33312
rect 12532 33260 12584 33312
rect 15384 33260 15436 33312
rect 18604 33260 18656 33312
rect 19064 33303 19116 33312
rect 19064 33269 19073 33303
rect 19073 33269 19107 33303
rect 19107 33269 19116 33303
rect 19064 33260 19116 33269
rect 21548 33303 21600 33312
rect 21548 33269 21557 33303
rect 21557 33269 21591 33303
rect 21591 33269 21600 33303
rect 21548 33260 21600 33269
rect 7210 33158 7262 33210
rect 7274 33158 7326 33210
rect 7338 33158 7390 33210
rect 7402 33158 7454 33210
rect 7466 33158 7518 33210
rect 15099 33158 15151 33210
rect 15163 33158 15215 33210
rect 15227 33158 15279 33210
rect 15291 33158 15343 33210
rect 15355 33158 15407 33210
rect 22988 33158 23040 33210
rect 23052 33158 23104 33210
rect 23116 33158 23168 33210
rect 23180 33158 23232 33210
rect 23244 33158 23296 33210
rect 30877 33158 30929 33210
rect 30941 33158 30993 33210
rect 31005 33158 31057 33210
rect 31069 33158 31121 33210
rect 31133 33158 31185 33210
rect 1952 33056 2004 33108
rect 5908 33056 5960 33108
rect 8944 33056 8996 33108
rect 3240 33031 3292 33040
rect 3240 32997 3249 33031
rect 3249 32997 3283 33031
rect 3283 32997 3292 33031
rect 3240 32988 3292 32997
rect 3792 32988 3844 33040
rect 11428 33056 11480 33108
rect 11704 33056 11756 33108
rect 11888 33031 11940 33040
rect 11888 32997 11897 33031
rect 11897 32997 11931 33031
rect 11931 32997 11940 33031
rect 11888 32988 11940 32997
rect 5724 32963 5776 32972
rect 5724 32929 5733 32963
rect 5733 32929 5767 32963
rect 5767 32929 5776 32963
rect 5724 32920 5776 32929
rect 7288 32920 7340 32972
rect 10048 32963 10100 32972
rect 10048 32929 10057 32963
rect 10057 32929 10091 32963
rect 10091 32929 10100 32963
rect 10048 32920 10100 32929
rect 10968 32920 11020 32972
rect 11060 32920 11112 32972
rect 5356 32784 5408 32836
rect 10140 32852 10192 32904
rect 10600 32784 10652 32836
rect 11980 32963 12032 32972
rect 11980 32929 11989 32963
rect 11989 32929 12023 32963
rect 12023 32929 12032 32963
rect 11980 32920 12032 32929
rect 12164 32920 12216 32972
rect 12532 33056 12584 33108
rect 13820 33056 13872 33108
rect 15016 33056 15068 33108
rect 11704 32784 11756 32836
rect 12256 32895 12308 32904
rect 12256 32861 12265 32895
rect 12265 32861 12299 32895
rect 12299 32861 12308 32895
rect 12256 32852 12308 32861
rect 7288 32759 7340 32768
rect 7288 32725 7297 32759
rect 7297 32725 7331 32759
rect 7331 32725 7340 32759
rect 7288 32716 7340 32725
rect 11060 32716 11112 32768
rect 11152 32716 11204 32768
rect 14004 32963 14056 32972
rect 14004 32929 14010 32963
rect 14010 32929 14044 32963
rect 14044 32929 14056 32963
rect 14004 32920 14056 32929
rect 14096 32920 14148 32972
rect 14832 32920 14884 32972
rect 15108 32920 15160 32972
rect 15476 32963 15528 32972
rect 15476 32929 15485 32963
rect 15485 32929 15519 32963
rect 15519 32929 15528 32963
rect 15476 32920 15528 32929
rect 15568 32963 15620 32972
rect 15568 32929 15577 32963
rect 15577 32929 15611 32963
rect 15611 32929 15620 32963
rect 15568 32920 15620 32929
rect 16120 32895 16172 32904
rect 16120 32861 16129 32895
rect 16129 32861 16163 32895
rect 16163 32861 16172 32895
rect 16120 32852 16172 32861
rect 18880 32895 18932 32904
rect 18880 32861 18889 32895
rect 18889 32861 18923 32895
rect 18923 32861 18932 32895
rect 18880 32852 18932 32861
rect 14924 32784 14976 32836
rect 13728 32716 13780 32768
rect 14280 32716 14332 32768
rect 15016 32716 15068 32768
rect 29276 32963 29328 32972
rect 29276 32929 29285 32963
rect 29285 32929 29319 32963
rect 29319 32929 29328 32963
rect 29276 32920 29328 32929
rect 34796 32988 34848 33040
rect 36084 32988 36136 33040
rect 32312 32963 32364 32972
rect 32312 32929 32321 32963
rect 32321 32929 32355 32963
rect 32355 32929 32364 32963
rect 32312 32920 32364 32929
rect 16764 32759 16816 32768
rect 16764 32725 16773 32759
rect 16773 32725 16807 32759
rect 16807 32725 16816 32759
rect 16764 32716 16816 32725
rect 18328 32759 18380 32768
rect 18328 32725 18337 32759
rect 18337 32725 18371 32759
rect 18371 32725 18380 32759
rect 18328 32716 18380 32725
rect 32404 32852 32456 32904
rect 32220 32784 32272 32836
rect 19616 32716 19668 32768
rect 6550 32614 6602 32666
rect 6614 32614 6666 32666
rect 6678 32614 6730 32666
rect 6742 32614 6794 32666
rect 6806 32614 6858 32666
rect 14439 32614 14491 32666
rect 14503 32614 14555 32666
rect 14567 32614 14619 32666
rect 14631 32614 14683 32666
rect 14695 32614 14747 32666
rect 22328 32614 22380 32666
rect 22392 32614 22444 32666
rect 22456 32614 22508 32666
rect 22520 32614 22572 32666
rect 22584 32614 22636 32666
rect 30217 32614 30269 32666
rect 30281 32614 30333 32666
rect 30345 32614 30397 32666
rect 30409 32614 30461 32666
rect 30473 32614 30525 32666
rect 10048 32512 10100 32564
rect 11888 32512 11940 32564
rect 664 32376 716 32428
rect 7288 32444 7340 32496
rect 13268 32512 13320 32564
rect 13728 32512 13780 32564
rect 12808 32444 12860 32496
rect 13820 32444 13872 32496
rect 16120 32512 16172 32564
rect 16764 32512 16816 32564
rect 6000 32419 6052 32428
rect 6000 32385 6009 32419
rect 6009 32385 6043 32419
rect 6043 32385 6052 32419
rect 6000 32376 6052 32385
rect 6460 32376 6512 32428
rect 4436 32351 4488 32360
rect 4436 32317 4445 32351
rect 4445 32317 4479 32351
rect 4479 32317 4488 32351
rect 4436 32308 4488 32317
rect 8944 32351 8996 32360
rect 8944 32317 8953 32351
rect 8953 32317 8987 32351
rect 8987 32317 8996 32351
rect 8944 32308 8996 32317
rect 10784 32376 10836 32428
rect 12256 32419 12308 32428
rect 12256 32385 12265 32419
rect 12265 32385 12299 32419
rect 12299 32385 12308 32419
rect 12256 32376 12308 32385
rect 11704 32308 11756 32360
rect 11060 32240 11112 32292
rect 12348 32351 12400 32360
rect 12348 32317 12357 32351
rect 12357 32317 12391 32351
rect 12391 32317 12400 32351
rect 12348 32308 12400 32317
rect 12532 32351 12584 32360
rect 12532 32317 12541 32351
rect 12541 32317 12575 32351
rect 12575 32317 12584 32351
rect 12532 32308 12584 32317
rect 12808 32308 12860 32360
rect 5080 32172 5132 32224
rect 5908 32215 5960 32224
rect 5908 32181 5917 32215
rect 5917 32181 5951 32215
rect 5951 32181 5960 32215
rect 5908 32172 5960 32181
rect 8392 32215 8444 32224
rect 8392 32181 8401 32215
rect 8401 32181 8435 32215
rect 8435 32181 8444 32215
rect 8392 32172 8444 32181
rect 9312 32172 9364 32224
rect 11888 32215 11940 32224
rect 11888 32181 11897 32215
rect 11897 32181 11931 32215
rect 11931 32181 11940 32215
rect 11888 32172 11940 32181
rect 14832 32444 14884 32496
rect 15568 32444 15620 32496
rect 19616 32444 19668 32496
rect 26792 32512 26844 32564
rect 16580 32376 16632 32428
rect 18328 32376 18380 32428
rect 14372 32351 14424 32360
rect 14372 32317 14381 32351
rect 14381 32317 14415 32351
rect 14415 32317 14424 32351
rect 14372 32308 14424 32317
rect 14280 32283 14332 32292
rect 14280 32249 14289 32283
rect 14289 32249 14323 32283
rect 14323 32249 14332 32283
rect 14280 32240 14332 32249
rect 14832 32351 14884 32360
rect 14832 32317 14841 32351
rect 14841 32317 14875 32351
rect 14875 32317 14884 32351
rect 14832 32308 14884 32317
rect 14924 32308 14976 32360
rect 19708 32376 19760 32428
rect 19800 32376 19852 32428
rect 24492 32376 24544 32428
rect 13084 32172 13136 32224
rect 14096 32215 14148 32224
rect 14096 32181 14105 32215
rect 14105 32181 14139 32215
rect 14139 32181 14148 32215
rect 14096 32172 14148 32181
rect 14188 32172 14240 32224
rect 15660 32172 15712 32224
rect 15936 32240 15988 32292
rect 18604 32240 18656 32292
rect 30380 32376 30432 32428
rect 31208 32376 31260 32428
rect 34888 32376 34940 32428
rect 33048 32308 33100 32360
rect 18788 32172 18840 32224
rect 23848 32172 23900 32224
rect 24032 32215 24084 32224
rect 24032 32181 24041 32215
rect 24041 32181 24075 32215
rect 24075 32181 24084 32215
rect 24032 32172 24084 32181
rect 24860 32215 24912 32224
rect 24860 32181 24869 32215
rect 24869 32181 24903 32215
rect 24903 32181 24912 32215
rect 24860 32172 24912 32181
rect 25228 32172 25280 32224
rect 28264 32215 28316 32224
rect 28264 32181 28273 32215
rect 28273 32181 28307 32215
rect 28307 32181 28316 32215
rect 28264 32172 28316 32181
rect 28816 32215 28868 32224
rect 28816 32181 28825 32215
rect 28825 32181 28859 32215
rect 28859 32181 28868 32215
rect 28816 32172 28868 32181
rect 29184 32215 29236 32224
rect 29184 32181 29193 32215
rect 29193 32181 29227 32215
rect 29227 32181 29236 32215
rect 29184 32172 29236 32181
rect 7210 32070 7262 32122
rect 7274 32070 7326 32122
rect 7338 32070 7390 32122
rect 7402 32070 7454 32122
rect 7466 32070 7518 32122
rect 15099 32070 15151 32122
rect 15163 32070 15215 32122
rect 15227 32070 15279 32122
rect 15291 32070 15343 32122
rect 15355 32070 15407 32122
rect 22988 32070 23040 32122
rect 23052 32070 23104 32122
rect 23116 32070 23168 32122
rect 23180 32070 23232 32122
rect 23244 32070 23296 32122
rect 30877 32070 30929 32122
rect 30941 32070 30993 32122
rect 31005 32070 31057 32122
rect 31069 32070 31121 32122
rect 31133 32070 31185 32122
rect 5080 31900 5132 31952
rect 9220 31968 9272 32020
rect 10140 32011 10192 32020
rect 10140 31977 10149 32011
rect 10149 31977 10183 32011
rect 10183 31977 10192 32011
rect 10140 31968 10192 31977
rect 15476 31968 15528 32020
rect 15936 31968 15988 32020
rect 18880 31968 18932 32020
rect 8392 31900 8444 31952
rect 9312 31900 9364 31952
rect 11060 31943 11112 31952
rect 11060 31909 11095 31943
rect 11095 31909 11112 31943
rect 11060 31900 11112 31909
rect 11888 31900 11940 31952
rect 12256 31900 12308 31952
rect 12532 31900 12584 31952
rect 14096 31900 14148 31952
rect 4620 31832 4672 31884
rect 4896 31875 4948 31884
rect 4896 31841 4905 31875
rect 4905 31841 4939 31875
rect 4939 31841 4948 31875
rect 4896 31832 4948 31841
rect 6920 31875 6972 31884
rect 6920 31841 6929 31875
rect 6929 31841 6963 31875
rect 6963 31841 6972 31875
rect 6920 31832 6972 31841
rect 7932 31832 7984 31884
rect 10692 31832 10744 31884
rect 10876 31875 10928 31884
rect 10876 31841 10885 31875
rect 10885 31841 10919 31875
rect 10919 31841 10928 31875
rect 10876 31832 10928 31841
rect 10968 31875 11020 31884
rect 10968 31841 10977 31875
rect 10977 31841 11011 31875
rect 11011 31841 11020 31875
rect 10968 31832 11020 31841
rect 3240 31807 3292 31816
rect 3240 31773 3249 31807
rect 3249 31773 3283 31807
rect 3283 31773 3292 31807
rect 3240 31764 3292 31773
rect 6184 31764 6236 31816
rect 11704 31832 11756 31884
rect 12164 31832 12216 31884
rect 14832 31900 14884 31952
rect 15384 31943 15436 31952
rect 15384 31909 15393 31943
rect 15393 31909 15427 31943
rect 15427 31909 15436 31943
rect 15384 31900 15436 31909
rect 15568 31900 15620 31952
rect 18788 31943 18840 31952
rect 18788 31909 18797 31943
rect 18797 31909 18831 31943
rect 18831 31909 18840 31943
rect 18788 31900 18840 31909
rect 14280 31832 14332 31884
rect 19156 31832 19208 31884
rect 15752 31764 15804 31816
rect 16580 31764 16632 31816
rect 17776 31807 17828 31816
rect 17776 31773 17785 31807
rect 17785 31773 17819 31807
rect 17819 31773 17828 31807
rect 17776 31764 17828 31773
rect 19800 31968 19852 32020
rect 25228 32011 25280 32020
rect 25228 31977 25237 32011
rect 25237 31977 25271 32011
rect 25271 31977 25280 32011
rect 25228 31968 25280 31977
rect 26056 31968 26108 32020
rect 30380 32011 30432 32020
rect 30380 31977 30389 32011
rect 30389 31977 30423 32011
rect 30423 31977 30432 32011
rect 30380 31968 30432 31977
rect 24032 31900 24084 31952
rect 29184 31900 29236 31952
rect 31300 31900 31352 31952
rect 33508 31900 33560 31952
rect 24860 31832 24912 31884
rect 27620 31875 27672 31884
rect 27620 31841 27629 31875
rect 27629 31841 27663 31875
rect 27663 31841 27672 31875
rect 27620 31832 27672 31841
rect 28540 31832 28592 31884
rect 32220 31875 32272 31884
rect 32220 31841 32229 31875
rect 32229 31841 32263 31875
rect 32263 31841 32272 31875
rect 32220 31832 32272 31841
rect 11336 31696 11388 31748
rect 14372 31696 14424 31748
rect 10600 31671 10652 31680
rect 10600 31637 10609 31671
rect 10609 31637 10643 31671
rect 10643 31637 10652 31671
rect 10600 31628 10652 31637
rect 10876 31628 10928 31680
rect 11980 31628 12032 31680
rect 14924 31628 14976 31680
rect 17224 31671 17276 31680
rect 17224 31637 17233 31671
rect 17233 31637 17267 31671
rect 17267 31637 17276 31671
rect 17224 31628 17276 31637
rect 17868 31628 17920 31680
rect 27528 31696 27580 31748
rect 30564 31764 30616 31816
rect 31852 31807 31904 31816
rect 31852 31773 31861 31807
rect 31861 31773 31895 31807
rect 31895 31773 31904 31807
rect 31852 31764 31904 31773
rect 32128 31807 32180 31816
rect 32128 31773 32137 31807
rect 32137 31773 32171 31807
rect 32171 31773 32180 31807
rect 32128 31764 32180 31773
rect 23296 31628 23348 31680
rect 26516 31628 26568 31680
rect 26884 31628 26936 31680
rect 27804 31671 27856 31680
rect 27804 31637 27813 31671
rect 27813 31637 27847 31671
rect 27847 31637 27856 31671
rect 27804 31628 27856 31637
rect 6550 31526 6602 31578
rect 6614 31526 6666 31578
rect 6678 31526 6730 31578
rect 6742 31526 6794 31578
rect 6806 31526 6858 31578
rect 14439 31526 14491 31578
rect 14503 31526 14555 31578
rect 14567 31526 14619 31578
rect 14631 31526 14683 31578
rect 14695 31526 14747 31578
rect 22328 31526 22380 31578
rect 22392 31526 22444 31578
rect 22456 31526 22508 31578
rect 22520 31526 22572 31578
rect 22584 31526 22636 31578
rect 30217 31526 30269 31578
rect 30281 31526 30333 31578
rect 30345 31526 30397 31578
rect 30409 31526 30461 31578
rect 30473 31526 30525 31578
rect 5448 31424 5500 31476
rect 15384 31424 15436 31476
rect 15476 31467 15528 31476
rect 15476 31433 15485 31467
rect 15485 31433 15519 31467
rect 15519 31433 15528 31467
rect 15476 31424 15528 31433
rect 18420 31424 18472 31476
rect 26792 31424 26844 31476
rect 5080 31356 5132 31408
rect 4896 31288 4948 31340
rect 7012 31356 7064 31408
rect 10600 31288 10652 31340
rect 11980 31288 12032 31340
rect 16580 31331 16632 31340
rect 16580 31297 16589 31331
rect 16589 31297 16623 31331
rect 16623 31297 16632 31331
rect 16580 31288 16632 31297
rect 17224 31288 17276 31340
rect 18788 31331 18840 31340
rect 18788 31297 18797 31331
rect 18797 31297 18831 31331
rect 18831 31297 18840 31331
rect 18788 31288 18840 31297
rect 23296 31288 23348 31340
rect 26516 31331 26568 31340
rect 26516 31297 26525 31331
rect 26525 31297 26559 31331
rect 26559 31297 26568 31331
rect 26516 31288 26568 31297
rect 26884 31288 26936 31340
rect 3332 31195 3384 31204
rect 3332 31161 3341 31195
rect 3341 31161 3375 31195
rect 3375 31161 3384 31195
rect 3332 31152 3384 31161
rect 5540 31263 5592 31272
rect 5540 31229 5549 31263
rect 5549 31229 5583 31263
rect 5583 31229 5592 31263
rect 5540 31220 5592 31229
rect 6920 31220 6972 31272
rect 7840 31220 7892 31272
rect 10140 31220 10192 31272
rect 10968 31220 11020 31272
rect 4896 31084 4948 31136
rect 6368 31152 6420 31204
rect 11888 31195 11940 31204
rect 11888 31161 11897 31195
rect 11897 31161 11931 31195
rect 11931 31161 11940 31195
rect 11888 31152 11940 31161
rect 7932 31084 7984 31136
rect 9772 31127 9824 31136
rect 9772 31093 9781 31127
rect 9781 31093 9815 31127
rect 9815 31093 9824 31127
rect 9772 31084 9824 31093
rect 10324 31084 10376 31136
rect 11152 31084 11204 31136
rect 11336 31127 11388 31136
rect 11336 31093 11345 31127
rect 11345 31093 11379 31127
rect 11379 31093 11388 31127
rect 12164 31263 12216 31272
rect 12164 31229 12173 31263
rect 12173 31229 12207 31263
rect 12207 31229 12216 31263
rect 12164 31220 12216 31229
rect 16488 31263 16540 31272
rect 16488 31229 16497 31263
rect 16497 31229 16531 31263
rect 16531 31229 16540 31263
rect 16488 31220 16540 31229
rect 11336 31084 11388 31093
rect 12256 31127 12308 31136
rect 12256 31093 12265 31127
rect 12265 31093 12299 31127
rect 12299 31093 12308 31127
rect 12256 31084 12308 31093
rect 12440 31127 12492 31136
rect 12440 31093 12449 31127
rect 12449 31093 12483 31127
rect 12483 31093 12492 31127
rect 12440 31084 12492 31093
rect 13360 31084 13412 31136
rect 16580 31152 16632 31204
rect 18144 31152 18196 31204
rect 16304 31127 16356 31136
rect 16304 31093 16313 31127
rect 16313 31093 16347 31127
rect 16347 31093 16356 31127
rect 16304 31084 16356 31093
rect 23664 31220 23716 31272
rect 31300 31467 31352 31476
rect 31300 31433 31309 31467
rect 31309 31433 31343 31467
rect 31343 31433 31352 31467
rect 31300 31424 31352 31433
rect 30012 31331 30064 31340
rect 30012 31297 30021 31331
rect 30021 31297 30055 31331
rect 30055 31297 30064 31331
rect 30012 31288 30064 31297
rect 33784 31331 33836 31340
rect 33784 31297 33793 31331
rect 33793 31297 33827 31331
rect 33827 31297 33836 31331
rect 33784 31288 33836 31297
rect 30748 31263 30800 31272
rect 30748 31229 30757 31263
rect 30757 31229 30791 31263
rect 30791 31229 30800 31263
rect 30748 31220 30800 31229
rect 32496 31263 32548 31272
rect 32496 31229 32505 31263
rect 32505 31229 32539 31263
rect 32539 31229 32548 31263
rect 32496 31220 32548 31229
rect 32772 31263 32824 31272
rect 32772 31229 32781 31263
rect 32781 31229 32815 31263
rect 32815 31229 32824 31263
rect 32772 31220 32824 31229
rect 22560 31195 22612 31204
rect 22560 31161 22569 31195
rect 22569 31161 22603 31195
rect 22603 31161 22612 31195
rect 22560 31152 22612 31161
rect 27804 31152 27856 31204
rect 28724 31152 28776 31204
rect 31576 31152 31628 31204
rect 32036 31152 32088 31204
rect 24124 31084 24176 31136
rect 24768 31084 24820 31136
rect 28540 31084 28592 31136
rect 30196 31127 30248 31136
rect 30196 31093 30205 31127
rect 30205 31093 30239 31127
rect 30239 31093 30248 31127
rect 30196 31084 30248 31093
rect 31852 31127 31904 31136
rect 31852 31093 31861 31127
rect 31861 31093 31895 31127
rect 31895 31093 31904 31127
rect 31852 31084 31904 31093
rect 7210 30982 7262 31034
rect 7274 30982 7326 31034
rect 7338 30982 7390 31034
rect 7402 30982 7454 31034
rect 7466 30982 7518 31034
rect 15099 30982 15151 31034
rect 15163 30982 15215 31034
rect 15227 30982 15279 31034
rect 15291 30982 15343 31034
rect 15355 30982 15407 31034
rect 22988 30982 23040 31034
rect 23052 30982 23104 31034
rect 23116 30982 23168 31034
rect 23180 30982 23232 31034
rect 23244 30982 23296 31034
rect 30877 30982 30929 31034
rect 30941 30982 30993 31034
rect 31005 30982 31057 31034
rect 31069 30982 31121 31034
rect 31133 30982 31185 31034
rect 4896 30880 4948 30932
rect 6368 30923 6420 30932
rect 6368 30889 6377 30923
rect 6377 30889 6411 30923
rect 6411 30889 6420 30923
rect 6368 30880 6420 30889
rect 8944 30880 8996 30932
rect 4712 30855 4764 30864
rect 4712 30821 4721 30855
rect 4721 30821 4755 30855
rect 4755 30821 4764 30855
rect 4712 30812 4764 30821
rect 5356 30812 5408 30864
rect 9220 30880 9272 30932
rect 9772 30880 9824 30932
rect 11704 30923 11756 30932
rect 11704 30889 11713 30923
rect 11713 30889 11747 30923
rect 11747 30889 11756 30923
rect 11704 30880 11756 30889
rect 12440 30880 12492 30932
rect 12624 30880 12676 30932
rect 13360 30880 13412 30932
rect 16488 30880 16540 30932
rect 17776 30880 17828 30932
rect 18420 30880 18472 30932
rect 18788 30880 18840 30932
rect 22560 30880 22612 30932
rect 27528 30880 27580 30932
rect 28540 30880 28592 30932
rect 8300 30787 8352 30796
rect 8300 30753 8309 30787
rect 8309 30753 8343 30787
rect 8343 30753 8352 30787
rect 8300 30744 8352 30753
rect 5264 30719 5316 30728
rect 5264 30685 5273 30719
rect 5273 30685 5307 30719
rect 5307 30685 5316 30719
rect 5264 30676 5316 30685
rect 9220 30787 9272 30796
rect 9220 30753 9229 30787
rect 9229 30753 9263 30787
rect 9263 30753 9272 30787
rect 9220 30744 9272 30753
rect 10784 30744 10836 30796
rect 11888 30812 11940 30864
rect 12256 30744 12308 30796
rect 12440 30744 12492 30796
rect 12624 30787 12676 30796
rect 12624 30753 12633 30787
rect 12633 30753 12667 30787
rect 12667 30753 12676 30787
rect 12624 30744 12676 30753
rect 4160 30540 4212 30592
rect 5816 30583 5868 30592
rect 5816 30549 5825 30583
rect 5825 30549 5859 30583
rect 5859 30549 5868 30583
rect 5816 30540 5868 30549
rect 8208 30583 8260 30592
rect 8208 30549 8217 30583
rect 8217 30549 8251 30583
rect 8251 30549 8260 30583
rect 8208 30540 8260 30549
rect 10692 30608 10744 30660
rect 12716 30719 12768 30728
rect 12716 30685 12725 30719
rect 12725 30685 12759 30719
rect 12759 30685 12768 30719
rect 12716 30676 12768 30685
rect 14188 30744 14240 30796
rect 16580 30744 16632 30796
rect 17684 30787 17736 30796
rect 17684 30753 17693 30787
rect 17693 30753 17727 30787
rect 17727 30753 17736 30787
rect 17684 30744 17736 30753
rect 30196 30880 30248 30932
rect 31576 30880 31628 30932
rect 15108 30719 15160 30728
rect 15108 30685 15117 30719
rect 15117 30685 15151 30719
rect 15151 30685 15160 30719
rect 15108 30676 15160 30685
rect 17868 30719 17920 30728
rect 14832 30608 14884 30660
rect 9588 30540 9640 30592
rect 9680 30540 9732 30592
rect 10784 30540 10836 30592
rect 11152 30540 11204 30592
rect 11980 30540 12032 30592
rect 12256 30583 12308 30592
rect 12256 30549 12265 30583
rect 12265 30549 12299 30583
rect 12299 30549 12308 30583
rect 12256 30540 12308 30549
rect 13268 30583 13320 30592
rect 13268 30549 13277 30583
rect 13277 30549 13311 30583
rect 13311 30549 13320 30583
rect 13268 30540 13320 30549
rect 14188 30540 14240 30592
rect 17868 30685 17877 30719
rect 17877 30685 17911 30719
rect 17911 30685 17920 30719
rect 17868 30676 17920 30685
rect 18144 30676 18196 30728
rect 17224 30540 17276 30592
rect 17868 30540 17920 30592
rect 24768 30787 24820 30796
rect 24768 30753 24777 30787
rect 24777 30753 24811 30787
rect 24811 30753 24820 30787
rect 24768 30744 24820 30753
rect 27804 30744 27856 30796
rect 31392 30787 31444 30796
rect 19708 30719 19760 30728
rect 19708 30685 19717 30719
rect 19717 30685 19751 30719
rect 19751 30685 19760 30719
rect 19708 30676 19760 30685
rect 24032 30719 24084 30728
rect 24032 30685 24041 30719
rect 24041 30685 24075 30719
rect 24075 30685 24084 30719
rect 24032 30676 24084 30685
rect 25504 30719 25556 30728
rect 25504 30685 25513 30719
rect 25513 30685 25547 30719
rect 25547 30685 25556 30719
rect 25504 30676 25556 30685
rect 19156 30583 19208 30592
rect 19156 30549 19165 30583
rect 19165 30549 19199 30583
rect 19199 30549 19208 30583
rect 19156 30540 19208 30549
rect 23480 30540 23532 30592
rect 24952 30583 25004 30592
rect 24952 30549 24961 30583
rect 24961 30549 24995 30583
rect 24995 30549 25004 30583
rect 24952 30540 25004 30549
rect 26240 30540 26292 30592
rect 28264 30676 28316 30728
rect 31392 30753 31401 30787
rect 31401 30753 31435 30787
rect 31435 30753 31444 30787
rect 31392 30744 31444 30753
rect 31852 30880 31904 30932
rect 33048 30880 33100 30932
rect 27620 30540 27672 30592
rect 29092 30540 29144 30592
rect 30840 30583 30892 30592
rect 30840 30549 30849 30583
rect 30849 30549 30883 30583
rect 30883 30549 30892 30583
rect 30840 30540 30892 30549
rect 31208 30540 31260 30592
rect 31392 30540 31444 30592
rect 31576 30540 31628 30592
rect 6550 30438 6602 30490
rect 6614 30438 6666 30490
rect 6678 30438 6730 30490
rect 6742 30438 6794 30490
rect 6806 30438 6858 30490
rect 14439 30438 14491 30490
rect 14503 30438 14555 30490
rect 14567 30438 14619 30490
rect 14631 30438 14683 30490
rect 14695 30438 14747 30490
rect 22328 30438 22380 30490
rect 22392 30438 22444 30490
rect 22456 30438 22508 30490
rect 22520 30438 22572 30490
rect 22584 30438 22636 30490
rect 30217 30438 30269 30490
rect 30281 30438 30333 30490
rect 30345 30438 30397 30490
rect 30409 30438 30461 30490
rect 30473 30438 30525 30490
rect 3332 30336 3384 30388
rect 5264 30336 5316 30388
rect 10324 30336 10376 30388
rect 14188 30336 14240 30388
rect 15108 30336 15160 30388
rect 24032 30336 24084 30388
rect 30748 30336 30800 30388
rect 32772 30336 32824 30388
rect 5448 30200 5500 30252
rect 4160 30175 4212 30184
rect 4160 30141 4169 30175
rect 4169 30141 4203 30175
rect 4203 30141 4212 30175
rect 6000 30200 6052 30252
rect 6368 30200 6420 30252
rect 4160 30132 4212 30141
rect 7012 30200 7064 30252
rect 7932 30243 7984 30252
rect 7932 30209 7941 30243
rect 7941 30209 7975 30243
rect 7975 30209 7984 30243
rect 7932 30200 7984 30209
rect 9220 30200 9272 30252
rect 12256 30243 12308 30252
rect 12256 30209 12265 30243
rect 12265 30209 12299 30243
rect 12299 30209 12308 30243
rect 12256 30200 12308 30209
rect 15660 30200 15712 30252
rect 23480 30268 23532 30320
rect 23664 30268 23716 30320
rect 25780 30268 25832 30320
rect 6828 30132 6880 30184
rect 7196 30175 7248 30184
rect 7196 30141 7205 30175
rect 7205 30141 7239 30175
rect 7239 30141 7248 30175
rect 7196 30132 7248 30141
rect 1308 30064 1360 30116
rect 5724 30064 5776 30116
rect 3240 30039 3292 30048
rect 3240 30005 3249 30039
rect 3249 30005 3283 30039
rect 3283 30005 3292 30039
rect 3240 29996 3292 30005
rect 8208 30107 8260 30116
rect 8208 30073 8217 30107
rect 8217 30073 8251 30107
rect 8251 30073 8260 30107
rect 8208 30064 8260 30073
rect 8852 30064 8904 30116
rect 13268 30132 13320 30184
rect 16028 30132 16080 30184
rect 16304 30132 16356 30184
rect 16856 30175 16908 30184
rect 16856 30141 16865 30175
rect 16865 30141 16899 30175
rect 16899 30141 16908 30175
rect 16856 30132 16908 30141
rect 14096 30064 14148 30116
rect 23388 30200 23440 30252
rect 24032 30243 24084 30252
rect 24032 30209 24041 30243
rect 24041 30209 24075 30243
rect 24075 30209 24084 30243
rect 24032 30200 24084 30209
rect 24952 30200 25004 30252
rect 25044 30200 25096 30252
rect 26792 30200 26844 30252
rect 7932 29996 7984 30048
rect 9680 30039 9732 30048
rect 9680 30005 9689 30039
rect 9689 30005 9723 30039
rect 9723 30005 9732 30039
rect 9680 29996 9732 30005
rect 9772 29996 9824 30048
rect 10140 30039 10192 30048
rect 10140 30005 10149 30039
rect 10149 30005 10183 30039
rect 10183 30005 10192 30039
rect 10140 29996 10192 30005
rect 10968 29996 11020 30048
rect 12256 29996 12308 30048
rect 12900 29996 12952 30048
rect 12992 29996 13044 30048
rect 16212 29996 16264 30048
rect 23388 29996 23440 30048
rect 23572 29996 23624 30048
rect 26700 30132 26752 30184
rect 28540 30175 28592 30184
rect 28540 30141 28549 30175
rect 28549 30141 28583 30175
rect 28583 30141 28592 30175
rect 28540 30132 28592 30141
rect 29368 30175 29420 30184
rect 29368 30141 29377 30175
rect 29377 30141 29411 30175
rect 29411 30141 29420 30175
rect 29368 30132 29420 30141
rect 30840 30200 30892 30252
rect 30380 30132 30432 30184
rect 30472 30175 30524 30184
rect 30472 30141 30481 30175
rect 30481 30141 30515 30175
rect 30515 30141 30524 30175
rect 30472 30132 30524 30141
rect 30656 30132 30708 30184
rect 31208 30175 31260 30184
rect 31208 30141 31217 30175
rect 31217 30141 31251 30175
rect 31251 30141 31260 30175
rect 31208 30132 31260 30141
rect 25044 29996 25096 30048
rect 25228 29996 25280 30048
rect 26884 29996 26936 30048
rect 27620 29996 27672 30048
rect 27712 30039 27764 30048
rect 27712 30005 27721 30039
rect 27721 30005 27755 30039
rect 27755 30005 27764 30039
rect 27712 29996 27764 30005
rect 27988 29996 28040 30048
rect 28908 29996 28960 30048
rect 32220 30064 32272 30116
rect 35164 30132 35216 30184
rect 34060 30064 34112 30116
rect 32128 29996 32180 30048
rect 7210 29894 7262 29946
rect 7274 29894 7326 29946
rect 7338 29894 7390 29946
rect 7402 29894 7454 29946
rect 7466 29894 7518 29946
rect 15099 29894 15151 29946
rect 15163 29894 15215 29946
rect 15227 29894 15279 29946
rect 15291 29894 15343 29946
rect 15355 29894 15407 29946
rect 22988 29894 23040 29946
rect 23052 29894 23104 29946
rect 23116 29894 23168 29946
rect 23180 29894 23232 29946
rect 23244 29894 23296 29946
rect 30877 29894 30929 29946
rect 30941 29894 30993 29946
rect 31005 29894 31057 29946
rect 31069 29894 31121 29946
rect 31133 29894 31185 29946
rect 5724 29792 5776 29844
rect 5816 29792 5868 29844
rect 8852 29835 8904 29844
rect 8852 29801 8861 29835
rect 8861 29801 8895 29835
rect 8895 29801 8904 29835
rect 8852 29792 8904 29801
rect 9588 29792 9640 29844
rect 10324 29792 10376 29844
rect 11060 29792 11112 29844
rect 12624 29792 12676 29844
rect 13544 29792 13596 29844
rect 14096 29835 14148 29844
rect 14096 29801 14105 29835
rect 14105 29801 14139 29835
rect 14139 29801 14148 29835
rect 14096 29792 14148 29801
rect 14280 29792 14332 29844
rect 16028 29835 16080 29844
rect 16028 29801 16037 29835
rect 16037 29801 16071 29835
rect 16071 29801 16080 29835
rect 16028 29792 16080 29801
rect 16856 29792 16908 29844
rect 25228 29792 25280 29844
rect 25504 29792 25556 29844
rect 27804 29792 27856 29844
rect 28540 29792 28592 29844
rect 28908 29792 28960 29844
rect 30472 29792 30524 29844
rect 32496 29792 32548 29844
rect 33048 29792 33100 29844
rect 4712 29656 4764 29708
rect 7932 29656 7984 29708
rect 9680 29724 9732 29776
rect 10416 29699 10468 29708
rect 10416 29665 10425 29699
rect 10425 29665 10459 29699
rect 10459 29665 10468 29699
rect 10416 29656 10468 29665
rect 10508 29656 10560 29708
rect 10784 29656 10836 29708
rect 12716 29724 12768 29776
rect 12900 29724 12952 29776
rect 5632 29588 5684 29640
rect 6828 29588 6880 29640
rect 6920 29631 6972 29640
rect 6920 29597 6929 29631
rect 6929 29597 6963 29631
rect 6963 29597 6972 29631
rect 6920 29588 6972 29597
rect 7564 29588 7616 29640
rect 8300 29588 8352 29640
rect 9864 29631 9916 29640
rect 9864 29597 9873 29631
rect 9873 29597 9907 29631
rect 9907 29597 9916 29631
rect 9864 29588 9916 29597
rect 10968 29588 11020 29640
rect 12256 29699 12308 29708
rect 12256 29665 12265 29699
rect 12265 29665 12299 29699
rect 12299 29665 12308 29699
rect 12256 29656 12308 29665
rect 4988 29520 5040 29572
rect 12992 29631 13044 29640
rect 12992 29597 13001 29631
rect 13001 29597 13035 29631
rect 13035 29597 13044 29631
rect 12992 29588 13044 29597
rect 14832 29724 14884 29776
rect 13912 29656 13964 29708
rect 15016 29656 15068 29708
rect 15476 29656 15528 29708
rect 17592 29699 17644 29708
rect 17592 29665 17601 29699
rect 17601 29665 17635 29699
rect 17635 29665 17644 29699
rect 17592 29656 17644 29665
rect 26240 29724 26292 29776
rect 26884 29724 26936 29776
rect 25136 29656 25188 29708
rect 12072 29520 12124 29572
rect 12440 29520 12492 29572
rect 5448 29452 5500 29504
rect 10232 29495 10284 29504
rect 10232 29461 10241 29495
rect 10241 29461 10275 29495
rect 10275 29461 10284 29495
rect 10232 29452 10284 29461
rect 13820 29520 13872 29572
rect 14004 29520 14056 29572
rect 20260 29588 20312 29640
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 23572 29520 23624 29572
rect 25780 29520 25832 29572
rect 14740 29452 14792 29504
rect 21180 29452 21232 29504
rect 23480 29452 23532 29504
rect 24768 29452 24820 29504
rect 24952 29452 25004 29504
rect 26148 29631 26200 29640
rect 26148 29597 26157 29631
rect 26157 29597 26191 29631
rect 26191 29597 26200 29631
rect 26148 29588 26200 29597
rect 26240 29588 26292 29640
rect 27896 29656 27948 29708
rect 29092 29724 29144 29776
rect 30380 29724 30432 29776
rect 31668 29724 31720 29776
rect 27712 29520 27764 29572
rect 30104 29656 30156 29708
rect 32036 29588 32088 29640
rect 32772 29656 32824 29708
rect 33048 29699 33100 29708
rect 33048 29665 33057 29699
rect 33057 29665 33091 29699
rect 33091 29665 33100 29699
rect 33048 29656 33100 29665
rect 27528 29452 27580 29504
rect 30656 29452 30708 29504
rect 6550 29350 6602 29402
rect 6614 29350 6666 29402
rect 6678 29350 6730 29402
rect 6742 29350 6794 29402
rect 6806 29350 6858 29402
rect 14439 29350 14491 29402
rect 14503 29350 14555 29402
rect 14567 29350 14619 29402
rect 14631 29350 14683 29402
rect 14695 29350 14747 29402
rect 22328 29350 22380 29402
rect 22392 29350 22444 29402
rect 22456 29350 22508 29402
rect 22520 29350 22572 29402
rect 22584 29350 22636 29402
rect 30217 29350 30269 29402
rect 30281 29350 30333 29402
rect 30345 29350 30397 29402
rect 30409 29350 30461 29402
rect 30473 29350 30525 29402
rect 4528 29248 4580 29300
rect 5448 29180 5500 29232
rect 5540 29155 5592 29164
rect 5540 29121 5549 29155
rect 5549 29121 5583 29155
rect 5583 29121 5592 29155
rect 5540 29112 5592 29121
rect 5724 29248 5776 29300
rect 6920 29248 6972 29300
rect 4988 29044 5040 29096
rect 5172 29044 5224 29096
rect 11980 29291 12032 29300
rect 11980 29257 11989 29291
rect 11989 29257 12023 29291
rect 12023 29257 12032 29291
rect 11980 29248 12032 29257
rect 13084 29248 13136 29300
rect 14096 29291 14148 29300
rect 14096 29257 14105 29291
rect 14105 29257 14139 29291
rect 14139 29257 14148 29291
rect 14096 29248 14148 29257
rect 7564 29112 7616 29164
rect 10140 29112 10192 29164
rect 12900 29180 12952 29232
rect 6368 28976 6420 29028
rect 5540 28908 5592 28960
rect 8300 28976 8352 29028
rect 10600 29019 10652 29028
rect 10600 28985 10609 29019
rect 10609 28985 10643 29019
rect 10643 28985 10652 29019
rect 10600 28976 10652 28985
rect 13728 29112 13780 29164
rect 14096 29112 14148 29164
rect 14648 29112 14700 29164
rect 14832 29155 14884 29164
rect 14832 29121 14841 29155
rect 14841 29121 14875 29155
rect 14875 29121 14884 29155
rect 14832 29112 14884 29121
rect 15016 29248 15068 29300
rect 15660 29248 15712 29300
rect 17592 29291 17644 29300
rect 17592 29257 17601 29291
rect 17601 29257 17635 29291
rect 17635 29257 17644 29291
rect 17592 29248 17644 29257
rect 19708 29248 19760 29300
rect 22560 29248 22612 29300
rect 23388 29248 23440 29300
rect 25044 29248 25096 29300
rect 26148 29248 26200 29300
rect 29368 29248 29420 29300
rect 32220 29248 32272 29300
rect 15844 29155 15896 29164
rect 15844 29121 15853 29155
rect 15853 29121 15887 29155
rect 15887 29121 15896 29155
rect 15844 29112 15896 29121
rect 16212 29112 16264 29164
rect 16488 29112 16540 29164
rect 12072 29087 12124 29096
rect 12072 29053 12081 29087
rect 12081 29053 12115 29087
rect 12115 29053 12124 29087
rect 12072 29044 12124 29053
rect 14004 29044 14056 29096
rect 17684 29087 17736 29096
rect 17684 29053 17693 29087
rect 17693 29053 17727 29087
rect 17727 29053 17736 29087
rect 17684 29044 17736 29053
rect 19708 29087 19760 29096
rect 19708 29053 19717 29087
rect 19717 29053 19751 29087
rect 19751 29053 19760 29087
rect 19708 29044 19760 29053
rect 8484 28908 8536 28960
rect 10416 28908 10468 28960
rect 10692 28908 10744 28960
rect 10876 28951 10928 28960
rect 10876 28917 10885 28951
rect 10885 28917 10919 28951
rect 10919 28917 10928 28951
rect 10876 28908 10928 28917
rect 10968 28951 11020 28960
rect 10968 28917 10977 28951
rect 10977 28917 11011 28951
rect 11011 28917 11020 28951
rect 10968 28908 11020 28917
rect 11152 28951 11204 28960
rect 11152 28917 11161 28951
rect 11161 28917 11195 28951
rect 11195 28917 11204 28951
rect 11152 28908 11204 28917
rect 11336 28908 11388 28960
rect 12992 28908 13044 28960
rect 13728 28976 13780 29028
rect 14372 28976 14424 29028
rect 14924 28976 14976 29028
rect 17132 28976 17184 29028
rect 17960 29019 18012 29028
rect 17960 28985 17969 29019
rect 17969 28985 18003 29019
rect 18003 28985 18012 29019
rect 17960 28976 18012 28985
rect 23480 29044 23532 29096
rect 23756 29044 23808 29096
rect 27528 29112 27580 29164
rect 27988 29155 28040 29164
rect 27988 29121 27997 29155
rect 27997 29121 28031 29155
rect 28031 29121 28040 29155
rect 27988 29112 28040 29121
rect 28448 29112 28500 29164
rect 21272 28976 21324 29028
rect 21548 29019 21600 29028
rect 21548 28985 21557 29019
rect 21557 28985 21591 29019
rect 21591 28985 21600 29019
rect 21548 28976 21600 28985
rect 22836 28976 22888 29028
rect 23388 28976 23440 29028
rect 27252 29087 27304 29096
rect 27252 29053 27261 29087
rect 27261 29053 27295 29087
rect 27295 29053 27304 29087
rect 27252 29044 27304 29053
rect 31208 29044 31260 29096
rect 31852 29087 31904 29096
rect 31852 29053 31861 29087
rect 31861 29053 31895 29087
rect 31895 29053 31904 29087
rect 31852 29044 31904 29053
rect 26792 28976 26844 29028
rect 20904 28908 20956 28960
rect 24676 28951 24728 28960
rect 24676 28917 24685 28951
rect 24685 28917 24719 28951
rect 24719 28917 24728 28951
rect 24676 28908 24728 28917
rect 26148 28908 26200 28960
rect 27436 28908 27488 28960
rect 29000 28976 29052 29028
rect 30104 28976 30156 29028
rect 28264 28908 28316 28960
rect 29368 28908 29420 28960
rect 31300 28951 31352 28960
rect 31300 28917 31309 28951
rect 31309 28917 31343 28951
rect 31343 28917 31352 28951
rect 31300 28908 31352 28917
rect 31392 28908 31444 28960
rect 32036 28908 32088 28960
rect 32588 29087 32640 29096
rect 32588 29053 32597 29087
rect 32597 29053 32631 29087
rect 32631 29053 32640 29087
rect 32588 29044 32640 29053
rect 33784 29019 33836 29028
rect 33784 28985 33793 29019
rect 33793 28985 33827 29019
rect 33827 28985 33836 29019
rect 33784 28976 33836 28985
rect 33140 28908 33192 28960
rect 7210 28806 7262 28858
rect 7274 28806 7326 28858
rect 7338 28806 7390 28858
rect 7402 28806 7454 28858
rect 7466 28806 7518 28858
rect 15099 28806 15151 28858
rect 15163 28806 15215 28858
rect 15227 28806 15279 28858
rect 15291 28806 15343 28858
rect 15355 28806 15407 28858
rect 22988 28806 23040 28858
rect 23052 28806 23104 28858
rect 23116 28806 23168 28858
rect 23180 28806 23232 28858
rect 23244 28806 23296 28858
rect 30877 28806 30929 28858
rect 30941 28806 30993 28858
rect 31005 28806 31057 28858
rect 31069 28806 31121 28858
rect 31133 28806 31185 28858
rect 5540 28704 5592 28756
rect 7932 28704 7984 28756
rect 8300 28747 8352 28756
rect 8300 28713 8309 28747
rect 8309 28713 8343 28747
rect 8343 28713 8352 28747
rect 8300 28704 8352 28713
rect 8484 28747 8536 28756
rect 8484 28713 8493 28747
rect 8493 28713 8527 28747
rect 8527 28713 8536 28747
rect 8484 28704 8536 28713
rect 10232 28704 10284 28756
rect 1308 28568 1360 28620
rect 4436 28611 4488 28620
rect 4436 28577 4445 28611
rect 4445 28577 4479 28611
rect 4479 28577 4488 28611
rect 4436 28568 4488 28577
rect 7564 28636 7616 28688
rect 10048 28636 10100 28688
rect 10784 28704 10836 28756
rect 10968 28704 11020 28756
rect 13636 28704 13688 28756
rect 14280 28704 14332 28756
rect 14832 28704 14884 28756
rect 8208 28611 8260 28620
rect 8208 28577 8217 28611
rect 8217 28577 8251 28611
rect 8251 28577 8260 28611
rect 8208 28568 8260 28577
rect 5356 28543 5408 28552
rect 5356 28509 5365 28543
rect 5365 28509 5399 28543
rect 5399 28509 5408 28543
rect 5356 28500 5408 28509
rect 7012 28500 7064 28552
rect 9864 28543 9916 28552
rect 9864 28509 9873 28543
rect 9873 28509 9907 28543
rect 9907 28509 9916 28543
rect 9864 28500 9916 28509
rect 10324 28679 10376 28688
rect 10324 28645 10333 28679
rect 10333 28645 10367 28679
rect 10367 28645 10376 28679
rect 10324 28636 10376 28645
rect 10416 28679 10468 28688
rect 10416 28645 10451 28679
rect 10451 28645 10468 28679
rect 10416 28636 10468 28645
rect 10692 28611 10744 28620
rect 10692 28577 10701 28611
rect 10701 28577 10735 28611
rect 10735 28577 10744 28611
rect 10692 28568 10744 28577
rect 10508 28500 10560 28552
rect 10968 28611 11020 28620
rect 10968 28577 10977 28611
rect 10977 28577 11011 28611
rect 11011 28577 11020 28611
rect 10968 28568 11020 28577
rect 11336 28568 11388 28620
rect 10600 28432 10652 28484
rect 13636 28568 13688 28620
rect 14740 28611 14792 28620
rect 14740 28577 14749 28611
rect 14749 28577 14783 28611
rect 14783 28577 14792 28611
rect 14740 28568 14792 28577
rect 14924 28611 14976 28620
rect 14924 28577 14933 28611
rect 14933 28577 14967 28611
rect 14967 28577 14976 28611
rect 14924 28568 14976 28577
rect 15016 28568 15068 28620
rect 16580 28704 16632 28756
rect 17132 28747 17184 28756
rect 17132 28713 17141 28747
rect 17141 28713 17175 28747
rect 17175 28713 17184 28747
rect 17132 28704 17184 28713
rect 17960 28704 18012 28756
rect 12440 28543 12492 28552
rect 12440 28509 12449 28543
rect 12449 28509 12483 28543
rect 12483 28509 12492 28543
rect 12440 28500 12492 28509
rect 15476 28500 15528 28552
rect 9220 28407 9272 28416
rect 9220 28373 9229 28407
rect 9229 28373 9263 28407
rect 9263 28373 9272 28407
rect 9220 28364 9272 28373
rect 10876 28364 10928 28416
rect 11612 28364 11664 28416
rect 12624 28407 12676 28416
rect 12624 28373 12633 28407
rect 12633 28373 12667 28407
rect 12667 28373 12676 28407
rect 12624 28364 12676 28373
rect 13820 28432 13872 28484
rect 14372 28432 14424 28484
rect 13176 28407 13228 28416
rect 13176 28373 13185 28407
rect 13185 28373 13219 28407
rect 13219 28373 13228 28407
rect 13176 28364 13228 28373
rect 13360 28364 13412 28416
rect 13912 28364 13964 28416
rect 15844 28568 15896 28620
rect 16396 28611 16448 28620
rect 16396 28577 16405 28611
rect 16405 28577 16439 28611
rect 16439 28577 16448 28611
rect 16396 28568 16448 28577
rect 19156 28636 19208 28688
rect 21548 28747 21600 28756
rect 21548 28713 21557 28747
rect 21557 28713 21591 28747
rect 21591 28713 21600 28747
rect 21548 28704 21600 28713
rect 19708 28636 19760 28688
rect 21916 28636 21968 28688
rect 22560 28679 22612 28688
rect 22560 28645 22569 28679
rect 22569 28645 22603 28679
rect 22603 28645 22612 28679
rect 22560 28636 22612 28645
rect 19248 28611 19300 28620
rect 19248 28577 19257 28611
rect 19257 28577 19291 28611
rect 19291 28577 19300 28611
rect 19248 28568 19300 28577
rect 19616 28611 19668 28620
rect 19616 28577 19625 28611
rect 19625 28577 19659 28611
rect 19659 28577 19668 28611
rect 19616 28568 19668 28577
rect 21088 28568 21140 28620
rect 22652 28611 22704 28620
rect 22652 28577 22661 28611
rect 22661 28577 22695 28611
rect 22695 28577 22704 28611
rect 22652 28568 22704 28577
rect 22836 28704 22888 28756
rect 23388 28704 23440 28756
rect 27252 28704 27304 28756
rect 27804 28704 27856 28756
rect 28264 28704 28316 28756
rect 29000 28704 29052 28756
rect 31208 28704 31260 28756
rect 22836 28611 22888 28620
rect 22836 28577 22845 28611
rect 22845 28577 22879 28611
rect 22879 28577 22888 28611
rect 22836 28568 22888 28577
rect 23480 28679 23532 28688
rect 23480 28645 23489 28679
rect 23489 28645 23523 28679
rect 23523 28645 23532 28679
rect 23480 28636 23532 28645
rect 24676 28636 24728 28688
rect 26884 28636 26936 28688
rect 27436 28568 27488 28620
rect 27528 28568 27580 28620
rect 27804 28611 27856 28620
rect 27804 28577 27813 28611
rect 27813 28577 27847 28611
rect 27847 28577 27856 28611
rect 27804 28568 27856 28577
rect 27896 28568 27948 28620
rect 31300 28679 31352 28688
rect 31300 28645 31309 28679
rect 31309 28645 31343 28679
rect 31343 28645 31352 28679
rect 31300 28636 31352 28645
rect 32036 28636 32088 28688
rect 28632 28568 28684 28620
rect 30564 28568 30616 28620
rect 33140 28568 33192 28620
rect 24768 28500 24820 28552
rect 25228 28543 25280 28552
rect 25228 28509 25237 28543
rect 25237 28509 25271 28543
rect 25271 28509 25280 28543
rect 25228 28500 25280 28509
rect 17500 28364 17552 28416
rect 24032 28364 24084 28416
rect 25872 28543 25924 28552
rect 25872 28509 25881 28543
rect 25881 28509 25915 28543
rect 25915 28509 25924 28543
rect 25872 28500 25924 28509
rect 29184 28543 29236 28552
rect 29184 28509 29193 28543
rect 29193 28509 29227 28543
rect 29227 28509 29236 28543
rect 29184 28500 29236 28509
rect 29460 28543 29512 28552
rect 29460 28509 29469 28543
rect 29469 28509 29503 28543
rect 29503 28509 29512 28543
rect 29460 28500 29512 28509
rect 28448 28432 28500 28484
rect 27804 28364 27856 28416
rect 30656 28500 30708 28552
rect 31024 28543 31076 28552
rect 31024 28509 31033 28543
rect 31033 28509 31067 28543
rect 31067 28509 31076 28543
rect 31024 28500 31076 28509
rect 33416 28543 33468 28552
rect 33416 28509 33425 28543
rect 33425 28509 33459 28543
rect 33459 28509 33468 28543
rect 33416 28500 33468 28509
rect 32312 28364 32364 28416
rect 32588 28364 32640 28416
rect 32864 28407 32916 28416
rect 32864 28373 32873 28407
rect 32873 28373 32907 28407
rect 32907 28373 32916 28407
rect 32864 28364 32916 28373
rect 33876 28407 33928 28416
rect 33876 28373 33885 28407
rect 33885 28373 33919 28407
rect 33919 28373 33928 28407
rect 33876 28364 33928 28373
rect 6550 28262 6602 28314
rect 6614 28262 6666 28314
rect 6678 28262 6730 28314
rect 6742 28262 6794 28314
rect 6806 28262 6858 28314
rect 14439 28262 14491 28314
rect 14503 28262 14555 28314
rect 14567 28262 14619 28314
rect 14631 28262 14683 28314
rect 14695 28262 14747 28314
rect 22328 28262 22380 28314
rect 22392 28262 22444 28314
rect 22456 28262 22508 28314
rect 22520 28262 22572 28314
rect 22584 28262 22636 28314
rect 30217 28262 30269 28314
rect 30281 28262 30333 28314
rect 30345 28262 30397 28314
rect 30409 28262 30461 28314
rect 30473 28262 30525 28314
rect 5356 28160 5408 28212
rect 9220 28160 9272 28212
rect 9864 28160 9916 28212
rect 12440 28160 12492 28212
rect 12992 28203 13044 28212
rect 12992 28169 13001 28203
rect 13001 28169 13035 28203
rect 13035 28169 13044 28203
rect 12992 28160 13044 28169
rect 13176 28160 13228 28212
rect 14096 28203 14148 28212
rect 14096 28169 14105 28203
rect 14105 28169 14139 28203
rect 14139 28169 14148 28203
rect 14096 28160 14148 28169
rect 3976 27999 4028 28008
rect 3976 27965 3985 27999
rect 3985 27965 4019 27999
rect 4019 27965 4028 27999
rect 3976 27956 4028 27965
rect 7840 28024 7892 28076
rect 11980 28092 12032 28144
rect 12256 28092 12308 28144
rect 11152 28024 11204 28076
rect 13360 28067 13412 28076
rect 13360 28033 13369 28067
rect 13369 28033 13403 28067
rect 13403 28033 13412 28067
rect 13360 28024 13412 28033
rect 13636 28024 13688 28076
rect 15752 28160 15804 28212
rect 16396 28160 16448 28212
rect 17500 28203 17552 28212
rect 17500 28169 17509 28203
rect 17509 28169 17543 28203
rect 17543 28169 17552 28203
rect 17500 28160 17552 28169
rect 20904 28160 20956 28212
rect 23388 28160 23440 28212
rect 24032 28160 24084 28212
rect 22836 28092 22888 28144
rect 25228 28160 25280 28212
rect 25872 28160 25924 28212
rect 26884 28160 26936 28212
rect 28356 28160 28408 28212
rect 28816 28160 28868 28212
rect 29276 28160 29328 28212
rect 29460 28160 29512 28212
rect 31852 28160 31904 28212
rect 14372 28067 14424 28076
rect 14372 28033 14381 28067
rect 14381 28033 14415 28067
rect 14415 28033 14424 28067
rect 14372 28024 14424 28033
rect 25044 28024 25096 28076
rect 28908 28092 28960 28144
rect 6736 27888 6788 27940
rect 4528 27863 4580 27872
rect 4528 27829 4537 27863
rect 4537 27829 4571 27863
rect 4571 27829 4580 27863
rect 4528 27820 4580 27829
rect 8392 27888 8444 27940
rect 10876 27956 10928 28008
rect 10508 27888 10560 27940
rect 11244 27999 11296 28008
rect 11244 27965 11253 27999
rect 11253 27965 11287 27999
rect 11287 27965 11296 27999
rect 11244 27956 11296 27965
rect 11428 27999 11480 28008
rect 11428 27965 11437 27999
rect 11437 27965 11471 27999
rect 11471 27965 11480 27999
rect 11428 27956 11480 27965
rect 13268 27999 13320 28008
rect 13268 27965 13277 27999
rect 13277 27965 13311 27999
rect 13311 27965 13320 27999
rect 13268 27956 13320 27965
rect 13544 27999 13596 28008
rect 13544 27965 13553 27999
rect 13553 27965 13587 27999
rect 13587 27965 13596 27999
rect 13544 27956 13596 27965
rect 11336 27888 11388 27940
rect 12900 27888 12952 27940
rect 14004 27956 14056 28008
rect 14280 27956 14332 28008
rect 17684 27956 17736 28008
rect 20076 27956 20128 28008
rect 20904 27956 20956 28008
rect 24216 27956 24268 28008
rect 15476 27888 15528 27940
rect 16028 27931 16080 27940
rect 16028 27897 16037 27931
rect 16037 27897 16071 27931
rect 16071 27897 16080 27931
rect 16028 27888 16080 27897
rect 16764 27888 16816 27940
rect 7564 27820 7616 27872
rect 8024 27820 8076 27872
rect 11704 27820 11756 27872
rect 13084 27863 13136 27872
rect 13084 27829 13093 27863
rect 13093 27829 13127 27863
rect 13127 27829 13136 27863
rect 13084 27820 13136 27829
rect 13820 27820 13872 27872
rect 14004 27820 14056 27872
rect 14648 27863 14700 27872
rect 14648 27829 14657 27863
rect 14657 27829 14691 27863
rect 14691 27829 14700 27863
rect 14648 27820 14700 27829
rect 15568 27820 15620 27872
rect 17776 27863 17828 27872
rect 17776 27829 17785 27863
rect 17785 27829 17819 27863
rect 17819 27829 17828 27863
rect 17776 27820 17828 27829
rect 18052 27820 18104 27872
rect 20996 27863 21048 27872
rect 20996 27829 21005 27863
rect 21005 27829 21039 27863
rect 21039 27829 21048 27863
rect 20996 27820 21048 27829
rect 21916 27863 21968 27872
rect 21916 27829 21925 27863
rect 21925 27829 21959 27863
rect 21959 27829 21968 27863
rect 21916 27820 21968 27829
rect 22192 27820 22244 27872
rect 22560 27820 22612 27872
rect 22652 27820 22704 27872
rect 25136 27820 25188 27872
rect 26148 27956 26200 28008
rect 26700 27999 26752 28008
rect 26700 27965 26709 27999
rect 26709 27965 26743 27999
rect 26743 27965 26752 27999
rect 26700 27956 26752 27965
rect 28724 27956 28776 28008
rect 30012 27956 30064 28008
rect 30380 27956 30432 28008
rect 31392 28024 31444 28076
rect 31668 28024 31720 28076
rect 32864 28024 32916 28076
rect 31024 27956 31076 28008
rect 33876 27956 33928 28008
rect 27528 27888 27580 27940
rect 27620 27931 27672 27940
rect 27620 27897 27629 27931
rect 27629 27897 27663 27931
rect 27663 27897 27672 27931
rect 27620 27888 27672 27897
rect 32312 27888 32364 27940
rect 32680 27888 32732 27940
rect 29368 27820 29420 27872
rect 30656 27820 30708 27872
rect 7210 27718 7262 27770
rect 7274 27718 7326 27770
rect 7338 27718 7390 27770
rect 7402 27718 7454 27770
rect 7466 27718 7518 27770
rect 15099 27718 15151 27770
rect 15163 27718 15215 27770
rect 15227 27718 15279 27770
rect 15291 27718 15343 27770
rect 15355 27718 15407 27770
rect 22988 27718 23040 27770
rect 23052 27718 23104 27770
rect 23116 27718 23168 27770
rect 23180 27718 23232 27770
rect 23244 27718 23296 27770
rect 30877 27718 30929 27770
rect 30941 27718 30993 27770
rect 31005 27718 31057 27770
rect 31069 27718 31121 27770
rect 31133 27718 31185 27770
rect 6736 27659 6788 27668
rect 6736 27625 6745 27659
rect 6745 27625 6779 27659
rect 6779 27625 6788 27659
rect 6736 27616 6788 27625
rect 8208 27616 8260 27668
rect 8392 27659 8444 27668
rect 8392 27625 8401 27659
rect 8401 27625 8435 27659
rect 8435 27625 8444 27659
rect 8392 27616 8444 27625
rect 11152 27616 11204 27668
rect 11244 27616 11296 27668
rect 11612 27616 11664 27668
rect 12624 27616 12676 27668
rect 4528 27591 4580 27600
rect 4528 27557 4537 27591
rect 4537 27557 4571 27591
rect 4571 27557 4580 27591
rect 4528 27548 4580 27557
rect 7012 27591 7064 27600
rect 7012 27557 7021 27591
rect 7021 27557 7055 27591
rect 7055 27557 7064 27591
rect 7012 27548 7064 27557
rect 5080 27523 5132 27532
rect 5080 27489 5089 27523
rect 5089 27489 5123 27523
rect 5123 27489 5132 27523
rect 5080 27480 5132 27489
rect 5540 27480 5592 27532
rect 5264 27455 5316 27464
rect 5264 27421 5273 27455
rect 5273 27421 5307 27455
rect 5307 27421 5316 27455
rect 5264 27412 5316 27421
rect 5356 27412 5408 27464
rect 7104 27523 7156 27532
rect 7104 27489 7113 27523
rect 7113 27489 7147 27523
rect 7147 27489 7156 27523
rect 7104 27480 7156 27489
rect 7564 27480 7616 27532
rect 10968 27548 11020 27600
rect 9956 27480 10008 27532
rect 10784 27480 10836 27532
rect 11980 27548 12032 27600
rect 13912 27548 13964 27600
rect 14096 27548 14148 27600
rect 14372 27659 14424 27668
rect 14372 27625 14381 27659
rect 14381 27625 14415 27659
rect 14415 27625 14424 27659
rect 14372 27616 14424 27625
rect 11796 27523 11848 27532
rect 4436 27276 4488 27328
rect 5816 27319 5868 27328
rect 5816 27285 5825 27319
rect 5825 27285 5859 27319
rect 5859 27285 5868 27319
rect 5816 27276 5868 27285
rect 6000 27276 6052 27328
rect 10968 27412 11020 27464
rect 11796 27489 11805 27523
rect 11805 27489 11839 27523
rect 11839 27489 11848 27523
rect 11796 27480 11848 27489
rect 12164 27480 12216 27532
rect 14372 27480 14424 27532
rect 15476 27616 15528 27668
rect 15568 27616 15620 27668
rect 16028 27616 16080 27668
rect 16580 27616 16632 27668
rect 16764 27659 16816 27668
rect 16764 27625 16773 27659
rect 16773 27625 16807 27659
rect 16807 27625 16816 27659
rect 16764 27616 16816 27625
rect 17040 27616 17092 27668
rect 17776 27659 17828 27668
rect 17776 27625 17785 27659
rect 17785 27625 17819 27659
rect 17819 27625 17828 27659
rect 17776 27616 17828 27625
rect 18052 27616 18104 27668
rect 17224 27591 17276 27600
rect 17224 27557 17233 27591
rect 17233 27557 17267 27591
rect 17267 27557 17276 27591
rect 17224 27548 17276 27557
rect 20076 27659 20128 27668
rect 20076 27625 20085 27659
rect 20085 27625 20119 27659
rect 20119 27625 20128 27659
rect 20076 27616 20128 27625
rect 28172 27659 28224 27668
rect 19064 27548 19116 27600
rect 20996 27548 21048 27600
rect 21824 27548 21876 27600
rect 14648 27412 14700 27464
rect 15844 27412 15896 27464
rect 17224 27412 17276 27464
rect 7748 27276 7800 27328
rect 9588 27319 9640 27328
rect 9588 27285 9597 27319
rect 9597 27285 9631 27319
rect 9631 27285 9640 27319
rect 9588 27276 9640 27285
rect 11060 27276 11112 27328
rect 11520 27276 11572 27328
rect 13820 27276 13872 27328
rect 14924 27344 14976 27396
rect 14280 27276 14332 27328
rect 15476 27276 15528 27328
rect 19248 27412 19300 27464
rect 21088 27412 21140 27464
rect 21732 27455 21784 27464
rect 21732 27421 21741 27455
rect 21741 27421 21775 27455
rect 21775 27421 21784 27455
rect 21732 27412 21784 27421
rect 23388 27548 23440 27600
rect 23756 27591 23808 27600
rect 23756 27557 23765 27591
rect 23765 27557 23799 27591
rect 23799 27557 23808 27591
rect 23756 27548 23808 27557
rect 24676 27548 24728 27600
rect 26148 27548 26200 27600
rect 28172 27625 28181 27659
rect 28181 27625 28215 27659
rect 28215 27625 28224 27659
rect 28172 27616 28224 27625
rect 28724 27659 28776 27668
rect 28724 27625 28733 27659
rect 28733 27625 28767 27659
rect 28767 27625 28776 27659
rect 28724 27616 28776 27625
rect 24216 27480 24268 27532
rect 28356 27548 28408 27600
rect 27712 27523 27764 27532
rect 27712 27489 27721 27523
rect 27721 27489 27755 27523
rect 27755 27489 27764 27523
rect 27712 27480 27764 27489
rect 18972 27276 19024 27328
rect 20260 27319 20312 27328
rect 20260 27285 20269 27319
rect 20269 27285 20303 27319
rect 20303 27285 20312 27319
rect 20260 27276 20312 27285
rect 24308 27455 24360 27464
rect 24308 27421 24317 27455
rect 24317 27421 24351 27455
rect 24351 27421 24360 27455
rect 24308 27412 24360 27421
rect 24860 27412 24912 27464
rect 26332 27455 26384 27464
rect 26332 27421 26341 27455
rect 26341 27421 26375 27455
rect 26375 27421 26384 27455
rect 26332 27412 26384 27421
rect 27160 27412 27212 27464
rect 28632 27480 28684 27532
rect 30104 27548 30156 27600
rect 30564 27616 30616 27668
rect 31668 27616 31720 27668
rect 32036 27616 32088 27668
rect 32496 27659 32548 27668
rect 32496 27625 32505 27659
rect 32505 27625 32539 27659
rect 32539 27625 32548 27659
rect 32496 27616 32548 27625
rect 32680 27616 32732 27668
rect 28908 27523 28960 27532
rect 28908 27489 28917 27523
rect 28917 27489 28951 27523
rect 28951 27489 28960 27523
rect 28908 27480 28960 27489
rect 29276 27523 29328 27532
rect 29276 27489 29285 27523
rect 29285 27489 29319 27523
rect 29319 27489 29328 27523
rect 29276 27480 29328 27489
rect 21272 27276 21324 27328
rect 22008 27276 22060 27328
rect 23296 27276 23348 27328
rect 24124 27276 24176 27328
rect 26700 27319 26752 27328
rect 26700 27285 26709 27319
rect 26709 27285 26743 27319
rect 26743 27285 26752 27319
rect 26700 27276 26752 27285
rect 27068 27319 27120 27328
rect 27068 27285 27077 27319
rect 27077 27285 27111 27319
rect 27111 27285 27120 27319
rect 27068 27276 27120 27285
rect 27620 27344 27672 27396
rect 30380 27480 30432 27532
rect 31392 27548 31444 27600
rect 29552 27455 29604 27464
rect 29552 27421 29561 27455
rect 29561 27421 29595 27455
rect 29595 27421 29604 27455
rect 29552 27412 29604 27421
rect 30104 27455 30156 27464
rect 30104 27421 30113 27455
rect 30113 27421 30147 27455
rect 30147 27421 30156 27455
rect 30104 27412 30156 27421
rect 30564 27455 30616 27464
rect 30564 27421 30573 27455
rect 30573 27421 30607 27455
rect 30607 27421 30616 27455
rect 30564 27412 30616 27421
rect 28172 27276 28224 27328
rect 29276 27276 29328 27328
rect 32036 27455 32088 27464
rect 32036 27421 32045 27455
rect 32045 27421 32079 27455
rect 32079 27421 32088 27455
rect 32036 27412 32088 27421
rect 32128 27412 32180 27464
rect 32404 27412 32456 27464
rect 33048 27412 33100 27464
rect 33416 27412 33468 27464
rect 32588 27344 32640 27396
rect 35164 27344 35216 27396
rect 30748 27276 30800 27328
rect 31392 27276 31444 27328
rect 32036 27276 32088 27328
rect 33784 27319 33836 27328
rect 33784 27285 33793 27319
rect 33793 27285 33827 27319
rect 33827 27285 33836 27319
rect 33784 27276 33836 27285
rect 6550 27174 6602 27226
rect 6614 27174 6666 27226
rect 6678 27174 6730 27226
rect 6742 27174 6794 27226
rect 6806 27174 6858 27226
rect 14439 27174 14491 27226
rect 14503 27174 14555 27226
rect 14567 27174 14619 27226
rect 14631 27174 14683 27226
rect 14695 27174 14747 27226
rect 22328 27174 22380 27226
rect 22392 27174 22444 27226
rect 22456 27174 22508 27226
rect 22520 27174 22572 27226
rect 22584 27174 22636 27226
rect 30217 27174 30269 27226
rect 30281 27174 30333 27226
rect 30345 27174 30397 27226
rect 30409 27174 30461 27226
rect 30473 27174 30525 27226
rect 3976 27115 4028 27124
rect 3976 27081 3985 27115
rect 3985 27081 4019 27115
rect 4019 27081 4028 27115
rect 3976 27072 4028 27081
rect 5264 27072 5316 27124
rect 6092 27072 6144 27124
rect 6368 27072 6420 27124
rect 7840 27115 7892 27124
rect 7840 27081 7849 27115
rect 7849 27081 7883 27115
rect 7883 27081 7892 27115
rect 7840 27072 7892 27081
rect 8208 27072 8260 27124
rect 10048 27072 10100 27124
rect 11428 27072 11480 27124
rect 4436 26979 4488 26988
rect 4436 26945 4445 26979
rect 4445 26945 4479 26979
rect 4479 26945 4488 26979
rect 4436 26936 4488 26945
rect 5632 27004 5684 27056
rect 1308 26868 1360 26920
rect 4620 26936 4672 26988
rect 11336 27004 11388 27056
rect 4896 26868 4948 26920
rect 6184 26868 6236 26920
rect 6276 26911 6328 26920
rect 6276 26877 6285 26911
rect 6285 26877 6319 26911
rect 6319 26877 6328 26911
rect 6276 26868 6328 26877
rect 8024 26868 8076 26920
rect 10600 26868 10652 26920
rect 11060 26936 11112 26988
rect 11520 27004 11572 27056
rect 12624 27072 12676 27124
rect 14096 27072 14148 27124
rect 14832 27072 14884 27124
rect 14280 27004 14332 27056
rect 11796 26936 11848 26988
rect 13084 26936 13136 26988
rect 13820 26936 13872 26988
rect 5540 26800 5592 26852
rect 5724 26800 5776 26852
rect 3608 26732 3660 26784
rect 4896 26732 4948 26784
rect 8852 26843 8904 26852
rect 8852 26809 8861 26843
rect 8861 26809 8895 26843
rect 8895 26809 8904 26843
rect 8852 26800 8904 26809
rect 9588 26800 9640 26852
rect 10416 26800 10468 26852
rect 12440 26868 12492 26920
rect 15844 27115 15896 27124
rect 15844 27081 15853 27115
rect 15853 27081 15887 27115
rect 15887 27081 15896 27115
rect 15844 27072 15896 27081
rect 15936 27072 15988 27124
rect 19064 27072 19116 27124
rect 21732 27072 21784 27124
rect 21824 27072 21876 27124
rect 22008 27072 22060 27124
rect 7196 26732 7248 26784
rect 10600 26775 10652 26784
rect 10600 26741 10609 26775
rect 10609 26741 10643 26775
rect 10643 26741 10652 26775
rect 10600 26732 10652 26741
rect 11888 26775 11940 26784
rect 11888 26741 11897 26775
rect 11897 26741 11931 26775
rect 11931 26741 11940 26775
rect 11888 26732 11940 26741
rect 11980 26775 12032 26784
rect 11980 26741 11989 26775
rect 11989 26741 12023 26775
rect 12023 26741 12032 26775
rect 11980 26732 12032 26741
rect 12716 26775 12768 26784
rect 12716 26741 12725 26775
rect 12725 26741 12759 26775
rect 12759 26741 12768 26775
rect 12716 26732 12768 26741
rect 13636 26843 13688 26852
rect 13636 26809 13645 26843
rect 13645 26809 13679 26843
rect 13679 26809 13688 26843
rect 13636 26800 13688 26809
rect 14648 26843 14700 26852
rect 14648 26809 14657 26843
rect 14657 26809 14691 26843
rect 14691 26809 14700 26843
rect 14648 26800 14700 26809
rect 15476 26911 15528 26920
rect 15476 26877 15485 26911
rect 15485 26877 15519 26911
rect 15519 26877 15528 26911
rect 15476 26868 15528 26877
rect 17684 26936 17736 26988
rect 18052 26936 18104 26988
rect 21916 26936 21968 26988
rect 24124 27072 24176 27124
rect 24860 27072 24912 27124
rect 26332 27072 26384 27124
rect 30564 27072 30616 27124
rect 32588 27072 32640 27124
rect 33048 27072 33100 27124
rect 24032 26936 24084 26988
rect 27068 26936 27120 26988
rect 28080 26936 28132 26988
rect 29184 26936 29236 26988
rect 33140 27004 33192 27056
rect 31852 26936 31904 26988
rect 32220 26936 32272 26988
rect 20904 26868 20956 26920
rect 21088 26911 21140 26920
rect 21088 26877 21097 26911
rect 21097 26877 21131 26911
rect 21131 26877 21140 26911
rect 21088 26868 21140 26877
rect 21180 26911 21232 26920
rect 21180 26877 21189 26911
rect 21189 26877 21223 26911
rect 21223 26877 21232 26911
rect 21180 26868 21232 26877
rect 21364 26868 21416 26920
rect 14832 26800 14884 26852
rect 15660 26800 15712 26852
rect 16304 26800 16356 26852
rect 17224 26800 17276 26852
rect 19064 26800 19116 26852
rect 14188 26732 14240 26784
rect 14740 26732 14792 26784
rect 21640 26800 21692 26852
rect 23296 26800 23348 26852
rect 21916 26732 21968 26784
rect 22192 26732 22244 26784
rect 24492 26868 24544 26920
rect 24676 26911 24728 26920
rect 24676 26877 24685 26911
rect 24685 26877 24719 26911
rect 24719 26877 24728 26911
rect 24676 26868 24728 26877
rect 24768 26911 24820 26920
rect 24768 26877 24777 26911
rect 24777 26877 24811 26911
rect 24811 26877 24820 26911
rect 24768 26868 24820 26877
rect 24584 26843 24636 26852
rect 24584 26809 24593 26843
rect 24593 26809 24627 26843
rect 24627 26809 24636 26843
rect 24584 26800 24636 26809
rect 25688 26911 25740 26920
rect 25688 26877 25697 26911
rect 25697 26877 25731 26911
rect 25731 26877 25740 26911
rect 25688 26868 25740 26877
rect 26240 26800 26292 26852
rect 26332 26843 26384 26852
rect 26332 26809 26341 26843
rect 26341 26809 26375 26843
rect 26375 26809 26384 26843
rect 26332 26800 26384 26809
rect 26884 26800 26936 26852
rect 24860 26732 24912 26784
rect 26976 26732 27028 26784
rect 28632 26911 28684 26920
rect 28632 26877 28641 26911
rect 28641 26877 28675 26911
rect 28675 26877 28684 26911
rect 28632 26868 28684 26877
rect 30656 26868 30708 26920
rect 33416 26868 33468 26920
rect 29552 26843 29604 26852
rect 29552 26809 29561 26843
rect 29561 26809 29595 26843
rect 29595 26809 29604 26843
rect 29552 26800 29604 26809
rect 31484 26843 31536 26852
rect 31484 26809 31493 26843
rect 31493 26809 31527 26843
rect 31527 26809 31536 26843
rect 31484 26800 31536 26809
rect 27988 26732 28040 26784
rect 29276 26732 29328 26784
rect 32496 26732 32548 26784
rect 7210 26630 7262 26682
rect 7274 26630 7326 26682
rect 7338 26630 7390 26682
rect 7402 26630 7454 26682
rect 7466 26630 7518 26682
rect 15099 26630 15151 26682
rect 15163 26630 15215 26682
rect 15227 26630 15279 26682
rect 15291 26630 15343 26682
rect 15355 26630 15407 26682
rect 22988 26630 23040 26682
rect 23052 26630 23104 26682
rect 23116 26630 23168 26682
rect 23180 26630 23232 26682
rect 23244 26630 23296 26682
rect 30877 26630 30929 26682
rect 30941 26630 30993 26682
rect 31005 26630 31057 26682
rect 31069 26630 31121 26682
rect 31133 26630 31185 26682
rect 4620 26528 4672 26580
rect 5724 26528 5776 26580
rect 5816 26528 5868 26580
rect 6184 26528 6236 26580
rect 8852 26528 8904 26580
rect 10692 26571 10744 26580
rect 10692 26537 10701 26571
rect 10701 26537 10735 26571
rect 10735 26537 10744 26571
rect 10692 26528 10744 26537
rect 11428 26528 11480 26580
rect 11888 26528 11940 26580
rect 13636 26528 13688 26580
rect 13728 26528 13780 26580
rect 13912 26528 13964 26580
rect 14096 26528 14148 26580
rect 15752 26528 15804 26580
rect 16304 26528 16356 26580
rect 17592 26528 17644 26580
rect 4252 26435 4304 26444
rect 4252 26401 4261 26435
rect 4261 26401 4295 26435
rect 4295 26401 4304 26435
rect 4252 26392 4304 26401
rect 8024 26392 8076 26444
rect 11704 26392 11756 26444
rect 12440 26392 12492 26444
rect 12624 26392 12676 26444
rect 21640 26460 21692 26512
rect 24584 26528 24636 26580
rect 26884 26571 26936 26580
rect 26884 26537 26893 26571
rect 26893 26537 26927 26571
rect 26927 26537 26936 26571
rect 26884 26528 26936 26537
rect 27160 26571 27212 26580
rect 27160 26537 27169 26571
rect 27169 26537 27203 26571
rect 27203 26537 27212 26571
rect 27160 26528 27212 26537
rect 30104 26528 30156 26580
rect 31484 26571 31536 26580
rect 31484 26537 31493 26571
rect 31493 26537 31527 26571
rect 31527 26537 31536 26571
rect 31484 26528 31536 26537
rect 32036 26528 32088 26580
rect 23848 26460 23900 26512
rect 25872 26460 25924 26512
rect 3240 26367 3292 26376
rect 3240 26333 3249 26367
rect 3249 26333 3283 26367
rect 3283 26333 3292 26367
rect 3240 26324 3292 26333
rect 6920 26367 6972 26376
rect 6920 26333 6929 26367
rect 6929 26333 6963 26367
rect 6963 26333 6972 26367
rect 6920 26324 6972 26333
rect 7656 26367 7708 26376
rect 7656 26333 7665 26367
rect 7665 26333 7699 26367
rect 7699 26333 7708 26367
rect 7656 26324 7708 26333
rect 9864 26367 9916 26376
rect 9864 26333 9873 26367
rect 9873 26333 9907 26367
rect 9907 26333 9916 26367
rect 9864 26324 9916 26333
rect 11888 26299 11940 26308
rect 11888 26265 11897 26299
rect 11897 26265 11931 26299
rect 11931 26265 11940 26299
rect 11888 26256 11940 26265
rect 14188 26392 14240 26444
rect 14740 26435 14792 26444
rect 14740 26401 14749 26435
rect 14749 26401 14783 26435
rect 14783 26401 14792 26435
rect 14740 26392 14792 26401
rect 15568 26435 15620 26444
rect 15568 26401 15577 26435
rect 15577 26401 15611 26435
rect 15611 26401 15620 26435
rect 15568 26392 15620 26401
rect 16580 26435 16632 26444
rect 16580 26401 16589 26435
rect 16589 26401 16623 26435
rect 16623 26401 16632 26435
rect 16580 26392 16632 26401
rect 17868 26392 17920 26444
rect 18972 26435 19024 26444
rect 18972 26401 18981 26435
rect 18981 26401 19015 26435
rect 19015 26401 19024 26435
rect 18972 26392 19024 26401
rect 13912 26256 13964 26308
rect 6368 26231 6420 26240
rect 6368 26197 6377 26231
rect 6377 26197 6411 26231
rect 6411 26197 6420 26231
rect 6368 26188 6420 26197
rect 18144 26367 18196 26376
rect 18144 26333 18153 26367
rect 18153 26333 18187 26367
rect 18187 26333 18196 26367
rect 18144 26324 18196 26333
rect 19248 26367 19300 26376
rect 19248 26333 19257 26367
rect 19257 26333 19291 26367
rect 19291 26333 19300 26367
rect 19248 26324 19300 26333
rect 20904 26324 20956 26376
rect 22192 26435 22244 26444
rect 22192 26401 22201 26435
rect 22201 26401 22235 26435
rect 22235 26401 22244 26435
rect 22192 26392 22244 26401
rect 23388 26392 23440 26444
rect 24860 26435 24912 26444
rect 24860 26401 24869 26435
rect 24869 26401 24903 26435
rect 24903 26401 24912 26435
rect 24860 26392 24912 26401
rect 26792 26435 26844 26444
rect 26792 26401 26801 26435
rect 26801 26401 26835 26435
rect 26835 26401 26844 26435
rect 26792 26392 26844 26401
rect 23480 26367 23532 26376
rect 23480 26333 23489 26367
rect 23489 26333 23523 26367
rect 23523 26333 23532 26367
rect 23480 26324 23532 26333
rect 17408 26299 17460 26308
rect 17408 26265 17417 26299
rect 17417 26265 17451 26299
rect 17451 26265 17460 26299
rect 17408 26256 17460 26265
rect 18052 26256 18104 26308
rect 14832 26188 14884 26240
rect 15844 26231 15896 26240
rect 15844 26197 15853 26231
rect 15853 26197 15887 26231
rect 15887 26197 15896 26231
rect 15844 26188 15896 26197
rect 17132 26188 17184 26240
rect 21548 26231 21600 26240
rect 21548 26197 21557 26231
rect 21557 26197 21591 26231
rect 21591 26197 21600 26231
rect 21548 26188 21600 26197
rect 24952 26324 25004 26376
rect 25964 26324 26016 26376
rect 27160 26392 27212 26444
rect 28080 26435 28132 26444
rect 28080 26401 28089 26435
rect 28089 26401 28123 26435
rect 28123 26401 28132 26435
rect 28080 26392 28132 26401
rect 28172 26392 28224 26444
rect 26792 26256 26844 26308
rect 30564 26324 30616 26376
rect 30932 26367 30984 26376
rect 30932 26333 30941 26367
rect 30941 26333 30975 26367
rect 30975 26333 30984 26367
rect 30932 26324 30984 26333
rect 33048 26367 33100 26376
rect 33048 26333 33057 26367
rect 33057 26333 33091 26367
rect 33091 26333 33100 26367
rect 33048 26324 33100 26333
rect 31852 26256 31904 26308
rect 24308 26188 24360 26240
rect 24860 26188 24912 26240
rect 25412 26188 25464 26240
rect 26056 26231 26108 26240
rect 26056 26197 26065 26231
rect 26065 26197 26099 26231
rect 26099 26197 26108 26231
rect 26056 26188 26108 26197
rect 26240 26188 26292 26240
rect 28172 26188 28224 26240
rect 6550 26086 6602 26138
rect 6614 26086 6666 26138
rect 6678 26086 6730 26138
rect 6742 26086 6794 26138
rect 6806 26086 6858 26138
rect 14439 26086 14491 26138
rect 14503 26086 14555 26138
rect 14567 26086 14619 26138
rect 14631 26086 14683 26138
rect 14695 26086 14747 26138
rect 22328 26086 22380 26138
rect 22392 26086 22444 26138
rect 22456 26086 22508 26138
rect 22520 26086 22572 26138
rect 22584 26086 22636 26138
rect 30217 26086 30269 26138
rect 30281 26086 30333 26138
rect 30345 26086 30397 26138
rect 30409 26086 30461 26138
rect 30473 26086 30525 26138
rect 7656 25984 7708 26036
rect 9864 25984 9916 26036
rect 10692 25984 10744 26036
rect 12624 25984 12676 26036
rect 19248 26027 19300 26036
rect 19248 25993 19257 26027
rect 19257 25993 19291 26027
rect 19291 25993 19300 26027
rect 19248 25984 19300 25993
rect 22836 25984 22888 26036
rect 23296 25984 23348 26036
rect 4988 25848 5040 25900
rect 6368 25848 6420 25900
rect 7656 25848 7708 25900
rect 4804 25780 4856 25832
rect 10324 25848 10376 25900
rect 13544 25916 13596 25968
rect 13452 25848 13504 25900
rect 10600 25780 10652 25832
rect 10692 25823 10744 25832
rect 10692 25789 10701 25823
rect 10701 25789 10735 25823
rect 10735 25789 10744 25823
rect 10692 25780 10744 25789
rect 11060 25780 11112 25832
rect 13636 25780 13688 25832
rect 13728 25780 13780 25832
rect 17408 25916 17460 25968
rect 14832 25848 14884 25900
rect 17684 25848 17736 25900
rect 17868 25848 17920 25900
rect 16396 25780 16448 25832
rect 17132 25780 17184 25832
rect 18052 25780 18104 25832
rect 21548 25891 21600 25900
rect 21548 25857 21557 25891
rect 21557 25857 21591 25891
rect 21591 25857 21600 25891
rect 21548 25848 21600 25857
rect 25872 26027 25924 26036
rect 25872 25993 25881 26027
rect 25881 25993 25915 26027
rect 25915 25993 25924 26027
rect 25872 25984 25924 25993
rect 26332 25984 26384 26036
rect 26424 25984 26476 26036
rect 27896 25984 27948 26036
rect 30932 25984 30984 26036
rect 26516 25916 26568 25968
rect 27344 25959 27396 25968
rect 27344 25925 27353 25959
rect 27353 25925 27387 25959
rect 27387 25925 27396 25959
rect 27344 25916 27396 25925
rect 29000 25916 29052 25968
rect 24032 25848 24084 25900
rect 24860 25848 24912 25900
rect 3884 25687 3936 25696
rect 3884 25653 3893 25687
rect 3893 25653 3927 25687
rect 3927 25653 3936 25687
rect 3884 25644 3936 25653
rect 10416 25644 10468 25696
rect 11980 25755 12032 25764
rect 11980 25721 11989 25755
rect 11989 25721 12023 25755
rect 12023 25721 12032 25755
rect 11980 25712 12032 25721
rect 13268 25712 13320 25764
rect 12072 25644 12124 25696
rect 15476 25712 15528 25764
rect 15844 25712 15896 25764
rect 16672 25712 16724 25764
rect 14188 25687 14240 25696
rect 14188 25653 14197 25687
rect 14197 25653 14231 25687
rect 14231 25653 14240 25687
rect 14188 25644 14240 25653
rect 14464 25644 14516 25696
rect 17776 25644 17828 25696
rect 18512 25644 18564 25696
rect 19156 25780 19208 25832
rect 18880 25755 18932 25764
rect 18880 25721 18889 25755
rect 18889 25721 18923 25755
rect 18923 25721 18932 25755
rect 18880 25712 18932 25721
rect 18972 25755 19024 25764
rect 18972 25721 18981 25755
rect 18981 25721 19015 25755
rect 19015 25721 19024 25755
rect 18972 25712 19024 25721
rect 21180 25780 21232 25832
rect 21272 25823 21324 25832
rect 21272 25789 21281 25823
rect 21281 25789 21315 25823
rect 21315 25789 21324 25823
rect 21272 25780 21324 25789
rect 26148 25780 26200 25832
rect 26516 25780 26568 25832
rect 21456 25712 21508 25764
rect 22560 25712 22612 25764
rect 19524 25687 19576 25696
rect 19524 25653 19533 25687
rect 19533 25653 19567 25687
rect 19567 25653 19576 25687
rect 19524 25644 19576 25653
rect 19616 25644 19668 25696
rect 20628 25644 20680 25696
rect 20996 25687 21048 25696
rect 20996 25653 21005 25687
rect 21005 25653 21039 25687
rect 21039 25653 21048 25687
rect 20996 25644 21048 25653
rect 22376 25644 22428 25696
rect 25412 25712 25464 25764
rect 26240 25644 26292 25696
rect 26608 25644 26660 25696
rect 26884 25644 26936 25696
rect 27160 25780 27212 25832
rect 29184 25848 29236 25900
rect 29368 25848 29420 25900
rect 28172 25712 28224 25764
rect 29276 25712 29328 25764
rect 30748 25712 30800 25764
rect 30564 25644 30616 25696
rect 32496 25644 32548 25696
rect 33048 25644 33100 25696
rect 7210 25542 7262 25594
rect 7274 25542 7326 25594
rect 7338 25542 7390 25594
rect 7402 25542 7454 25594
rect 7466 25542 7518 25594
rect 15099 25542 15151 25594
rect 15163 25542 15215 25594
rect 15227 25542 15279 25594
rect 15291 25542 15343 25594
rect 15355 25542 15407 25594
rect 22988 25542 23040 25594
rect 23052 25542 23104 25594
rect 23116 25542 23168 25594
rect 23180 25542 23232 25594
rect 23244 25542 23296 25594
rect 30877 25542 30929 25594
rect 30941 25542 30993 25594
rect 31005 25542 31057 25594
rect 31069 25542 31121 25594
rect 31133 25542 31185 25594
rect 6920 25440 6972 25492
rect 9680 25440 9732 25492
rect 10692 25440 10744 25492
rect 11336 25440 11388 25492
rect 12164 25440 12216 25492
rect 13268 25440 13320 25492
rect 13452 25440 13504 25492
rect 3884 25372 3936 25424
rect 4252 25372 4304 25424
rect 6184 25372 6236 25424
rect 8208 25372 8260 25424
rect 8760 25372 8812 25424
rect 11428 25372 11480 25424
rect 4804 25347 4856 25356
rect 4804 25313 4813 25347
rect 4813 25313 4847 25347
rect 4847 25313 4856 25347
rect 4804 25304 4856 25313
rect 6552 25304 6604 25356
rect 5632 25236 5684 25288
rect 6460 25168 6512 25220
rect 5908 25143 5960 25152
rect 5908 25109 5917 25143
rect 5917 25109 5951 25143
rect 5951 25109 5960 25143
rect 8024 25347 8076 25356
rect 8024 25313 8033 25347
rect 8033 25313 8067 25347
rect 8067 25313 8076 25347
rect 8024 25304 8076 25313
rect 12256 25372 12308 25424
rect 8852 25236 8904 25288
rect 12072 25347 12124 25356
rect 12072 25313 12081 25347
rect 12081 25313 12115 25347
rect 12115 25313 12124 25347
rect 12072 25304 12124 25313
rect 13728 25347 13780 25356
rect 13728 25313 13737 25347
rect 13737 25313 13771 25347
rect 13771 25313 13780 25347
rect 13728 25304 13780 25313
rect 14924 25440 14976 25492
rect 17684 25440 17736 25492
rect 19616 25440 19668 25492
rect 14188 25372 14240 25424
rect 16396 25372 16448 25424
rect 17408 25372 17460 25424
rect 14464 25236 14516 25288
rect 16672 25236 16724 25288
rect 17776 25236 17828 25288
rect 18604 25236 18656 25288
rect 18696 25236 18748 25288
rect 19156 25304 19208 25356
rect 19524 25304 19576 25356
rect 19984 25440 20036 25492
rect 21272 25440 21324 25492
rect 21456 25483 21508 25492
rect 21456 25449 21465 25483
rect 21465 25449 21499 25483
rect 21499 25449 21508 25483
rect 21456 25440 21508 25449
rect 20996 25372 21048 25424
rect 22376 25440 22428 25492
rect 22560 25440 22612 25492
rect 22192 25372 22244 25424
rect 23112 25440 23164 25492
rect 23388 25372 23440 25424
rect 20536 25236 20588 25288
rect 20628 25236 20680 25288
rect 22100 25279 22152 25288
rect 22100 25245 22109 25279
rect 22109 25245 22143 25279
rect 22143 25245 22152 25279
rect 22100 25236 22152 25245
rect 5908 25100 5960 25109
rect 6920 25100 6972 25152
rect 7748 25100 7800 25152
rect 10416 25100 10468 25152
rect 11612 25143 11664 25152
rect 11612 25109 11621 25143
rect 11621 25109 11655 25143
rect 11655 25109 11664 25143
rect 11612 25100 11664 25109
rect 12256 25168 12308 25220
rect 12440 25168 12492 25220
rect 13636 25168 13688 25220
rect 15568 25211 15620 25220
rect 15568 25177 15577 25211
rect 15577 25177 15611 25211
rect 15611 25177 15620 25211
rect 15568 25168 15620 25177
rect 15844 25168 15896 25220
rect 16580 25168 16632 25220
rect 18512 25168 18564 25220
rect 19616 25143 19668 25152
rect 19616 25109 19625 25143
rect 19625 25109 19659 25143
rect 19659 25109 19668 25143
rect 19616 25100 19668 25109
rect 22928 25347 22980 25356
rect 22928 25313 22937 25347
rect 22937 25313 22971 25347
rect 22971 25313 22980 25347
rect 22928 25304 22980 25313
rect 24768 25440 24820 25492
rect 25688 25440 25740 25492
rect 26976 25440 27028 25492
rect 27344 25440 27396 25492
rect 28908 25440 28960 25492
rect 24860 25304 24912 25356
rect 23480 25279 23532 25288
rect 23480 25245 23489 25279
rect 23489 25245 23523 25279
rect 23523 25245 23532 25279
rect 23480 25236 23532 25245
rect 23756 25279 23808 25288
rect 23756 25245 23765 25279
rect 23765 25245 23799 25279
rect 23799 25245 23808 25279
rect 23756 25236 23808 25245
rect 25320 25279 25372 25288
rect 25320 25245 25329 25279
rect 25329 25245 25363 25279
rect 25363 25245 25372 25279
rect 25320 25236 25372 25245
rect 27528 25304 27580 25356
rect 26700 25236 26752 25288
rect 27068 25279 27120 25288
rect 27068 25245 27077 25279
rect 27077 25245 27111 25279
rect 27111 25245 27120 25279
rect 27068 25236 27120 25245
rect 23296 25143 23348 25152
rect 23296 25109 23305 25143
rect 23305 25109 23339 25143
rect 23339 25109 23348 25143
rect 23296 25100 23348 25109
rect 28632 25304 28684 25356
rect 30104 25304 30156 25356
rect 27804 25279 27856 25288
rect 27804 25245 27813 25279
rect 27813 25245 27847 25279
rect 27847 25245 27856 25279
rect 27804 25236 27856 25245
rect 27896 25236 27948 25288
rect 29828 25279 29880 25288
rect 29828 25245 29837 25279
rect 29837 25245 29871 25279
rect 29871 25245 29880 25279
rect 29828 25236 29880 25245
rect 27712 25100 27764 25152
rect 28448 25143 28500 25152
rect 28448 25109 28457 25143
rect 28457 25109 28491 25143
rect 28491 25109 28500 25143
rect 28448 25100 28500 25109
rect 29368 25100 29420 25152
rect 30564 25100 30616 25152
rect 6550 24998 6602 25050
rect 6614 24998 6666 25050
rect 6678 24998 6730 25050
rect 6742 24998 6794 25050
rect 6806 24998 6858 25050
rect 14439 24998 14491 25050
rect 14503 24998 14555 25050
rect 14567 24998 14619 25050
rect 14631 24998 14683 25050
rect 14695 24998 14747 25050
rect 22328 24998 22380 25050
rect 22392 24998 22444 25050
rect 22456 24998 22508 25050
rect 22520 24998 22572 25050
rect 22584 24998 22636 25050
rect 30217 24998 30269 25050
rect 30281 24998 30333 25050
rect 30345 24998 30397 25050
rect 30409 24998 30461 25050
rect 30473 24998 30525 25050
rect 5632 24896 5684 24948
rect 8760 24896 8812 24948
rect 8852 24896 8904 24948
rect 11428 24896 11480 24948
rect 13728 24896 13780 24948
rect 15844 24896 15896 24948
rect 18236 24896 18288 24948
rect 18604 24939 18656 24948
rect 18604 24905 18613 24939
rect 18613 24905 18647 24939
rect 18647 24905 18656 24939
rect 18604 24896 18656 24905
rect 20536 24939 20588 24948
rect 20536 24905 20545 24939
rect 20545 24905 20579 24939
rect 20579 24905 20588 24939
rect 20536 24896 20588 24905
rect 6368 24828 6420 24880
rect 6552 24828 6604 24880
rect 4252 24803 4304 24812
rect 4252 24769 4261 24803
rect 4261 24769 4295 24803
rect 4295 24769 4304 24803
rect 4252 24760 4304 24769
rect 4896 24760 4948 24812
rect 5540 24760 5592 24812
rect 7840 24760 7892 24812
rect 9128 24760 9180 24812
rect 1308 24692 1360 24744
rect 4344 24735 4396 24744
rect 4344 24701 4353 24735
rect 4353 24701 4387 24735
rect 4387 24701 4396 24735
rect 4344 24692 4396 24701
rect 6736 24692 6788 24744
rect 7656 24692 7708 24744
rect 10600 24760 10652 24812
rect 21732 24828 21784 24880
rect 23480 24896 23532 24948
rect 23756 24896 23808 24948
rect 25412 24939 25464 24948
rect 25412 24905 25421 24939
rect 25421 24905 25455 24939
rect 25455 24905 25464 24939
rect 25412 24896 25464 24905
rect 27068 24896 27120 24948
rect 27804 24939 27856 24948
rect 27804 24905 27813 24939
rect 27813 24905 27847 24939
rect 27847 24905 27856 24939
rect 27804 24896 27856 24905
rect 10232 24735 10284 24744
rect 10232 24701 10241 24735
rect 10241 24701 10275 24735
rect 10275 24701 10284 24735
rect 10232 24692 10284 24701
rect 10508 24692 10560 24744
rect 4896 24556 4948 24608
rect 5448 24556 5500 24608
rect 5632 24556 5684 24608
rect 6184 24556 6236 24608
rect 6368 24599 6420 24608
rect 6368 24565 6377 24599
rect 6377 24565 6411 24599
rect 6411 24565 6420 24599
rect 6368 24556 6420 24565
rect 6920 24599 6972 24608
rect 6920 24565 6929 24599
rect 6929 24565 6963 24599
rect 6963 24565 6972 24599
rect 6920 24556 6972 24565
rect 7012 24556 7064 24608
rect 8576 24556 8628 24608
rect 11336 24692 11388 24744
rect 13636 24760 13688 24812
rect 15660 24760 15712 24812
rect 16396 24803 16448 24812
rect 16396 24769 16405 24803
rect 16405 24769 16439 24803
rect 16439 24769 16448 24803
rect 16396 24760 16448 24769
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 16856 24760 16908 24812
rect 18512 24760 18564 24812
rect 19616 24760 19668 24812
rect 20904 24760 20956 24812
rect 11520 24692 11572 24744
rect 11704 24692 11756 24744
rect 15752 24735 15804 24744
rect 15752 24701 15761 24735
rect 15761 24701 15795 24735
rect 15795 24701 15804 24735
rect 15752 24692 15804 24701
rect 11428 24667 11480 24676
rect 11428 24633 11437 24667
rect 11437 24633 11471 24667
rect 11471 24633 11480 24667
rect 11428 24624 11480 24633
rect 16948 24735 17000 24744
rect 16948 24701 16957 24735
rect 16957 24701 16991 24735
rect 16991 24701 17000 24735
rect 16948 24692 17000 24701
rect 18696 24735 18748 24744
rect 18696 24701 18705 24735
rect 18705 24701 18739 24735
rect 18739 24701 18748 24735
rect 18696 24692 18748 24701
rect 18880 24735 18932 24744
rect 18880 24701 18889 24735
rect 18889 24701 18923 24735
rect 18923 24701 18932 24735
rect 18880 24692 18932 24701
rect 19432 24692 19484 24744
rect 19708 24692 19760 24744
rect 21456 24760 21508 24812
rect 22100 24760 22152 24812
rect 22836 24803 22888 24812
rect 22836 24769 22845 24803
rect 22845 24769 22879 24803
rect 22879 24769 22888 24803
rect 22836 24760 22888 24769
rect 23296 24760 23348 24812
rect 21180 24692 21232 24744
rect 23112 24692 23164 24744
rect 18604 24624 18656 24676
rect 12716 24556 12768 24608
rect 15568 24599 15620 24608
rect 15568 24565 15577 24599
rect 15577 24565 15611 24599
rect 15611 24565 15620 24599
rect 15568 24556 15620 24565
rect 17592 24599 17644 24608
rect 17592 24565 17601 24599
rect 17601 24565 17635 24599
rect 17635 24565 17644 24599
rect 17592 24556 17644 24565
rect 18328 24556 18380 24608
rect 18420 24599 18472 24608
rect 18420 24565 18429 24599
rect 18429 24565 18463 24599
rect 18463 24565 18472 24599
rect 18420 24556 18472 24565
rect 19616 24556 19668 24608
rect 22928 24624 22980 24676
rect 24860 24692 24912 24744
rect 28632 24760 28684 24812
rect 29000 24803 29052 24812
rect 29000 24769 29009 24803
rect 29009 24769 29043 24803
rect 29043 24769 29052 24803
rect 29000 24760 29052 24769
rect 29368 24760 29420 24812
rect 25596 24624 25648 24676
rect 28816 24735 28868 24744
rect 28816 24701 28825 24735
rect 28825 24701 28859 24735
rect 28859 24701 28868 24735
rect 28816 24692 28868 24701
rect 30564 24692 30616 24744
rect 22560 24599 22612 24608
rect 22560 24565 22569 24599
rect 22569 24565 22603 24599
rect 22603 24565 22612 24599
rect 22560 24556 22612 24565
rect 23756 24556 23808 24608
rect 27712 24624 27764 24676
rect 28540 24624 28592 24676
rect 27160 24556 27212 24608
rect 27988 24556 28040 24608
rect 28264 24599 28316 24608
rect 28264 24565 28273 24599
rect 28273 24565 28307 24599
rect 28307 24565 28316 24599
rect 28264 24556 28316 24565
rect 30564 24556 30616 24608
rect 7210 24454 7262 24506
rect 7274 24454 7326 24506
rect 7338 24454 7390 24506
rect 7402 24454 7454 24506
rect 7466 24454 7518 24506
rect 15099 24454 15151 24506
rect 15163 24454 15215 24506
rect 15227 24454 15279 24506
rect 15291 24454 15343 24506
rect 15355 24454 15407 24506
rect 22988 24454 23040 24506
rect 23052 24454 23104 24506
rect 23116 24454 23168 24506
rect 23180 24454 23232 24506
rect 23244 24454 23296 24506
rect 30877 24454 30929 24506
rect 30941 24454 30993 24506
rect 31005 24454 31057 24506
rect 31069 24454 31121 24506
rect 31133 24454 31185 24506
rect 6276 24352 6328 24404
rect 6460 24352 6512 24404
rect 6736 24352 6788 24404
rect 11060 24352 11112 24404
rect 5080 24284 5132 24336
rect 5816 24216 5868 24268
rect 6184 24259 6236 24268
rect 6184 24225 6193 24259
rect 6193 24225 6227 24259
rect 6227 24225 6236 24259
rect 6184 24216 6236 24225
rect 6092 24080 6144 24132
rect 6920 24148 6972 24200
rect 7472 24080 7524 24132
rect 4804 24012 4856 24064
rect 6276 24012 6328 24064
rect 7012 24012 7064 24064
rect 9680 24284 9732 24336
rect 11428 24284 11480 24336
rect 11888 24327 11940 24336
rect 11888 24293 11897 24327
rect 11897 24293 11931 24327
rect 11931 24293 11940 24327
rect 11888 24284 11940 24293
rect 10324 24259 10376 24268
rect 10324 24225 10333 24259
rect 10333 24225 10367 24259
rect 10367 24225 10376 24259
rect 10324 24216 10376 24225
rect 10508 24216 10560 24268
rect 11520 24259 11572 24268
rect 13452 24284 13504 24336
rect 14004 24284 14056 24336
rect 11520 24225 11558 24259
rect 11558 24225 11572 24259
rect 11520 24216 11572 24225
rect 8024 24191 8076 24200
rect 8024 24157 8033 24191
rect 8033 24157 8067 24191
rect 8067 24157 8076 24191
rect 8024 24148 8076 24157
rect 8300 24191 8352 24200
rect 8300 24157 8309 24191
rect 8309 24157 8343 24191
rect 8343 24157 8352 24191
rect 8300 24148 8352 24157
rect 12348 24148 12400 24200
rect 7656 24080 7708 24132
rect 8484 24012 8536 24064
rect 10876 24012 10928 24064
rect 11612 24055 11664 24064
rect 11612 24021 11621 24055
rect 11621 24021 11655 24055
rect 11655 24021 11664 24055
rect 11612 24012 11664 24021
rect 11704 24055 11756 24064
rect 11704 24021 11732 24055
rect 11732 24021 11756 24055
rect 11704 24012 11756 24021
rect 12164 24012 12216 24064
rect 14464 24216 14516 24268
rect 18604 24352 18656 24404
rect 22008 24352 22060 24404
rect 22100 24352 22152 24404
rect 17316 24284 17368 24336
rect 22560 24284 22612 24336
rect 23388 24284 23440 24336
rect 13452 24191 13504 24200
rect 13452 24157 13461 24191
rect 13461 24157 13495 24191
rect 13495 24157 13504 24191
rect 13452 24148 13504 24157
rect 19524 24216 19576 24268
rect 26240 24284 26292 24336
rect 27896 24284 27948 24336
rect 28264 24352 28316 24404
rect 29828 24352 29880 24404
rect 28724 24284 28776 24336
rect 15660 24148 15712 24200
rect 16948 24148 17000 24200
rect 17592 24123 17644 24132
rect 17592 24089 17601 24123
rect 17601 24089 17635 24123
rect 17635 24089 17644 24123
rect 17592 24080 17644 24089
rect 18236 24148 18288 24200
rect 22652 24148 22704 24200
rect 28540 24216 28592 24268
rect 29552 24259 29604 24268
rect 29552 24225 29561 24259
rect 29561 24225 29595 24259
rect 29595 24225 29604 24259
rect 29552 24216 29604 24225
rect 29644 24259 29696 24268
rect 29644 24225 29653 24259
rect 29653 24225 29687 24259
rect 29687 24225 29696 24259
rect 29644 24216 29696 24225
rect 23756 24148 23808 24200
rect 27712 24148 27764 24200
rect 29184 24148 29236 24200
rect 18420 24080 18472 24132
rect 27160 24080 27212 24132
rect 29828 24216 29880 24268
rect 30564 24216 30616 24268
rect 18052 24012 18104 24064
rect 18328 24012 18380 24064
rect 18972 24012 19024 24064
rect 19892 24012 19944 24064
rect 21732 24012 21784 24064
rect 22192 24012 22244 24064
rect 23572 24055 23624 24064
rect 23572 24021 23581 24055
rect 23581 24021 23615 24055
rect 23615 24021 23624 24055
rect 23572 24012 23624 24021
rect 26608 24055 26660 24064
rect 26608 24021 26617 24055
rect 26617 24021 26651 24055
rect 26651 24021 26660 24055
rect 26608 24012 26660 24021
rect 27620 24012 27672 24064
rect 34704 24148 34756 24200
rect 28724 24012 28776 24064
rect 29920 24012 29972 24064
rect 6550 23910 6602 23962
rect 6614 23910 6666 23962
rect 6678 23910 6730 23962
rect 6742 23910 6794 23962
rect 6806 23910 6858 23962
rect 14439 23910 14491 23962
rect 14503 23910 14555 23962
rect 14567 23910 14619 23962
rect 14631 23910 14683 23962
rect 14695 23910 14747 23962
rect 22328 23910 22380 23962
rect 22392 23910 22444 23962
rect 22456 23910 22508 23962
rect 22520 23910 22572 23962
rect 22584 23910 22636 23962
rect 30217 23910 30269 23962
rect 30281 23910 30333 23962
rect 30345 23910 30397 23962
rect 30409 23910 30461 23962
rect 30473 23910 30525 23962
rect 5080 23808 5132 23860
rect 6000 23808 6052 23860
rect 6276 23808 6328 23860
rect 6460 23808 6512 23860
rect 6828 23808 6880 23860
rect 8300 23808 8352 23860
rect 9956 23851 10008 23860
rect 9956 23817 9965 23851
rect 9965 23817 9999 23851
rect 9999 23817 10008 23851
rect 9956 23808 10008 23817
rect 10324 23851 10376 23860
rect 10324 23817 10333 23851
rect 10333 23817 10367 23851
rect 10367 23817 10376 23851
rect 10324 23808 10376 23817
rect 11060 23808 11112 23860
rect 11612 23851 11664 23860
rect 11612 23817 11621 23851
rect 11621 23817 11655 23851
rect 11655 23817 11664 23851
rect 11612 23808 11664 23817
rect 13452 23808 13504 23860
rect 13728 23808 13780 23860
rect 14004 23851 14056 23860
rect 14004 23817 14013 23851
rect 14013 23817 14047 23851
rect 14047 23817 14056 23851
rect 14004 23808 14056 23817
rect 15752 23808 15804 23860
rect 3516 23715 3568 23724
rect 3516 23681 3525 23715
rect 3525 23681 3559 23715
rect 3559 23681 3568 23715
rect 3516 23672 3568 23681
rect 4988 23672 5040 23724
rect 3056 23647 3108 23656
rect 3056 23613 3065 23647
rect 3065 23613 3099 23647
rect 3099 23613 3108 23647
rect 3056 23604 3108 23613
rect 5908 23672 5960 23724
rect 6368 23672 6420 23724
rect 10232 23740 10284 23792
rect 11152 23740 11204 23792
rect 7656 23604 7708 23656
rect 7840 23604 7892 23656
rect 8576 23672 8628 23724
rect 10508 23672 10560 23724
rect 8300 23647 8352 23656
rect 8300 23613 8309 23647
rect 8309 23613 8343 23647
rect 8343 23613 8352 23647
rect 8300 23604 8352 23613
rect 9220 23604 9272 23656
rect 9864 23604 9916 23656
rect 10048 23647 10100 23656
rect 10048 23613 10057 23647
rect 10057 23613 10091 23647
rect 10091 23613 10100 23647
rect 10048 23604 10100 23613
rect 10416 23604 10468 23656
rect 12440 23672 12492 23724
rect 11704 23647 11756 23656
rect 11704 23613 11713 23647
rect 11713 23613 11747 23647
rect 11747 23613 11756 23647
rect 11704 23604 11756 23613
rect 11796 23604 11848 23656
rect 11980 23647 12032 23656
rect 11980 23613 11989 23647
rect 11989 23613 12023 23647
rect 12023 23613 12032 23647
rect 11980 23604 12032 23613
rect 12072 23647 12124 23656
rect 12072 23613 12082 23647
rect 12082 23613 12116 23647
rect 12116 23613 12124 23647
rect 12072 23604 12124 23613
rect 16396 23740 16448 23792
rect 18604 23740 18656 23792
rect 19340 23740 19392 23792
rect 18420 23672 18472 23724
rect 14832 23647 14884 23656
rect 14832 23613 14841 23647
rect 14841 23613 14875 23647
rect 14875 23613 14884 23647
rect 14832 23604 14884 23613
rect 16856 23604 16908 23656
rect 19616 23647 19668 23656
rect 5816 23468 5868 23520
rect 7012 23511 7064 23520
rect 7012 23477 7021 23511
rect 7021 23477 7055 23511
rect 7055 23477 7064 23511
rect 7012 23468 7064 23477
rect 7472 23511 7524 23520
rect 7472 23477 7481 23511
rect 7481 23477 7515 23511
rect 7515 23477 7524 23511
rect 7472 23468 7524 23477
rect 7656 23468 7708 23520
rect 8944 23468 8996 23520
rect 9220 23511 9272 23520
rect 9220 23477 9229 23511
rect 9229 23477 9263 23511
rect 9263 23477 9272 23511
rect 9220 23468 9272 23477
rect 10140 23536 10192 23588
rect 12900 23579 12952 23588
rect 12900 23545 12909 23579
rect 12909 23545 12943 23579
rect 12943 23545 12952 23579
rect 12900 23536 12952 23545
rect 10600 23468 10652 23520
rect 11796 23468 11848 23520
rect 12348 23468 12400 23520
rect 13820 23468 13872 23520
rect 14096 23468 14148 23520
rect 14188 23511 14240 23520
rect 14188 23477 14197 23511
rect 14197 23477 14231 23511
rect 14231 23477 14240 23511
rect 14188 23468 14240 23477
rect 14280 23468 14332 23520
rect 15660 23468 15712 23520
rect 15752 23511 15804 23520
rect 15752 23477 15761 23511
rect 15761 23477 15795 23511
rect 15795 23477 15804 23511
rect 15752 23468 15804 23477
rect 17316 23511 17368 23520
rect 17316 23477 17325 23511
rect 17325 23477 17359 23511
rect 17359 23477 17368 23511
rect 17316 23468 17368 23477
rect 17868 23579 17920 23588
rect 17868 23545 17877 23579
rect 17877 23545 17911 23579
rect 17911 23545 17920 23579
rect 17868 23536 17920 23545
rect 18052 23468 18104 23520
rect 19064 23468 19116 23520
rect 19340 23468 19392 23520
rect 19616 23613 19625 23647
rect 19625 23613 19659 23647
rect 19659 23613 19668 23647
rect 19616 23604 19668 23613
rect 19892 23647 19944 23656
rect 19892 23613 19901 23647
rect 19901 23613 19935 23647
rect 19935 23613 19944 23647
rect 19892 23604 19944 23613
rect 23572 23740 23624 23792
rect 23664 23783 23716 23792
rect 23664 23749 23673 23783
rect 23673 23749 23707 23783
rect 23707 23749 23716 23783
rect 23664 23740 23716 23749
rect 25412 23808 25464 23860
rect 28080 23808 28132 23860
rect 28816 23808 28868 23860
rect 28908 23808 28960 23860
rect 29552 23808 29604 23860
rect 29644 23740 29696 23792
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 20536 23604 20588 23656
rect 19800 23579 19852 23588
rect 19800 23545 19809 23579
rect 19809 23545 19843 23579
rect 19843 23545 19852 23579
rect 19800 23536 19852 23545
rect 21088 23604 21140 23656
rect 21732 23604 21784 23656
rect 24032 23715 24084 23724
rect 24032 23681 24041 23715
rect 24041 23681 24075 23715
rect 24075 23681 24084 23715
rect 24032 23672 24084 23681
rect 25596 23672 25648 23724
rect 26332 23604 26384 23656
rect 26700 23604 26752 23656
rect 27436 23647 27488 23656
rect 27436 23613 27445 23647
rect 27445 23613 27479 23647
rect 27479 23613 27488 23647
rect 27436 23604 27488 23613
rect 20168 23511 20220 23520
rect 20168 23477 20177 23511
rect 20177 23477 20211 23511
rect 20211 23477 20220 23511
rect 20168 23468 20220 23477
rect 20996 23468 21048 23520
rect 25044 23536 25096 23588
rect 27712 23604 27764 23656
rect 27620 23536 27672 23588
rect 27344 23468 27396 23520
rect 28080 23647 28132 23656
rect 28080 23613 28089 23647
rect 28089 23613 28123 23647
rect 28123 23613 28132 23647
rect 28080 23604 28132 23613
rect 28356 23604 28408 23656
rect 33784 23604 33836 23656
rect 29920 23536 29972 23588
rect 28540 23468 28592 23520
rect 28908 23468 28960 23520
rect 7210 23366 7262 23418
rect 7274 23366 7326 23418
rect 7338 23366 7390 23418
rect 7402 23366 7454 23418
rect 7466 23366 7518 23418
rect 15099 23366 15151 23418
rect 15163 23366 15215 23418
rect 15227 23366 15279 23418
rect 15291 23366 15343 23418
rect 15355 23366 15407 23418
rect 22988 23366 23040 23418
rect 23052 23366 23104 23418
rect 23116 23366 23168 23418
rect 23180 23366 23232 23418
rect 23244 23366 23296 23418
rect 30877 23366 30929 23418
rect 30941 23366 30993 23418
rect 31005 23366 31057 23418
rect 31069 23366 31121 23418
rect 31133 23366 31185 23418
rect 8300 23264 8352 23316
rect 5540 23196 5592 23248
rect 7012 23196 7064 23248
rect 7840 23196 7892 23248
rect 5448 23128 5500 23180
rect 9864 23264 9916 23316
rect 9956 23264 10008 23316
rect 8576 23128 8628 23180
rect 9036 23196 9088 23248
rect 9220 23196 9272 23248
rect 9864 23128 9916 23180
rect 10140 23239 10192 23248
rect 10140 23205 10149 23239
rect 10149 23205 10183 23239
rect 10183 23205 10192 23239
rect 10140 23196 10192 23205
rect 10232 23196 10284 23248
rect 10600 23171 10652 23180
rect 10600 23137 10609 23171
rect 10609 23137 10643 23171
rect 10643 23137 10652 23171
rect 10600 23128 10652 23137
rect 3424 23103 3476 23112
rect 3424 23069 3433 23103
rect 3433 23069 3467 23103
rect 3467 23069 3476 23103
rect 3424 23060 3476 23069
rect 7840 23060 7892 23112
rect 9036 23060 9088 23112
rect 9496 23060 9548 23112
rect 9588 23060 9640 23112
rect 11336 23128 11388 23180
rect 14280 23264 14332 23316
rect 15292 23264 15344 23316
rect 19708 23264 19760 23316
rect 20352 23264 20404 23316
rect 22652 23264 22704 23316
rect 25044 23307 25096 23316
rect 25044 23273 25053 23307
rect 25053 23273 25087 23307
rect 25087 23273 25096 23307
rect 25044 23264 25096 23273
rect 26332 23264 26384 23316
rect 26608 23264 26660 23316
rect 27436 23264 27488 23316
rect 11888 23171 11940 23180
rect 11888 23137 11897 23171
rect 11897 23137 11931 23171
rect 11931 23137 11940 23171
rect 11888 23128 11940 23137
rect 14188 23196 14240 23248
rect 16488 23196 16540 23248
rect 12440 23128 12492 23180
rect 12716 23171 12768 23180
rect 12716 23137 12725 23171
rect 12725 23137 12759 23171
rect 12759 23137 12768 23171
rect 12716 23128 12768 23137
rect 14924 23171 14976 23180
rect 14924 23137 14933 23171
rect 14933 23137 14967 23171
rect 14967 23137 14976 23171
rect 14924 23128 14976 23137
rect 16580 23128 16632 23180
rect 3792 22924 3844 22976
rect 4068 22967 4120 22976
rect 4068 22933 4077 22967
rect 4077 22933 4111 22967
rect 4111 22933 4120 22967
rect 4068 22924 4120 22933
rect 4804 22924 4856 22976
rect 5448 22967 5500 22976
rect 5448 22933 5457 22967
rect 5457 22933 5491 22967
rect 5491 22933 5500 22967
rect 5448 22924 5500 22933
rect 9220 22924 9272 22976
rect 9496 22967 9548 22976
rect 9496 22933 9505 22967
rect 9505 22933 9539 22967
rect 9539 22933 9548 22967
rect 9496 22924 9548 22933
rect 9772 23035 9824 23044
rect 9772 23001 9781 23035
rect 9781 23001 9815 23035
rect 9815 23001 9824 23035
rect 9772 22992 9824 23001
rect 10968 22992 11020 23044
rect 11060 23035 11112 23044
rect 11060 23001 11069 23035
rect 11069 23001 11103 23035
rect 11103 23001 11112 23035
rect 11060 22992 11112 23001
rect 12164 23035 12216 23044
rect 12164 23001 12173 23035
rect 12173 23001 12207 23035
rect 12207 23001 12216 23035
rect 12164 22992 12216 23001
rect 11612 22967 11664 22976
rect 11612 22933 11621 22967
rect 11621 22933 11655 22967
rect 11655 22933 11664 22967
rect 11612 22924 11664 22933
rect 13728 23103 13780 23112
rect 13728 23069 13737 23103
rect 13737 23069 13771 23103
rect 13771 23069 13780 23103
rect 13728 23060 13780 23069
rect 13820 23060 13872 23112
rect 14188 23103 14240 23112
rect 14188 23069 14197 23103
rect 14197 23069 14231 23103
rect 14231 23069 14240 23103
rect 14188 23060 14240 23069
rect 15200 23103 15252 23112
rect 15200 23069 15209 23103
rect 15209 23069 15243 23103
rect 15243 23069 15252 23103
rect 15200 23060 15252 23069
rect 15292 23060 15344 23112
rect 15752 23060 15804 23112
rect 17408 23060 17460 23112
rect 18696 23171 18748 23180
rect 18696 23137 18705 23171
rect 18705 23137 18739 23171
rect 18739 23137 18748 23171
rect 18696 23128 18748 23137
rect 20168 23196 20220 23248
rect 20996 23196 21048 23248
rect 19248 23128 19300 23180
rect 19984 23171 20036 23180
rect 19984 23137 19993 23171
rect 19993 23137 20027 23171
rect 20027 23137 20036 23171
rect 19984 23128 20036 23137
rect 21824 23128 21876 23180
rect 23664 23128 23716 23180
rect 19156 23060 19208 23112
rect 12624 22967 12676 22976
rect 12624 22933 12633 22967
rect 12633 22933 12667 22967
rect 12667 22933 12676 22967
rect 12624 22924 12676 22933
rect 13084 22924 13136 22976
rect 16304 22924 16356 22976
rect 16856 22924 16908 22976
rect 17776 22967 17828 22976
rect 17776 22933 17785 22967
rect 17785 22933 17819 22967
rect 17819 22933 17828 22967
rect 17776 22924 17828 22933
rect 18328 22967 18380 22976
rect 18328 22933 18337 22967
rect 18337 22933 18371 22967
rect 18371 22933 18380 22967
rect 18328 22924 18380 22933
rect 19340 22924 19392 22976
rect 23572 23060 23624 23112
rect 25412 23060 25464 23112
rect 25872 23103 25924 23112
rect 25872 23069 25881 23103
rect 25881 23069 25915 23103
rect 25915 23069 25924 23103
rect 25872 23060 25924 23069
rect 25320 22992 25372 23044
rect 25688 22992 25740 23044
rect 24768 22924 24820 22976
rect 28080 23264 28132 23316
rect 30104 23264 30156 23316
rect 27344 23171 27396 23180
rect 27344 23137 27353 23171
rect 27353 23137 27387 23171
rect 27387 23137 27396 23171
rect 27344 23128 27396 23137
rect 27620 23128 27672 23180
rect 27804 23128 27856 23180
rect 28356 23128 28408 23180
rect 28724 23128 28776 23180
rect 29092 23128 29144 23180
rect 26516 23060 26568 23112
rect 28172 23103 28224 23112
rect 28172 23069 28181 23103
rect 28181 23069 28215 23103
rect 28215 23069 28224 23103
rect 28172 23060 28224 23069
rect 29828 23128 29880 23180
rect 27712 22992 27764 23044
rect 27988 22992 28040 23044
rect 31116 23171 31168 23180
rect 31116 23137 31125 23171
rect 31125 23137 31159 23171
rect 31159 23137 31168 23171
rect 31116 23128 31168 23137
rect 31760 23171 31812 23180
rect 30012 23060 30064 23112
rect 31760 23137 31769 23171
rect 31769 23137 31803 23171
rect 31803 23137 31812 23171
rect 31760 23128 31812 23137
rect 29644 22967 29696 22976
rect 29644 22933 29653 22967
rect 29653 22933 29687 22967
rect 29687 22933 29696 22967
rect 29644 22924 29696 22933
rect 29828 22967 29880 22976
rect 29828 22933 29837 22967
rect 29837 22933 29871 22967
rect 29871 22933 29880 22967
rect 29828 22924 29880 22933
rect 30104 22924 30156 22976
rect 30932 22967 30984 22976
rect 30932 22933 30941 22967
rect 30941 22933 30975 22967
rect 30975 22933 30984 22967
rect 30932 22924 30984 22933
rect 6550 22822 6602 22874
rect 6614 22822 6666 22874
rect 6678 22822 6730 22874
rect 6742 22822 6794 22874
rect 6806 22822 6858 22874
rect 14439 22822 14491 22874
rect 14503 22822 14555 22874
rect 14567 22822 14619 22874
rect 14631 22822 14683 22874
rect 14695 22822 14747 22874
rect 22328 22822 22380 22874
rect 22392 22822 22444 22874
rect 22456 22822 22508 22874
rect 22520 22822 22572 22874
rect 22584 22822 22636 22874
rect 30217 22822 30269 22874
rect 30281 22822 30333 22874
rect 30345 22822 30397 22874
rect 30409 22822 30461 22874
rect 30473 22822 30525 22874
rect 3056 22763 3108 22772
rect 3056 22729 3065 22763
rect 3065 22729 3099 22763
rect 3099 22729 3108 22763
rect 3056 22720 3108 22729
rect 5632 22720 5684 22772
rect 9220 22763 9272 22772
rect 9220 22729 9229 22763
rect 9229 22729 9263 22763
rect 9263 22729 9272 22763
rect 9220 22720 9272 22729
rect 9864 22720 9916 22772
rect 10324 22720 10376 22772
rect 13728 22720 13780 22772
rect 14832 22720 14884 22772
rect 15200 22720 15252 22772
rect 16304 22720 16356 22772
rect 16580 22763 16632 22772
rect 16580 22729 16589 22763
rect 16589 22729 16623 22763
rect 16623 22729 16632 22763
rect 16580 22720 16632 22729
rect 17868 22720 17920 22772
rect 18328 22720 18380 22772
rect 19616 22720 19668 22772
rect 19984 22720 20036 22772
rect 24768 22720 24820 22772
rect 25872 22720 25924 22772
rect 8944 22652 8996 22704
rect 4068 22584 4120 22636
rect 4804 22559 4856 22568
rect 4804 22525 4813 22559
rect 4813 22525 4847 22559
rect 4847 22525 4856 22559
rect 4804 22516 4856 22525
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 5448 22559 5500 22568
rect 5448 22525 5457 22559
rect 5457 22525 5491 22559
rect 5491 22525 5500 22559
rect 5448 22516 5500 22525
rect 4712 22380 4764 22432
rect 7748 22448 7800 22500
rect 9496 22516 9548 22568
rect 9772 22559 9824 22568
rect 9772 22525 9781 22559
rect 9781 22525 9815 22559
rect 9815 22525 9824 22559
rect 9772 22516 9824 22525
rect 10968 22695 11020 22704
rect 10968 22661 10977 22695
rect 10977 22661 11011 22695
rect 11011 22661 11020 22695
rect 10968 22652 11020 22661
rect 11888 22652 11940 22704
rect 11980 22627 12032 22636
rect 11980 22593 11989 22627
rect 11989 22593 12023 22627
rect 12023 22593 12032 22627
rect 11980 22584 12032 22593
rect 13084 22584 13136 22636
rect 10876 22516 10928 22568
rect 11244 22516 11296 22568
rect 11428 22516 11480 22568
rect 11612 22516 11664 22568
rect 9588 22448 9640 22500
rect 12624 22516 12676 22568
rect 12716 22559 12768 22568
rect 12716 22525 12725 22559
rect 12725 22525 12759 22559
rect 12759 22525 12768 22559
rect 12716 22516 12768 22525
rect 14096 22516 14148 22568
rect 15016 22516 15068 22568
rect 16672 22559 16724 22568
rect 16672 22525 16681 22559
rect 16681 22525 16715 22559
rect 16715 22525 16724 22559
rect 16672 22516 16724 22525
rect 17224 22559 17276 22568
rect 17224 22525 17233 22559
rect 17233 22525 17267 22559
rect 17267 22525 17276 22559
rect 17224 22516 17276 22525
rect 17868 22516 17920 22568
rect 6000 22380 6052 22432
rect 6460 22380 6512 22432
rect 9036 22380 9088 22432
rect 9956 22380 10008 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 11796 22380 11848 22432
rect 12440 22380 12492 22432
rect 14832 22380 14884 22432
rect 17960 22380 18012 22432
rect 18236 22516 18288 22568
rect 18420 22516 18472 22568
rect 19064 22448 19116 22500
rect 19708 22448 19760 22500
rect 20352 22559 20404 22568
rect 20352 22525 20361 22559
rect 20361 22525 20395 22559
rect 20395 22525 20404 22559
rect 20352 22516 20404 22525
rect 20536 22559 20588 22568
rect 20536 22525 20545 22559
rect 20545 22525 20579 22559
rect 20579 22525 20588 22559
rect 20536 22516 20588 22525
rect 21088 22559 21140 22568
rect 21088 22525 21097 22559
rect 21097 22525 21131 22559
rect 21131 22525 21140 22559
rect 21088 22516 21140 22525
rect 21180 22559 21232 22568
rect 21180 22525 21189 22559
rect 21189 22525 21223 22559
rect 21223 22525 21232 22559
rect 21180 22516 21232 22525
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 26700 22652 26752 22704
rect 22652 22516 22704 22568
rect 23756 22559 23808 22568
rect 23756 22525 23765 22559
rect 23765 22525 23799 22559
rect 23799 22525 23808 22559
rect 23756 22516 23808 22525
rect 21824 22491 21876 22500
rect 21824 22457 21833 22491
rect 21833 22457 21867 22491
rect 21867 22457 21876 22491
rect 21824 22448 21876 22457
rect 20996 22423 21048 22432
rect 20996 22389 21005 22423
rect 21005 22389 21039 22423
rect 21039 22389 21048 22423
rect 20996 22380 21048 22389
rect 21916 22423 21968 22432
rect 21916 22389 21925 22423
rect 21925 22389 21959 22423
rect 21959 22389 21968 22423
rect 21916 22380 21968 22389
rect 22836 22423 22888 22432
rect 22836 22389 22845 22423
rect 22845 22389 22879 22423
rect 22879 22389 22888 22423
rect 22836 22380 22888 22389
rect 23848 22423 23900 22432
rect 23848 22389 23857 22423
rect 23857 22389 23891 22423
rect 23891 22389 23900 22423
rect 23848 22380 23900 22389
rect 25412 22516 25464 22568
rect 26332 22559 26384 22568
rect 26332 22525 26341 22559
rect 26341 22525 26375 22559
rect 26375 22525 26384 22559
rect 26332 22516 26384 22525
rect 28172 22720 28224 22772
rect 31116 22720 31168 22772
rect 31208 22720 31260 22772
rect 31760 22720 31812 22772
rect 27896 22695 27948 22704
rect 27896 22661 27905 22695
rect 27905 22661 27939 22695
rect 27939 22661 27948 22695
rect 27896 22652 27948 22661
rect 28356 22652 28408 22704
rect 26424 22491 26476 22500
rect 26424 22457 26433 22491
rect 26433 22457 26467 22491
rect 26467 22457 26476 22491
rect 26424 22448 26476 22457
rect 26516 22491 26568 22500
rect 26516 22457 26525 22491
rect 26525 22457 26559 22491
rect 26559 22457 26568 22491
rect 26516 22448 26568 22457
rect 29184 22584 29236 22636
rect 31576 22584 31628 22636
rect 27068 22448 27120 22500
rect 28448 22516 28500 22568
rect 33416 22584 33468 22636
rect 35164 22516 35216 22568
rect 29552 22491 29604 22500
rect 29552 22457 29561 22491
rect 29561 22457 29595 22491
rect 29595 22457 29604 22491
rect 29552 22448 29604 22457
rect 30104 22448 30156 22500
rect 25688 22380 25740 22432
rect 27160 22380 27212 22432
rect 28172 22423 28224 22432
rect 28172 22389 28181 22423
rect 28181 22389 28215 22423
rect 28215 22389 28224 22423
rect 28172 22380 28224 22389
rect 28448 22423 28500 22432
rect 28448 22389 28457 22423
rect 28457 22389 28491 22423
rect 28491 22389 28500 22423
rect 28448 22380 28500 22389
rect 32772 22491 32824 22500
rect 32772 22457 32781 22491
rect 32781 22457 32815 22491
rect 32815 22457 32824 22491
rect 32772 22448 32824 22457
rect 33784 22423 33836 22432
rect 33784 22389 33793 22423
rect 33793 22389 33827 22423
rect 33827 22389 33836 22423
rect 33784 22380 33836 22389
rect 7210 22278 7262 22330
rect 7274 22278 7326 22330
rect 7338 22278 7390 22330
rect 7402 22278 7454 22330
rect 7466 22278 7518 22330
rect 15099 22278 15151 22330
rect 15163 22278 15215 22330
rect 15227 22278 15279 22330
rect 15291 22278 15343 22330
rect 15355 22278 15407 22330
rect 22988 22278 23040 22330
rect 23052 22278 23104 22330
rect 23116 22278 23168 22330
rect 23180 22278 23232 22330
rect 23244 22278 23296 22330
rect 30877 22278 30929 22330
rect 30941 22278 30993 22330
rect 31005 22278 31057 22330
rect 31069 22278 31121 22330
rect 31133 22278 31185 22330
rect 3056 22176 3108 22228
rect 3424 22219 3476 22228
rect 3424 22185 3433 22219
rect 3433 22185 3467 22219
rect 3467 22185 3476 22219
rect 3424 22176 3476 22185
rect 3792 22151 3844 22160
rect 3792 22117 3801 22151
rect 3801 22117 3835 22151
rect 3835 22117 3844 22151
rect 3792 22108 3844 22117
rect 4712 22176 4764 22228
rect 5356 22176 5408 22228
rect 7748 22219 7800 22228
rect 7748 22185 7757 22219
rect 7757 22185 7791 22219
rect 7791 22185 7800 22219
rect 7748 22176 7800 22185
rect 7840 22176 7892 22228
rect 8944 22176 8996 22228
rect 9496 22176 9548 22228
rect 9772 22176 9824 22228
rect 4804 22108 4856 22160
rect 8116 22108 8168 22160
rect 3240 21879 3292 21888
rect 3240 21845 3249 21879
rect 3249 21845 3283 21879
rect 3283 21845 3292 21879
rect 3240 21836 3292 21845
rect 4252 21836 4304 21888
rect 4528 22015 4580 22024
rect 4528 21981 4537 22015
rect 4537 21981 4571 22015
rect 4571 21981 4580 22015
rect 4528 21972 4580 21981
rect 5080 21972 5132 22024
rect 5264 21972 5316 22024
rect 8300 22040 8352 22092
rect 10232 22108 10284 22160
rect 11060 22108 11112 22160
rect 9036 22015 9088 22024
rect 9036 21981 9045 22015
rect 9045 21981 9079 22015
rect 9079 21981 9088 22015
rect 9036 21972 9088 21981
rect 9496 21972 9548 22024
rect 10324 22083 10376 22092
rect 10324 22049 10333 22083
rect 10333 22049 10367 22083
rect 10367 22049 10376 22083
rect 10324 22040 10376 22049
rect 12164 22176 12216 22228
rect 17224 22176 17276 22228
rect 17776 22176 17828 22228
rect 14832 22108 14884 22160
rect 18328 22108 18380 22160
rect 21180 22176 21232 22228
rect 20996 22108 21048 22160
rect 21916 22176 21968 22228
rect 11520 22040 11572 22092
rect 12348 22083 12400 22092
rect 12348 22049 12357 22083
rect 12357 22049 12391 22083
rect 12391 22049 12400 22083
rect 12348 22040 12400 22049
rect 13544 22040 13596 22092
rect 15844 22040 15896 22092
rect 10508 21972 10560 22024
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 12256 21972 12308 21981
rect 12624 21972 12676 22024
rect 13820 22015 13872 22024
rect 13820 21981 13829 22015
rect 13829 21981 13863 22015
rect 13863 21981 13872 22015
rect 13820 21972 13872 21981
rect 14004 22015 14056 22024
rect 14004 21981 14013 22015
rect 14013 21981 14047 22015
rect 14047 21981 14056 22015
rect 14004 21972 14056 21981
rect 6000 21904 6052 21956
rect 14832 21972 14884 22024
rect 4896 21836 4948 21888
rect 9588 21879 9640 21888
rect 9588 21845 9597 21879
rect 9597 21845 9631 21879
rect 9631 21845 9640 21879
rect 9588 21836 9640 21845
rect 10324 21879 10376 21888
rect 10324 21845 10333 21879
rect 10333 21845 10367 21879
rect 10367 21845 10376 21879
rect 10324 21836 10376 21845
rect 11152 21836 11204 21888
rect 11520 21836 11572 21888
rect 11704 21836 11756 21888
rect 12072 21836 12124 21888
rect 17500 22040 17552 22092
rect 18880 22083 18932 22092
rect 18880 22049 18889 22083
rect 18889 22049 18923 22083
rect 18923 22049 18932 22083
rect 18880 22040 18932 22049
rect 22652 22176 22704 22228
rect 25136 22176 25188 22228
rect 17408 21972 17460 22024
rect 18972 21972 19024 22024
rect 19064 22015 19116 22024
rect 19064 21981 19073 22015
rect 19073 21981 19107 22015
rect 19107 21981 19116 22015
rect 19064 21972 19116 21981
rect 16672 21879 16724 21888
rect 16672 21845 16681 21879
rect 16681 21845 16715 21879
rect 16715 21845 16724 21879
rect 16672 21836 16724 21845
rect 17592 21947 17644 21956
rect 17592 21913 17601 21947
rect 17601 21913 17635 21947
rect 17635 21913 17644 21947
rect 17592 21904 17644 21913
rect 17868 21836 17920 21888
rect 17960 21879 18012 21888
rect 17960 21845 17969 21879
rect 17969 21845 18003 21879
rect 18003 21845 18012 21879
rect 17960 21836 18012 21845
rect 18696 21904 18748 21956
rect 19616 21972 19668 22024
rect 21732 22015 21784 22024
rect 21732 21981 21741 22015
rect 21741 21981 21775 22015
rect 21775 21981 21784 22015
rect 21732 21972 21784 21981
rect 18236 21836 18288 21888
rect 18420 21836 18472 21888
rect 18788 21879 18840 21888
rect 18788 21845 18797 21879
rect 18797 21845 18831 21879
rect 18831 21845 18840 21879
rect 18788 21836 18840 21845
rect 19708 21836 19760 21888
rect 21916 21836 21968 21888
rect 22008 21879 22060 21888
rect 22008 21845 22017 21879
rect 22017 21845 22051 21879
rect 22051 21845 22060 21879
rect 22008 21836 22060 21845
rect 22192 21836 22244 21888
rect 23296 22108 23348 22160
rect 22928 22083 22980 22092
rect 22928 22049 22937 22083
rect 22937 22049 22971 22083
rect 22971 22049 22980 22083
rect 22928 22040 22980 22049
rect 23848 22108 23900 22160
rect 25412 22176 25464 22228
rect 25964 22176 26016 22228
rect 26332 22176 26384 22228
rect 26424 22176 26476 22228
rect 26700 22176 26752 22228
rect 27436 22176 27488 22228
rect 22744 21972 22796 22024
rect 23204 21972 23256 22024
rect 25688 21972 25740 22024
rect 26700 22040 26752 22092
rect 27068 22083 27120 22092
rect 27068 22049 27077 22083
rect 27077 22049 27111 22083
rect 27111 22049 27120 22083
rect 27620 22108 27672 22160
rect 31576 22176 31628 22228
rect 32772 22176 32824 22228
rect 27068 22040 27120 22049
rect 27896 22040 27948 22092
rect 29276 22108 29328 22160
rect 28080 21972 28132 22024
rect 29092 22040 29144 22092
rect 30656 22108 30708 22160
rect 29552 22083 29604 22092
rect 29552 22049 29561 22083
rect 29561 22049 29595 22083
rect 29595 22049 29604 22083
rect 29552 22040 29604 22049
rect 31944 22108 31996 22160
rect 30104 22015 30156 22024
rect 30104 21981 30113 22015
rect 30113 21981 30147 22015
rect 30147 21981 30156 22015
rect 30104 21972 30156 21981
rect 26976 21904 27028 21956
rect 27068 21904 27120 21956
rect 22560 21836 22612 21888
rect 22744 21836 22796 21888
rect 23296 21836 23348 21888
rect 24124 21836 24176 21888
rect 27620 21879 27672 21888
rect 27620 21845 27629 21879
rect 27629 21845 27663 21879
rect 27663 21845 27672 21879
rect 27620 21836 27672 21845
rect 28172 21836 28224 21888
rect 29000 21836 29052 21888
rect 30564 21836 30616 21888
rect 32404 21879 32456 21888
rect 32404 21845 32413 21879
rect 32413 21845 32447 21879
rect 32447 21845 32456 21879
rect 32404 21836 32456 21845
rect 6550 21734 6602 21786
rect 6614 21734 6666 21786
rect 6678 21734 6730 21786
rect 6742 21734 6794 21786
rect 6806 21734 6858 21786
rect 14439 21734 14491 21786
rect 14503 21734 14555 21786
rect 14567 21734 14619 21786
rect 14631 21734 14683 21786
rect 14695 21734 14747 21786
rect 22328 21734 22380 21786
rect 22392 21734 22444 21786
rect 22456 21734 22508 21786
rect 22520 21734 22572 21786
rect 22584 21734 22636 21786
rect 30217 21734 30269 21786
rect 30281 21734 30333 21786
rect 30345 21734 30397 21786
rect 30409 21734 30461 21786
rect 30473 21734 30525 21786
rect 4528 21632 4580 21684
rect 5816 21632 5868 21684
rect 8024 21632 8076 21684
rect 9680 21632 9732 21684
rect 10508 21632 10560 21684
rect 12348 21632 12400 21684
rect 6920 21564 6972 21616
rect 12256 21564 12308 21616
rect 14372 21632 14424 21684
rect 15016 21632 15068 21684
rect 15844 21675 15896 21684
rect 15844 21641 15853 21675
rect 15853 21641 15887 21675
rect 15887 21641 15896 21675
rect 15844 21632 15896 21641
rect 18144 21675 18196 21684
rect 18144 21641 18153 21675
rect 18153 21641 18187 21675
rect 18187 21641 18196 21675
rect 18144 21632 18196 21641
rect 17868 21564 17920 21616
rect 21364 21632 21416 21684
rect 23388 21632 23440 21684
rect 19524 21564 19576 21616
rect 22560 21564 22612 21616
rect 22928 21564 22980 21616
rect 6000 21496 6052 21548
rect 6092 21539 6144 21548
rect 6092 21505 6101 21539
rect 6101 21505 6135 21539
rect 6135 21505 6144 21539
rect 6092 21496 6144 21505
rect 4804 21471 4856 21480
rect 4804 21437 4813 21471
rect 4813 21437 4847 21471
rect 4847 21437 4856 21471
rect 4804 21428 4856 21437
rect 3240 21360 3292 21412
rect 4528 21403 4580 21412
rect 4528 21369 4537 21403
rect 4537 21369 4571 21403
rect 4571 21369 4580 21403
rect 4528 21360 4580 21369
rect 9864 21496 9916 21548
rect 10600 21496 10652 21548
rect 12072 21496 12124 21548
rect 10140 21428 10192 21480
rect 4344 21292 4396 21344
rect 5632 21292 5684 21344
rect 6092 21360 6144 21412
rect 7656 21360 7708 21412
rect 9128 21403 9180 21412
rect 9128 21369 9137 21403
rect 9137 21369 9171 21403
rect 9171 21369 9180 21403
rect 9128 21360 9180 21369
rect 9772 21403 9824 21412
rect 9772 21369 9781 21403
rect 9781 21369 9815 21403
rect 9815 21369 9824 21403
rect 9772 21360 9824 21369
rect 11336 21360 11388 21412
rect 11612 21471 11664 21480
rect 11612 21437 11621 21471
rect 11621 21437 11655 21471
rect 11655 21437 11664 21471
rect 11612 21428 11664 21437
rect 11704 21428 11756 21480
rect 12624 21496 12676 21548
rect 14004 21496 14056 21548
rect 14188 21496 14240 21548
rect 14648 21539 14700 21548
rect 14648 21505 14657 21539
rect 14657 21505 14691 21539
rect 14691 21505 14700 21539
rect 14648 21496 14700 21505
rect 14924 21496 14976 21548
rect 16672 21539 16724 21548
rect 16672 21505 16681 21539
rect 16681 21505 16715 21539
rect 16715 21505 16724 21539
rect 16672 21496 16724 21505
rect 17132 21496 17184 21548
rect 13912 21428 13964 21480
rect 6184 21292 6236 21344
rect 7012 21292 7064 21344
rect 7840 21292 7892 21344
rect 11060 21292 11112 21344
rect 11612 21292 11664 21344
rect 18788 21428 18840 21480
rect 18972 21428 19024 21480
rect 23480 21496 23532 21548
rect 16764 21360 16816 21412
rect 12256 21292 12308 21344
rect 15016 21292 15068 21344
rect 15660 21292 15712 21344
rect 16672 21292 16724 21344
rect 18788 21292 18840 21344
rect 19064 21292 19116 21344
rect 19524 21292 19576 21344
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 29276 21632 29328 21684
rect 30104 21632 30156 21684
rect 31944 21632 31996 21684
rect 32404 21632 32456 21684
rect 24032 21564 24084 21616
rect 26056 21539 26108 21548
rect 26056 21505 26065 21539
rect 26065 21505 26099 21539
rect 26099 21505 26108 21539
rect 26056 21496 26108 21505
rect 29644 21539 29696 21548
rect 29644 21505 29653 21539
rect 29653 21505 29687 21539
rect 29687 21505 29696 21539
rect 29644 21496 29696 21505
rect 23756 21428 23808 21480
rect 21272 21403 21324 21412
rect 21272 21369 21281 21403
rect 21281 21369 21315 21403
rect 21315 21369 21324 21403
rect 21272 21360 21324 21369
rect 22008 21360 22060 21412
rect 20628 21292 20680 21344
rect 22652 21292 22704 21344
rect 25780 21428 25832 21480
rect 26148 21428 26200 21480
rect 28172 21428 28224 21480
rect 29828 21471 29880 21480
rect 29828 21437 29837 21471
rect 29837 21437 29871 21471
rect 29871 21437 29880 21471
rect 29828 21428 29880 21437
rect 26516 21360 26568 21412
rect 30656 21428 30708 21480
rect 31116 21428 31168 21480
rect 31300 21360 31352 21412
rect 29460 21292 29512 21344
rect 32588 21471 32640 21480
rect 32588 21437 32597 21471
rect 32597 21437 32631 21471
rect 32631 21437 32640 21471
rect 32588 21428 32640 21437
rect 34888 21360 34940 21412
rect 7210 21190 7262 21242
rect 7274 21190 7326 21242
rect 7338 21190 7390 21242
rect 7402 21190 7454 21242
rect 7466 21190 7518 21242
rect 15099 21190 15151 21242
rect 15163 21190 15215 21242
rect 15227 21190 15279 21242
rect 15291 21190 15343 21242
rect 15355 21190 15407 21242
rect 22988 21190 23040 21242
rect 23052 21190 23104 21242
rect 23116 21190 23168 21242
rect 23180 21190 23232 21242
rect 23244 21190 23296 21242
rect 30877 21190 30929 21242
rect 30941 21190 30993 21242
rect 31005 21190 31057 21242
rect 31069 21190 31121 21242
rect 31133 21190 31185 21242
rect 4528 21088 4580 21140
rect 1308 21020 1360 21072
rect 5172 21020 5224 21072
rect 6092 21088 6144 21140
rect 8116 21088 8168 21140
rect 9588 21088 9640 21140
rect 10876 21088 10928 21140
rect 4436 20995 4488 21004
rect 4436 20961 4445 20995
rect 4445 20961 4479 20995
rect 4479 20961 4488 20995
rect 4436 20952 4488 20961
rect 5540 20995 5592 21004
rect 5540 20961 5549 20995
rect 5549 20961 5583 20995
rect 5583 20961 5592 20995
rect 5540 20952 5592 20961
rect 5816 20952 5868 21004
rect 8024 21020 8076 21072
rect 14188 21088 14240 21140
rect 15476 21088 15528 21140
rect 17960 21088 18012 21140
rect 11520 21020 11572 21072
rect 11612 21063 11664 21072
rect 11612 21029 11621 21063
rect 11621 21029 11655 21063
rect 11655 21029 11664 21063
rect 11612 21020 11664 21029
rect 14372 21020 14424 21072
rect 9864 20952 9916 21004
rect 9956 20884 10008 20936
rect 10140 20884 10192 20936
rect 10232 20927 10284 20936
rect 10232 20893 10241 20927
rect 10241 20893 10275 20927
rect 10275 20893 10284 20927
rect 10232 20884 10284 20893
rect 10784 20884 10836 20936
rect 10968 20952 11020 21004
rect 11336 20952 11388 21004
rect 11980 20952 12032 21004
rect 12256 20952 12308 21004
rect 12440 20952 12492 21004
rect 14648 21020 14700 21072
rect 16856 20995 16908 21004
rect 16856 20961 16865 20995
rect 16865 20961 16899 20995
rect 16899 20961 16908 20995
rect 16856 20952 16908 20961
rect 10968 20816 11020 20868
rect 6460 20748 6512 20800
rect 8484 20748 8536 20800
rect 9680 20748 9732 20800
rect 11520 20884 11572 20936
rect 13636 20927 13688 20936
rect 13636 20893 13645 20927
rect 13645 20893 13679 20927
rect 13679 20893 13688 20927
rect 13636 20884 13688 20893
rect 19616 21088 19668 21140
rect 21272 21088 21324 21140
rect 20720 21020 20772 21072
rect 20628 20952 20680 21004
rect 22376 21063 22428 21072
rect 22376 21029 22385 21063
rect 22385 21029 22419 21063
rect 22419 21029 22428 21063
rect 26884 21088 26936 21140
rect 27988 21088 28040 21140
rect 28448 21088 28500 21140
rect 29552 21088 29604 21140
rect 31300 21088 31352 21140
rect 22376 21020 22428 21029
rect 18604 20927 18656 20936
rect 18604 20893 18613 20927
rect 18613 20893 18647 20927
rect 18647 20893 18656 20927
rect 18604 20884 18656 20893
rect 12900 20816 12952 20868
rect 16672 20816 16724 20868
rect 16764 20816 16816 20868
rect 17960 20816 18012 20868
rect 18328 20816 18380 20868
rect 20904 20884 20956 20936
rect 21272 20952 21324 21004
rect 21364 20952 21416 21004
rect 22652 20995 22704 21004
rect 22652 20961 22661 20995
rect 22661 20961 22695 20995
rect 22695 20961 22704 20995
rect 22652 20952 22704 20961
rect 24492 21020 24544 21072
rect 24768 21020 24820 21072
rect 24032 20995 24084 21004
rect 24032 20961 24041 20995
rect 24041 20961 24075 20995
rect 24075 20961 24084 20995
rect 24032 20952 24084 20961
rect 25596 20995 25648 21004
rect 25596 20961 25605 20995
rect 25605 20961 25639 20995
rect 25639 20961 25648 20995
rect 25596 20952 25648 20961
rect 26056 21020 26108 21072
rect 21916 20927 21968 20936
rect 21916 20893 21925 20927
rect 21925 20893 21959 20927
rect 21959 20893 21968 20927
rect 21916 20884 21968 20893
rect 23664 20884 23716 20936
rect 26976 20995 27028 21004
rect 26976 20961 26985 20995
rect 26985 20961 27019 20995
rect 27019 20961 27028 20995
rect 26976 20952 27028 20961
rect 27068 20995 27120 21004
rect 27068 20961 27077 20995
rect 27077 20961 27111 20995
rect 27111 20961 27120 20995
rect 27068 20952 27120 20961
rect 27344 20952 27396 21004
rect 27712 20995 27764 21004
rect 27712 20961 27721 20995
rect 27721 20961 27755 20995
rect 27755 20961 27764 20995
rect 27712 20952 27764 20961
rect 27804 20952 27856 21004
rect 28172 21063 28224 21072
rect 28172 21029 28181 21063
rect 28181 21029 28215 21063
rect 28215 21029 28224 21063
rect 28172 21020 28224 21029
rect 28356 21020 28408 21072
rect 29368 21020 29420 21072
rect 29920 21020 29972 21072
rect 30656 21063 30708 21072
rect 30656 21029 30665 21063
rect 30665 21029 30699 21063
rect 30699 21029 30708 21063
rect 30656 21020 30708 21029
rect 32588 21088 32640 21140
rect 26700 20884 26752 20936
rect 27252 20884 27304 20936
rect 33416 20952 33468 21004
rect 30472 20884 30524 20936
rect 30656 20884 30708 20936
rect 31024 20884 31076 20936
rect 31760 20927 31812 20936
rect 31760 20893 31769 20927
rect 31769 20893 31803 20927
rect 31803 20893 31812 20927
rect 31760 20884 31812 20893
rect 32312 20884 32364 20936
rect 33140 20884 33192 20936
rect 33324 20927 33376 20936
rect 33324 20893 33333 20927
rect 33333 20893 33367 20927
rect 33367 20893 33376 20927
rect 33324 20884 33376 20893
rect 11520 20748 11572 20800
rect 13084 20748 13136 20800
rect 13360 20748 13412 20800
rect 14280 20791 14332 20800
rect 14280 20757 14289 20791
rect 14289 20757 14323 20791
rect 14323 20757 14332 20791
rect 14280 20748 14332 20757
rect 15936 20748 15988 20800
rect 18144 20791 18196 20800
rect 18144 20757 18153 20791
rect 18153 20757 18187 20791
rect 18187 20757 18196 20791
rect 18144 20748 18196 20757
rect 18696 20748 18748 20800
rect 20260 20791 20312 20800
rect 20260 20757 20269 20791
rect 20269 20757 20303 20791
rect 20303 20757 20312 20791
rect 20260 20748 20312 20757
rect 21180 20791 21232 20800
rect 21180 20757 21189 20791
rect 21189 20757 21223 20791
rect 21223 20757 21232 20791
rect 21180 20748 21232 20757
rect 21272 20748 21324 20800
rect 22376 20748 22428 20800
rect 22652 20748 22704 20800
rect 24032 20748 24084 20800
rect 24492 20748 24544 20800
rect 25780 20748 25832 20800
rect 26332 20748 26384 20800
rect 27988 20748 28040 20800
rect 28356 20748 28408 20800
rect 30932 20748 30984 20800
rect 31208 20748 31260 20800
rect 32036 20791 32088 20800
rect 32036 20757 32045 20791
rect 32045 20757 32079 20791
rect 32079 20757 32088 20791
rect 32036 20748 32088 20757
rect 32588 20748 32640 20800
rect 33876 20791 33928 20800
rect 33876 20757 33885 20791
rect 33885 20757 33919 20791
rect 33919 20757 33928 20791
rect 33876 20748 33928 20757
rect 6550 20646 6602 20698
rect 6614 20646 6666 20698
rect 6678 20646 6730 20698
rect 6742 20646 6794 20698
rect 6806 20646 6858 20698
rect 14439 20646 14491 20698
rect 14503 20646 14555 20698
rect 14567 20646 14619 20698
rect 14631 20646 14683 20698
rect 14695 20646 14747 20698
rect 22328 20646 22380 20698
rect 22392 20646 22444 20698
rect 22456 20646 22508 20698
rect 22520 20646 22572 20698
rect 22584 20646 22636 20698
rect 30217 20646 30269 20698
rect 30281 20646 30333 20698
rect 30345 20646 30397 20698
rect 30409 20646 30461 20698
rect 30473 20646 30525 20698
rect 5172 20587 5224 20596
rect 5172 20553 5181 20587
rect 5181 20553 5215 20587
rect 5215 20553 5224 20587
rect 5172 20544 5224 20553
rect 6828 20544 6880 20596
rect 9864 20587 9916 20596
rect 9864 20553 9873 20587
rect 9873 20553 9907 20587
rect 9907 20553 9916 20587
rect 9864 20544 9916 20553
rect 10232 20544 10284 20596
rect 10784 20544 10836 20596
rect 4252 20451 4304 20460
rect 4252 20417 4261 20451
rect 4261 20417 4295 20451
rect 4295 20417 4304 20451
rect 4252 20408 4304 20417
rect 4344 20408 4396 20460
rect 9496 20519 9548 20528
rect 9496 20485 9505 20519
rect 9505 20485 9539 20519
rect 9539 20485 9548 20519
rect 9496 20476 9548 20485
rect 9680 20476 9732 20528
rect 10968 20476 11020 20528
rect 5632 20408 5684 20460
rect 5908 20408 5960 20460
rect 7104 20408 7156 20460
rect 8024 20408 8076 20460
rect 8484 20451 8536 20460
rect 8484 20417 8493 20451
rect 8493 20417 8527 20451
rect 8527 20417 8536 20451
rect 8484 20408 8536 20417
rect 8852 20408 8904 20460
rect 10048 20408 10100 20460
rect 10692 20408 10744 20460
rect 10876 20408 10928 20460
rect 11336 20544 11388 20596
rect 13820 20587 13872 20596
rect 13820 20553 13829 20587
rect 13829 20553 13863 20587
rect 13863 20553 13872 20587
rect 13820 20544 13872 20553
rect 18604 20587 18656 20596
rect 18604 20553 18613 20587
rect 18613 20553 18647 20587
rect 18647 20553 18656 20587
rect 18604 20544 18656 20553
rect 19064 20544 19116 20596
rect 19892 20544 19944 20596
rect 20720 20544 20772 20596
rect 21548 20544 21600 20596
rect 21824 20544 21876 20596
rect 23572 20544 23624 20596
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 12348 20408 12400 20460
rect 14832 20408 14884 20460
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 18052 20408 18104 20460
rect 19156 20451 19208 20460
rect 19156 20417 19165 20451
rect 19165 20417 19199 20451
rect 19199 20417 19208 20451
rect 19156 20408 19208 20417
rect 7840 20383 7892 20392
rect 7840 20349 7849 20383
rect 7849 20349 7883 20383
rect 7883 20349 7892 20383
rect 7840 20340 7892 20349
rect 8116 20340 8168 20392
rect 9956 20340 10008 20392
rect 7656 20272 7708 20324
rect 7932 20272 7984 20324
rect 10048 20272 10100 20324
rect 10416 20272 10468 20324
rect 11428 20383 11480 20392
rect 11428 20349 11437 20383
rect 11437 20349 11471 20383
rect 11471 20349 11480 20383
rect 11428 20340 11480 20349
rect 17960 20340 18012 20392
rect 18880 20340 18932 20392
rect 20260 20408 20312 20460
rect 21456 20408 21508 20460
rect 19432 20383 19484 20392
rect 19432 20349 19441 20383
rect 19441 20349 19475 20383
rect 19475 20349 19484 20383
rect 19432 20340 19484 20349
rect 19708 20340 19760 20392
rect 21088 20383 21140 20392
rect 21088 20349 21097 20383
rect 21097 20349 21131 20383
rect 21131 20349 21140 20383
rect 21088 20340 21140 20349
rect 21272 20340 21324 20392
rect 3700 20247 3752 20256
rect 3700 20213 3709 20247
rect 3709 20213 3743 20247
rect 3743 20213 3752 20247
rect 3700 20204 3752 20213
rect 5356 20204 5408 20256
rect 5724 20247 5776 20256
rect 5724 20213 5733 20247
rect 5733 20213 5767 20247
rect 5767 20213 5776 20247
rect 5724 20204 5776 20213
rect 6368 20204 6420 20256
rect 6828 20204 6880 20256
rect 7012 20204 7064 20256
rect 8024 20247 8076 20256
rect 8024 20213 8033 20247
rect 8033 20213 8067 20247
rect 8067 20213 8076 20247
rect 8024 20204 8076 20213
rect 9404 20204 9456 20256
rect 10600 20204 10652 20256
rect 10876 20204 10928 20256
rect 12992 20272 13044 20324
rect 15200 20272 15252 20324
rect 12072 20204 12124 20256
rect 13452 20247 13504 20256
rect 13452 20213 13461 20247
rect 13461 20213 13495 20247
rect 13495 20213 13504 20247
rect 13452 20204 13504 20213
rect 14280 20204 14332 20256
rect 16028 20315 16080 20324
rect 16028 20281 16037 20315
rect 16037 20281 16071 20315
rect 16071 20281 16080 20315
rect 16028 20272 16080 20281
rect 19984 20272 20036 20324
rect 16764 20204 16816 20256
rect 17868 20204 17920 20256
rect 18880 20204 18932 20256
rect 19892 20204 19944 20256
rect 21824 20340 21876 20392
rect 21916 20383 21968 20392
rect 21916 20349 21925 20383
rect 21925 20349 21959 20383
rect 21959 20349 21968 20383
rect 21916 20340 21968 20349
rect 22560 20408 22612 20460
rect 23940 20408 23992 20460
rect 24124 20451 24176 20460
rect 24124 20417 24133 20451
rect 24133 20417 24167 20451
rect 24167 20417 24176 20451
rect 24124 20408 24176 20417
rect 24492 20408 24544 20460
rect 25596 20544 25648 20596
rect 26240 20544 26292 20596
rect 26424 20587 26476 20596
rect 26424 20553 26433 20587
rect 26433 20553 26467 20587
rect 26467 20553 26476 20587
rect 26424 20544 26476 20553
rect 26700 20544 26752 20596
rect 27160 20544 27212 20596
rect 27620 20587 27672 20596
rect 27620 20553 27629 20587
rect 27629 20553 27663 20587
rect 27663 20553 27672 20587
rect 27620 20544 27672 20553
rect 27712 20544 27764 20596
rect 29460 20587 29512 20596
rect 29460 20553 29469 20587
rect 29469 20553 29503 20587
rect 29503 20553 29512 20587
rect 29460 20544 29512 20553
rect 29828 20544 29880 20596
rect 31760 20544 31812 20596
rect 23848 20204 23900 20256
rect 24124 20204 24176 20256
rect 24676 20204 24728 20256
rect 25780 20272 25832 20324
rect 26332 20408 26384 20460
rect 26056 20340 26108 20392
rect 26608 20340 26660 20392
rect 26148 20272 26200 20324
rect 26332 20272 26384 20324
rect 27528 20340 27580 20392
rect 27620 20383 27672 20392
rect 27620 20349 27629 20383
rect 27629 20349 27663 20383
rect 27663 20349 27672 20383
rect 27620 20340 27672 20349
rect 31484 20476 31536 20528
rect 29368 20408 29420 20460
rect 27436 20315 27488 20324
rect 27436 20281 27445 20315
rect 27445 20281 27479 20315
rect 27479 20281 27488 20315
rect 27436 20272 27488 20281
rect 29644 20383 29696 20392
rect 29644 20349 29653 20383
rect 29653 20349 29687 20383
rect 29687 20349 29696 20383
rect 29644 20340 29696 20349
rect 30656 20340 30708 20392
rect 30932 20408 30984 20460
rect 30840 20340 30892 20392
rect 31024 20383 31076 20392
rect 31024 20349 31033 20383
rect 31033 20349 31067 20383
rect 31067 20349 31076 20383
rect 31024 20340 31076 20349
rect 31392 20340 31444 20392
rect 32588 20408 32640 20460
rect 32036 20340 32088 20392
rect 33876 20340 33928 20392
rect 29920 20315 29972 20324
rect 29920 20281 29961 20315
rect 29961 20281 29972 20315
rect 29920 20272 29972 20281
rect 31576 20315 31628 20324
rect 31576 20281 31585 20315
rect 31585 20281 31619 20315
rect 31619 20281 31628 20315
rect 31576 20272 31628 20281
rect 29828 20204 29880 20256
rect 30104 20247 30156 20256
rect 30104 20213 30113 20247
rect 30113 20213 30147 20247
rect 30147 20213 30156 20247
rect 30104 20204 30156 20213
rect 30564 20204 30616 20256
rect 30748 20204 30800 20256
rect 31024 20204 31076 20256
rect 7210 20102 7262 20154
rect 7274 20102 7326 20154
rect 7338 20102 7390 20154
rect 7402 20102 7454 20154
rect 7466 20102 7518 20154
rect 15099 20102 15151 20154
rect 15163 20102 15215 20154
rect 15227 20102 15279 20154
rect 15291 20102 15343 20154
rect 15355 20102 15407 20154
rect 22988 20102 23040 20154
rect 23052 20102 23104 20154
rect 23116 20102 23168 20154
rect 23180 20102 23232 20154
rect 23244 20102 23296 20154
rect 30877 20102 30929 20154
rect 30941 20102 30993 20154
rect 31005 20102 31057 20154
rect 31069 20102 31121 20154
rect 31133 20102 31185 20154
rect 5356 20000 5408 20052
rect 7656 20000 7708 20052
rect 7932 20000 7984 20052
rect 8024 20000 8076 20052
rect 9036 20000 9088 20052
rect 10416 20000 10468 20052
rect 11428 20000 11480 20052
rect 11520 20000 11572 20052
rect 4620 19932 4672 19984
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 4804 19839 4856 19848
rect 4804 19805 4813 19839
rect 4813 19805 4847 19839
rect 4847 19805 4856 19839
rect 4804 19796 4856 19805
rect 5264 19864 5316 19916
rect 5816 19864 5868 19916
rect 6184 19864 6236 19916
rect 5540 19796 5592 19848
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 9496 19932 9548 19984
rect 12072 19975 12124 19984
rect 12072 19941 12081 19975
rect 12081 19941 12115 19975
rect 12115 19941 12124 19975
rect 12072 19932 12124 19941
rect 5724 19728 5776 19780
rect 7656 19728 7708 19780
rect 9036 19839 9088 19848
rect 9036 19805 9045 19839
rect 9045 19805 9079 19839
rect 9079 19805 9088 19839
rect 9036 19796 9088 19805
rect 10324 19864 10376 19916
rect 10508 19864 10560 19916
rect 10876 19907 10928 19916
rect 10876 19873 10885 19907
rect 10885 19873 10919 19907
rect 10919 19873 10928 19907
rect 10876 19864 10928 19873
rect 10968 19907 11020 19916
rect 10968 19873 10977 19907
rect 10977 19873 11011 19907
rect 11011 19873 11020 19907
rect 10968 19864 11020 19873
rect 10784 19796 10836 19848
rect 11704 19907 11756 19916
rect 11704 19873 11713 19907
rect 11713 19873 11747 19907
rect 11747 19873 11756 19907
rect 11704 19864 11756 19873
rect 12992 20000 13044 20052
rect 13636 20000 13688 20052
rect 15568 20000 15620 20052
rect 16028 20000 16080 20052
rect 16764 20043 16816 20052
rect 16764 20009 16773 20043
rect 16773 20009 16807 20043
rect 16807 20009 16816 20043
rect 16764 20000 16816 20009
rect 17040 20000 17092 20052
rect 18972 20000 19024 20052
rect 19156 20000 19208 20052
rect 20904 20000 20956 20052
rect 21272 20000 21324 20052
rect 13820 19975 13872 19984
rect 13820 19941 13829 19975
rect 13829 19941 13863 19975
rect 13863 19941 13872 19975
rect 13820 19932 13872 19941
rect 14004 19932 14056 19984
rect 14188 19975 14240 19984
rect 14188 19941 14197 19975
rect 14197 19941 14231 19975
rect 14231 19941 14240 19975
rect 14188 19932 14240 19941
rect 16396 19932 16448 19984
rect 12348 19907 12400 19916
rect 12348 19873 12357 19907
rect 12357 19873 12391 19907
rect 12391 19873 12400 19907
rect 12348 19864 12400 19873
rect 13544 19864 13596 19916
rect 4988 19660 5040 19712
rect 5816 19660 5868 19712
rect 8300 19660 8352 19712
rect 8392 19660 8444 19712
rect 10048 19728 10100 19780
rect 10876 19728 10928 19780
rect 12164 19796 12216 19848
rect 13912 19839 13964 19848
rect 13912 19805 13921 19839
rect 13921 19805 13955 19839
rect 13955 19805 13964 19839
rect 13912 19796 13964 19805
rect 10692 19660 10744 19712
rect 11428 19703 11480 19712
rect 11428 19669 11437 19703
rect 11437 19669 11471 19703
rect 11471 19669 11480 19703
rect 11428 19660 11480 19669
rect 13268 19728 13320 19780
rect 16488 19796 16540 19848
rect 17960 19864 18012 19916
rect 17224 19796 17276 19848
rect 19432 19932 19484 19984
rect 19892 19932 19944 19984
rect 20536 19932 20588 19984
rect 22192 20000 22244 20052
rect 26332 20000 26384 20052
rect 27436 20000 27488 20052
rect 18696 19864 18748 19916
rect 19156 19864 19208 19916
rect 22100 19932 22152 19984
rect 24676 19932 24728 19984
rect 18420 19796 18472 19848
rect 18236 19728 18288 19780
rect 19064 19839 19116 19848
rect 19064 19805 19073 19839
rect 19073 19805 19107 19839
rect 19107 19805 19116 19839
rect 19064 19796 19116 19805
rect 19984 19796 20036 19848
rect 20076 19839 20128 19848
rect 20076 19805 20085 19839
rect 20085 19805 20119 19839
rect 20119 19805 20128 19839
rect 20076 19796 20128 19805
rect 20996 19796 21048 19848
rect 12532 19703 12584 19712
rect 12532 19669 12541 19703
rect 12541 19669 12575 19703
rect 12575 19669 12584 19703
rect 12532 19660 12584 19669
rect 17040 19660 17092 19712
rect 17316 19660 17368 19712
rect 17408 19660 17460 19712
rect 17960 19660 18012 19712
rect 18328 19660 18380 19712
rect 19248 19728 19300 19780
rect 19892 19660 19944 19712
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 22560 19728 22612 19780
rect 23664 19864 23716 19916
rect 23848 19864 23900 19916
rect 25320 19975 25372 19984
rect 25320 19941 25329 19975
rect 25329 19941 25363 19975
rect 25363 19941 25372 19975
rect 25320 19932 25372 19941
rect 25688 19864 25740 19916
rect 26240 19864 26292 19916
rect 26792 19864 26844 19916
rect 30748 20000 30800 20052
rect 32312 20043 32364 20052
rect 32312 20009 32321 20043
rect 32321 20009 32355 20043
rect 32355 20009 32364 20043
rect 32312 20000 32364 20009
rect 32404 20000 32456 20052
rect 27344 19864 27396 19916
rect 27896 19864 27948 19916
rect 29368 19932 29420 19984
rect 29644 19932 29696 19984
rect 32772 19932 32824 19984
rect 29736 19864 29788 19916
rect 30564 19907 30616 19916
rect 30564 19873 30573 19907
rect 30573 19873 30607 19907
rect 30607 19873 30616 19907
rect 30564 19864 30616 19873
rect 33140 19864 33192 19916
rect 23480 19796 23532 19848
rect 23572 19728 23624 19780
rect 28080 19796 28132 19848
rect 29000 19796 29052 19848
rect 32312 19796 32364 19848
rect 33048 19796 33100 19848
rect 33324 19796 33376 19848
rect 26056 19728 26108 19780
rect 27068 19728 27120 19780
rect 29644 19728 29696 19780
rect 24952 19703 25004 19712
rect 24952 19669 24973 19703
rect 24973 19669 25004 19703
rect 24952 19660 25004 19669
rect 25780 19660 25832 19712
rect 26608 19660 26660 19712
rect 27528 19660 27580 19712
rect 27988 19703 28040 19712
rect 27988 19669 27997 19703
rect 27997 19669 28031 19703
rect 28031 19669 28040 19703
rect 27988 19660 28040 19669
rect 29000 19660 29052 19712
rect 30656 19660 30708 19712
rect 6550 19558 6602 19610
rect 6614 19558 6666 19610
rect 6678 19558 6730 19610
rect 6742 19558 6794 19610
rect 6806 19558 6858 19610
rect 14439 19558 14491 19610
rect 14503 19558 14555 19610
rect 14567 19558 14619 19610
rect 14631 19558 14683 19610
rect 14695 19558 14747 19610
rect 22328 19558 22380 19610
rect 22392 19558 22444 19610
rect 22456 19558 22508 19610
rect 22520 19558 22572 19610
rect 22584 19558 22636 19610
rect 30217 19558 30269 19610
rect 30281 19558 30333 19610
rect 30345 19558 30397 19610
rect 30409 19558 30461 19610
rect 30473 19558 30525 19610
rect 5172 19456 5224 19508
rect 5540 19456 5592 19508
rect 10968 19456 11020 19508
rect 11336 19499 11388 19508
rect 11336 19465 11345 19499
rect 11345 19465 11379 19499
rect 11379 19465 11388 19499
rect 11336 19456 11388 19465
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 13820 19456 13872 19508
rect 15476 19456 15528 19508
rect 16396 19456 16448 19508
rect 3240 19295 3292 19304
rect 3240 19261 3249 19295
rect 3249 19261 3283 19295
rect 3283 19261 3292 19295
rect 3240 19252 3292 19261
rect 4620 19252 4672 19304
rect 5632 19388 5684 19440
rect 6736 19388 6788 19440
rect 8116 19388 8168 19440
rect 17224 19456 17276 19508
rect 21180 19456 21232 19508
rect 21456 19456 21508 19508
rect 22100 19499 22152 19508
rect 22100 19465 22109 19499
rect 22109 19465 22143 19499
rect 22143 19465 22152 19499
rect 22100 19456 22152 19465
rect 24952 19456 25004 19508
rect 26424 19456 26476 19508
rect 26792 19456 26844 19508
rect 29184 19456 29236 19508
rect 30104 19456 30156 19508
rect 26332 19388 26384 19440
rect 26700 19388 26752 19440
rect 28080 19431 28132 19440
rect 28080 19397 28089 19431
rect 28089 19397 28123 19431
rect 28123 19397 28132 19431
rect 28080 19388 28132 19397
rect 28816 19388 28868 19440
rect 29460 19388 29512 19440
rect 29920 19388 29972 19440
rect 5264 19320 5316 19372
rect 5724 19320 5776 19372
rect 7104 19320 7156 19372
rect 9772 19320 9824 19372
rect 9128 19295 9180 19304
rect 9128 19261 9137 19295
rect 9137 19261 9171 19295
rect 9171 19261 9180 19295
rect 9128 19252 9180 19261
rect 5540 19159 5592 19168
rect 5540 19125 5549 19159
rect 5549 19125 5583 19159
rect 5583 19125 5592 19159
rect 5540 19116 5592 19125
rect 6920 19116 6972 19168
rect 7748 19184 7800 19236
rect 8576 19184 8628 19236
rect 9496 19227 9548 19236
rect 9496 19193 9505 19227
rect 9505 19193 9539 19227
rect 9539 19193 9548 19227
rect 9496 19184 9548 19193
rect 10784 19320 10836 19372
rect 11980 19320 12032 19372
rect 12532 19320 12584 19372
rect 13452 19320 13504 19372
rect 9956 19295 10008 19304
rect 9956 19261 9965 19295
rect 9965 19261 9999 19295
rect 9999 19261 10008 19295
rect 9956 19252 10008 19261
rect 11152 19252 11204 19304
rect 11612 19252 11664 19304
rect 8484 19159 8536 19168
rect 8484 19125 8493 19159
rect 8493 19125 8527 19159
rect 8527 19125 8536 19159
rect 8484 19116 8536 19125
rect 10784 19116 10836 19168
rect 11336 19184 11388 19236
rect 11520 19227 11572 19236
rect 11520 19193 11529 19227
rect 11529 19193 11563 19227
rect 11563 19193 11572 19227
rect 11520 19184 11572 19193
rect 12348 19252 12400 19304
rect 12164 19116 12216 19168
rect 12440 19159 12492 19168
rect 12440 19125 12449 19159
rect 12449 19125 12483 19159
rect 12483 19125 12492 19159
rect 12440 19116 12492 19125
rect 14004 19320 14056 19372
rect 15752 19320 15804 19372
rect 16396 19320 16448 19372
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 19248 19363 19300 19372
rect 19248 19329 19257 19363
rect 19257 19329 19291 19363
rect 19291 19329 19300 19363
rect 19248 19320 19300 19329
rect 23480 19320 23532 19372
rect 23756 19363 23808 19372
rect 23756 19329 23765 19363
rect 23765 19329 23799 19363
rect 23799 19329 23808 19363
rect 23756 19320 23808 19329
rect 14924 19252 14976 19304
rect 16488 19252 16540 19304
rect 17132 19295 17184 19304
rect 17132 19261 17141 19295
rect 17141 19261 17175 19295
rect 17175 19261 17184 19295
rect 17132 19252 17184 19261
rect 21088 19295 21140 19304
rect 21088 19261 21097 19295
rect 21097 19261 21131 19295
rect 21131 19261 21140 19295
rect 21088 19252 21140 19261
rect 14556 19159 14608 19168
rect 14556 19125 14565 19159
rect 14565 19125 14599 19159
rect 14599 19125 14608 19159
rect 14556 19116 14608 19125
rect 15568 19116 15620 19168
rect 23664 19184 23716 19236
rect 20260 19116 20312 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 25320 19295 25372 19304
rect 25320 19261 25329 19295
rect 25329 19261 25363 19295
rect 25363 19261 25372 19295
rect 25320 19252 25372 19261
rect 27160 19295 27212 19304
rect 27160 19261 27169 19295
rect 27169 19261 27203 19295
rect 27203 19261 27212 19295
rect 27160 19252 27212 19261
rect 27344 19320 27396 19372
rect 27896 19320 27948 19372
rect 28264 19295 28316 19304
rect 28264 19261 28273 19295
rect 28273 19261 28307 19295
rect 28307 19261 28316 19295
rect 28264 19252 28316 19261
rect 33784 19363 33836 19372
rect 33784 19329 33793 19363
rect 33793 19329 33827 19363
rect 33827 19329 33836 19363
rect 33784 19320 33836 19329
rect 30656 19252 30708 19304
rect 31300 19252 31352 19304
rect 32772 19295 32824 19304
rect 32772 19261 32781 19295
rect 32781 19261 32815 19295
rect 32815 19261 32824 19295
rect 32772 19252 32824 19261
rect 26056 19159 26108 19168
rect 26056 19125 26065 19159
rect 26065 19125 26099 19159
rect 26099 19125 26108 19159
rect 26056 19116 26108 19125
rect 27252 19227 27304 19236
rect 27252 19193 27287 19227
rect 27287 19193 27304 19227
rect 27252 19184 27304 19193
rect 27436 19116 27488 19168
rect 27712 19159 27764 19168
rect 27712 19125 27721 19159
rect 27721 19125 27755 19159
rect 27755 19125 27764 19159
rect 27712 19116 27764 19125
rect 27804 19159 27856 19168
rect 27804 19125 27813 19159
rect 27813 19125 27847 19159
rect 27847 19125 27856 19159
rect 27804 19116 27856 19125
rect 27896 19159 27948 19168
rect 27896 19125 27905 19159
rect 27905 19125 27939 19159
rect 27939 19125 27948 19159
rect 27896 19116 27948 19125
rect 29828 19184 29880 19236
rect 29092 19159 29144 19168
rect 29092 19125 29101 19159
rect 29101 19125 29135 19159
rect 29135 19125 29144 19159
rect 29092 19116 29144 19125
rect 29276 19159 29328 19168
rect 29276 19125 29285 19159
rect 29285 19125 29319 19159
rect 29319 19125 29328 19159
rect 29276 19116 29328 19125
rect 29368 19159 29420 19168
rect 29368 19125 29377 19159
rect 29377 19125 29411 19159
rect 29411 19125 29420 19159
rect 29368 19116 29420 19125
rect 29552 19116 29604 19168
rect 30012 19116 30064 19168
rect 30288 19116 30340 19168
rect 32496 19159 32548 19168
rect 32496 19125 32505 19159
rect 32505 19125 32539 19159
rect 32539 19125 32548 19159
rect 32496 19116 32548 19125
rect 33048 19116 33100 19168
rect 33692 19116 33744 19168
rect 7210 19014 7262 19066
rect 7274 19014 7326 19066
rect 7338 19014 7390 19066
rect 7402 19014 7454 19066
rect 7466 19014 7518 19066
rect 15099 19014 15151 19066
rect 15163 19014 15215 19066
rect 15227 19014 15279 19066
rect 15291 19014 15343 19066
rect 15355 19014 15407 19066
rect 22988 19014 23040 19066
rect 23052 19014 23104 19066
rect 23116 19014 23168 19066
rect 23180 19014 23232 19066
rect 23244 19014 23296 19066
rect 30877 19014 30929 19066
rect 30941 19014 30993 19066
rect 31005 19014 31057 19066
rect 31069 19014 31121 19066
rect 31133 19014 31185 19066
rect 4528 18912 4580 18964
rect 5264 18912 5316 18964
rect 1308 18776 1360 18828
rect 3700 18776 3752 18828
rect 4804 18844 4856 18896
rect 5540 18844 5592 18896
rect 5816 18844 5868 18896
rect 6368 18844 6420 18896
rect 7012 18912 7064 18964
rect 7656 18912 7708 18964
rect 7748 18955 7800 18964
rect 7748 18921 7757 18955
rect 7757 18921 7791 18955
rect 7791 18921 7800 18955
rect 7748 18912 7800 18921
rect 8484 18912 8536 18964
rect 9128 18912 9180 18964
rect 9496 18912 9548 18964
rect 11888 18912 11940 18964
rect 12164 18912 12216 18964
rect 12256 18955 12308 18964
rect 12256 18921 12265 18955
rect 12265 18921 12299 18955
rect 12299 18921 12308 18955
rect 12256 18912 12308 18921
rect 4988 18708 5040 18760
rect 3240 18615 3292 18624
rect 3240 18581 3249 18615
rect 3249 18581 3283 18615
rect 3283 18581 3292 18615
rect 3240 18572 3292 18581
rect 6184 18572 6236 18624
rect 8576 18819 8628 18828
rect 8576 18785 8585 18819
rect 8585 18785 8619 18819
rect 8619 18785 8628 18819
rect 9956 18887 10008 18896
rect 9956 18853 9965 18887
rect 9965 18853 9999 18887
rect 9999 18853 10008 18887
rect 9956 18844 10008 18853
rect 10876 18844 10928 18896
rect 11520 18844 11572 18896
rect 14832 18912 14884 18964
rect 8576 18776 8628 18785
rect 8392 18751 8444 18760
rect 8392 18717 8401 18751
rect 8401 18717 8435 18751
rect 8435 18717 8444 18751
rect 8392 18708 8444 18717
rect 8484 18751 8536 18760
rect 8484 18717 8493 18751
rect 8493 18717 8527 18751
rect 8527 18717 8536 18751
rect 8484 18708 8536 18717
rect 9404 18708 9456 18760
rect 8668 18640 8720 18692
rect 12900 18776 12952 18828
rect 13912 18819 13964 18828
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 13912 18785 13921 18819
rect 13921 18785 13955 18819
rect 13955 18785 13964 18819
rect 13912 18776 13964 18785
rect 9680 18572 9732 18624
rect 10600 18615 10652 18624
rect 10600 18581 10609 18615
rect 10609 18581 10643 18615
rect 10643 18581 10652 18615
rect 10600 18572 10652 18581
rect 14004 18640 14056 18692
rect 11428 18572 11480 18624
rect 11796 18615 11848 18624
rect 11796 18581 11805 18615
rect 11805 18581 11839 18615
rect 11839 18581 11848 18615
rect 11796 18572 11848 18581
rect 12164 18572 12216 18624
rect 12900 18615 12952 18624
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 13820 18615 13872 18624
rect 13820 18581 13829 18615
rect 13829 18581 13863 18615
rect 13863 18581 13872 18615
rect 13820 18572 13872 18581
rect 15568 18844 15620 18896
rect 16120 18776 16172 18828
rect 14556 18751 14608 18760
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 17500 18912 17552 18964
rect 17408 18844 17460 18896
rect 19432 18955 19484 18964
rect 19432 18921 19441 18955
rect 19441 18921 19475 18955
rect 19475 18921 19484 18955
rect 19432 18912 19484 18921
rect 19524 18912 19576 18964
rect 19800 18912 19852 18964
rect 18512 18776 18564 18828
rect 19156 18776 19208 18828
rect 16396 18751 16448 18760
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 16672 18751 16724 18760
rect 16672 18717 16681 18751
rect 16681 18717 16715 18751
rect 16715 18717 16724 18751
rect 16672 18708 16724 18717
rect 19800 18819 19852 18828
rect 19800 18785 19809 18819
rect 19809 18785 19843 18819
rect 19843 18785 19852 18819
rect 19800 18776 19852 18785
rect 20720 18912 20772 18964
rect 26056 18912 26108 18964
rect 27988 18912 28040 18964
rect 28908 18912 28960 18964
rect 29460 18912 29512 18964
rect 29552 18912 29604 18964
rect 20352 18776 20404 18828
rect 20996 18751 21048 18760
rect 20996 18717 21005 18751
rect 21005 18717 21039 18751
rect 21039 18717 21048 18751
rect 20996 18708 21048 18717
rect 23480 18751 23532 18760
rect 23480 18717 23489 18751
rect 23489 18717 23523 18751
rect 23523 18717 23532 18751
rect 23480 18708 23532 18717
rect 24124 18776 24176 18828
rect 25688 18776 25740 18828
rect 27712 18844 27764 18896
rect 28448 18844 28500 18896
rect 28816 18844 28868 18896
rect 27344 18776 27396 18828
rect 16764 18572 16816 18624
rect 17776 18572 17828 18624
rect 19524 18572 19576 18624
rect 23940 18640 23992 18692
rect 29000 18776 29052 18828
rect 29644 18844 29696 18896
rect 32496 18912 32548 18964
rect 30656 18844 30708 18896
rect 30012 18819 30064 18828
rect 30012 18785 30021 18819
rect 30021 18785 30055 18819
rect 30055 18785 30064 18819
rect 30012 18776 30064 18785
rect 30104 18819 30156 18828
rect 30104 18785 30113 18819
rect 30113 18785 30147 18819
rect 30147 18785 30156 18819
rect 30104 18776 30156 18785
rect 30288 18776 30340 18828
rect 32956 18776 33008 18828
rect 33508 18819 33560 18828
rect 33508 18785 33517 18819
rect 33517 18785 33551 18819
rect 33551 18785 33560 18819
rect 33508 18776 33560 18785
rect 29644 18751 29696 18760
rect 29644 18717 29653 18751
rect 29653 18717 29687 18751
rect 29687 18717 29696 18751
rect 29644 18708 29696 18717
rect 27896 18640 27948 18692
rect 29828 18640 29880 18692
rect 21364 18615 21416 18624
rect 21364 18581 21373 18615
rect 21373 18581 21407 18615
rect 21407 18581 21416 18615
rect 21364 18572 21416 18581
rect 21640 18572 21692 18624
rect 23388 18572 23440 18624
rect 24400 18572 24452 18624
rect 27436 18572 27488 18624
rect 28172 18572 28224 18624
rect 28816 18572 28868 18624
rect 29920 18572 29972 18624
rect 34520 18708 34572 18760
rect 30840 18615 30892 18624
rect 30840 18581 30849 18615
rect 30849 18581 30883 18615
rect 30883 18581 30892 18615
rect 30840 18572 30892 18581
rect 32036 18615 32088 18624
rect 32036 18581 32045 18615
rect 32045 18581 32079 18615
rect 32079 18581 32088 18615
rect 32036 18572 32088 18581
rect 6550 18470 6602 18522
rect 6614 18470 6666 18522
rect 6678 18470 6730 18522
rect 6742 18470 6794 18522
rect 6806 18470 6858 18522
rect 14439 18470 14491 18522
rect 14503 18470 14555 18522
rect 14567 18470 14619 18522
rect 14631 18470 14683 18522
rect 14695 18470 14747 18522
rect 22328 18470 22380 18522
rect 22392 18470 22444 18522
rect 22456 18470 22508 18522
rect 22520 18470 22572 18522
rect 22584 18470 22636 18522
rect 30217 18470 30269 18522
rect 30281 18470 30333 18522
rect 30345 18470 30397 18522
rect 30409 18470 30461 18522
rect 30473 18470 30525 18522
rect 3240 18368 3292 18420
rect 3608 18368 3660 18420
rect 6552 18368 6604 18420
rect 8576 18368 8628 18420
rect 11796 18368 11848 18420
rect 13820 18368 13872 18420
rect 14004 18368 14056 18420
rect 5724 18275 5776 18284
rect 5724 18241 5733 18275
rect 5733 18241 5767 18275
rect 5767 18241 5776 18275
rect 5724 18232 5776 18241
rect 5816 18232 5868 18284
rect 6552 18275 6604 18284
rect 6552 18241 6586 18275
rect 6586 18241 6604 18275
rect 6552 18232 6604 18241
rect 4712 18164 4764 18216
rect 5080 18164 5132 18216
rect 5264 18096 5316 18148
rect 3424 18071 3476 18080
rect 3424 18037 3433 18071
rect 3433 18037 3467 18071
rect 3467 18037 3476 18071
rect 3424 18028 3476 18037
rect 7656 18164 7708 18216
rect 8852 18232 8904 18284
rect 10600 18232 10652 18284
rect 10784 18232 10836 18284
rect 13084 18232 13136 18284
rect 14924 18368 14976 18420
rect 16672 18368 16724 18420
rect 6000 18028 6052 18080
rect 6368 18028 6420 18080
rect 8024 18096 8076 18148
rect 7748 18028 7800 18080
rect 9128 18071 9180 18080
rect 9128 18037 9137 18071
rect 9137 18037 9171 18071
rect 9171 18037 9180 18071
rect 9128 18028 9180 18037
rect 9772 18028 9824 18080
rect 10876 18071 10928 18080
rect 10876 18037 10885 18071
rect 10885 18037 10919 18071
rect 10919 18037 10928 18071
rect 10876 18028 10928 18037
rect 13820 18096 13872 18148
rect 12900 18028 12952 18080
rect 12992 18028 13044 18080
rect 16304 18232 16356 18284
rect 17316 18275 17368 18284
rect 17316 18241 17325 18275
rect 17325 18241 17359 18275
rect 17359 18241 17368 18275
rect 17316 18232 17368 18241
rect 17776 18275 17828 18284
rect 17776 18241 17794 18275
rect 17794 18241 17828 18275
rect 17776 18232 17828 18241
rect 17868 18275 17920 18284
rect 17868 18241 17877 18275
rect 17877 18241 17911 18275
rect 17911 18241 17920 18275
rect 17868 18232 17920 18241
rect 16764 18164 16816 18216
rect 16948 18164 17000 18216
rect 19064 18411 19116 18420
rect 19064 18377 19073 18411
rect 19073 18377 19107 18411
rect 19107 18377 19116 18411
rect 19064 18368 19116 18377
rect 23480 18368 23532 18420
rect 18788 18300 18840 18352
rect 19800 18300 19852 18352
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 19064 18232 19116 18284
rect 20260 18232 20312 18284
rect 20812 18232 20864 18284
rect 23572 18275 23624 18284
rect 23572 18241 23581 18275
rect 23581 18241 23615 18275
rect 23615 18241 23624 18275
rect 23572 18232 23624 18241
rect 18512 18207 18564 18216
rect 18512 18173 18521 18207
rect 18521 18173 18555 18207
rect 18555 18173 18564 18207
rect 18512 18164 18564 18173
rect 18604 18207 18656 18216
rect 18604 18173 18613 18207
rect 18613 18173 18647 18207
rect 18647 18173 18656 18207
rect 18604 18164 18656 18173
rect 18788 18207 18840 18216
rect 18788 18173 18797 18207
rect 18797 18173 18831 18207
rect 18831 18173 18840 18207
rect 18788 18164 18840 18173
rect 18972 18207 19024 18216
rect 18972 18173 18981 18207
rect 18981 18173 19015 18207
rect 19015 18173 19024 18207
rect 18972 18164 19024 18173
rect 24400 18232 24452 18284
rect 25688 18368 25740 18420
rect 27804 18368 27856 18420
rect 28356 18368 28408 18420
rect 27528 18300 27580 18352
rect 28080 18300 28132 18352
rect 26608 18207 26660 18216
rect 26608 18173 26617 18207
rect 26617 18173 26651 18207
rect 26651 18173 26660 18207
rect 26608 18164 26660 18173
rect 26792 18207 26844 18216
rect 26792 18173 26801 18207
rect 26801 18173 26835 18207
rect 26835 18173 26844 18207
rect 26792 18164 26844 18173
rect 21548 18139 21600 18148
rect 21548 18105 21557 18139
rect 21557 18105 21591 18139
rect 21591 18105 21600 18139
rect 21548 18096 21600 18105
rect 23480 18096 23532 18148
rect 27436 18164 27488 18216
rect 28448 18207 28500 18216
rect 28448 18173 28458 18207
rect 28458 18173 28500 18207
rect 28448 18164 28500 18173
rect 29276 18368 29328 18420
rect 30748 18368 30800 18420
rect 29368 18300 29420 18352
rect 29828 18300 29880 18352
rect 31208 18300 31260 18352
rect 28908 18232 28960 18284
rect 29644 18164 29696 18216
rect 30104 18164 30156 18216
rect 30840 18164 30892 18216
rect 31300 18164 31352 18216
rect 32956 18207 33008 18216
rect 32956 18173 32965 18207
rect 32965 18173 32999 18207
rect 32999 18173 33008 18207
rect 32956 18164 33008 18173
rect 33508 18275 33560 18284
rect 33508 18241 33517 18275
rect 33517 18241 33551 18275
rect 33551 18241 33560 18275
rect 33508 18232 33560 18241
rect 33692 18275 33744 18284
rect 33692 18241 33701 18275
rect 33701 18241 33735 18275
rect 33735 18241 33744 18275
rect 33692 18232 33744 18241
rect 27988 18096 28040 18148
rect 17132 18071 17184 18080
rect 17132 18037 17141 18071
rect 17141 18037 17175 18071
rect 17175 18037 17184 18071
rect 17132 18028 17184 18037
rect 17224 18028 17276 18080
rect 17684 18028 17736 18080
rect 18052 18028 18104 18080
rect 18604 18028 18656 18080
rect 20536 18071 20588 18080
rect 20536 18037 20545 18071
rect 20545 18037 20579 18071
rect 20579 18037 20588 18071
rect 20536 18028 20588 18037
rect 22192 18028 22244 18080
rect 24952 18071 25004 18080
rect 24952 18037 24961 18071
rect 24961 18037 24995 18071
rect 24995 18037 25004 18071
rect 24952 18028 25004 18037
rect 26884 18071 26936 18080
rect 26884 18037 26893 18071
rect 26893 18037 26927 18071
rect 26927 18037 26936 18071
rect 26884 18028 26936 18037
rect 26976 18028 27028 18080
rect 27068 18028 27120 18080
rect 29368 18096 29420 18148
rect 29552 18096 29604 18148
rect 30564 18096 30616 18148
rect 28448 18028 28500 18080
rect 28724 18071 28776 18080
rect 28724 18037 28733 18071
rect 28733 18037 28767 18071
rect 28767 18037 28776 18071
rect 28724 18028 28776 18037
rect 28816 18028 28868 18080
rect 29460 18028 29512 18080
rect 29920 18028 29972 18080
rect 30104 18071 30156 18080
rect 30104 18037 30113 18071
rect 30113 18037 30147 18071
rect 30147 18037 30156 18071
rect 30104 18028 30156 18037
rect 32036 18096 32088 18148
rect 32404 18096 32456 18148
rect 33600 18028 33652 18080
rect 7210 17926 7262 17978
rect 7274 17926 7326 17978
rect 7338 17926 7390 17978
rect 7402 17926 7454 17978
rect 7466 17926 7518 17978
rect 15099 17926 15151 17978
rect 15163 17926 15215 17978
rect 15227 17926 15279 17978
rect 15291 17926 15343 17978
rect 15355 17926 15407 17978
rect 22988 17926 23040 17978
rect 23052 17926 23104 17978
rect 23116 17926 23168 17978
rect 23180 17926 23232 17978
rect 23244 17926 23296 17978
rect 30877 17926 30929 17978
rect 30941 17926 30993 17978
rect 31005 17926 31057 17978
rect 31069 17926 31121 17978
rect 31133 17926 31185 17978
rect 5448 17824 5500 17876
rect 6920 17799 6972 17808
rect 6920 17765 6929 17799
rect 6929 17765 6963 17799
rect 6963 17765 6972 17799
rect 6920 17756 6972 17765
rect 9128 17824 9180 17876
rect 9588 17756 9640 17808
rect 18880 17824 18932 17876
rect 20904 17824 20956 17876
rect 12900 17799 12952 17808
rect 12900 17765 12909 17799
rect 12909 17765 12943 17799
rect 12943 17765 12952 17799
rect 12900 17756 12952 17765
rect 13452 17799 13504 17808
rect 13452 17765 13461 17799
rect 13461 17765 13495 17799
rect 13495 17765 13504 17799
rect 13452 17756 13504 17765
rect 16028 17799 16080 17808
rect 16028 17765 16037 17799
rect 16037 17765 16071 17799
rect 16071 17765 16080 17799
rect 16028 17756 16080 17765
rect 16120 17756 16172 17808
rect 17408 17756 17460 17808
rect 17776 17799 17828 17808
rect 17776 17765 17785 17799
rect 17785 17765 17819 17799
rect 17819 17765 17828 17799
rect 17776 17756 17828 17765
rect 17868 17756 17920 17808
rect 3424 17688 3476 17740
rect 5356 17688 5408 17740
rect 4528 17663 4580 17672
rect 4528 17629 4537 17663
rect 4537 17629 4571 17663
rect 4571 17629 4580 17663
rect 4528 17620 4580 17629
rect 3056 17527 3108 17536
rect 3056 17493 3065 17527
rect 3065 17493 3099 17527
rect 3099 17493 3108 17527
rect 3056 17484 3108 17493
rect 4160 17484 4212 17536
rect 6368 17620 6420 17672
rect 6460 17484 6512 17536
rect 7104 17595 7156 17604
rect 7104 17561 7113 17595
rect 7113 17561 7147 17595
rect 7147 17561 7156 17595
rect 12256 17663 12308 17672
rect 12256 17629 12265 17663
rect 12265 17629 12299 17663
rect 12299 17629 12308 17663
rect 12256 17620 12308 17629
rect 12348 17620 12400 17672
rect 12992 17688 13044 17740
rect 13084 17688 13136 17740
rect 14832 17620 14884 17672
rect 16580 17620 16632 17672
rect 16856 17620 16908 17672
rect 17224 17663 17276 17672
rect 17224 17629 17233 17663
rect 17233 17629 17267 17663
rect 17267 17629 17276 17663
rect 17224 17620 17276 17629
rect 17592 17620 17644 17672
rect 20812 17756 20864 17808
rect 21916 17756 21968 17808
rect 22744 17824 22796 17876
rect 23296 17824 23348 17876
rect 18236 17688 18288 17740
rect 18328 17620 18380 17672
rect 19064 17688 19116 17740
rect 19524 17731 19576 17740
rect 19524 17697 19533 17731
rect 19533 17697 19567 17731
rect 19567 17697 19576 17731
rect 19524 17688 19576 17697
rect 20536 17688 20588 17740
rect 21272 17688 21324 17740
rect 21640 17688 21692 17740
rect 24216 17756 24268 17808
rect 26884 17824 26936 17876
rect 28264 17824 28316 17876
rect 28080 17756 28132 17808
rect 27620 17688 27672 17740
rect 28264 17688 28316 17740
rect 29368 17824 29420 17876
rect 30104 17824 30156 17876
rect 32404 17824 32456 17876
rect 33508 17824 33560 17876
rect 28540 17688 28592 17740
rect 7104 17552 7156 17561
rect 7656 17484 7708 17536
rect 9772 17527 9824 17536
rect 9772 17493 9781 17527
rect 9781 17493 9815 17527
rect 9815 17493 9824 17527
rect 9772 17484 9824 17493
rect 10508 17484 10560 17536
rect 11060 17484 11112 17536
rect 15476 17484 15528 17536
rect 17684 17552 17736 17604
rect 19248 17620 19300 17672
rect 20076 17620 20128 17672
rect 20260 17663 20312 17672
rect 20260 17629 20269 17663
rect 20269 17629 20303 17663
rect 20303 17629 20312 17663
rect 20260 17620 20312 17629
rect 16672 17484 16724 17536
rect 17132 17484 17184 17536
rect 17868 17484 17920 17536
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 18420 17484 18472 17536
rect 19800 17527 19852 17536
rect 19800 17493 19809 17527
rect 19809 17493 19843 17527
rect 19843 17493 19852 17527
rect 19800 17484 19852 17493
rect 23020 17620 23072 17672
rect 24952 17620 25004 17672
rect 20996 17484 21048 17536
rect 21272 17484 21324 17536
rect 23480 17484 23532 17536
rect 25228 17527 25280 17536
rect 25228 17493 25237 17527
rect 25237 17493 25271 17527
rect 25271 17493 25280 17527
rect 25228 17484 25280 17493
rect 27620 17484 27672 17536
rect 28540 17484 28592 17536
rect 28632 17527 28684 17536
rect 28632 17493 28641 17527
rect 28641 17493 28675 17527
rect 28675 17493 28684 17527
rect 28632 17484 28684 17493
rect 29184 17663 29236 17672
rect 29184 17629 29193 17663
rect 29193 17629 29227 17663
rect 29227 17629 29236 17663
rect 29184 17620 29236 17629
rect 29368 17731 29420 17740
rect 29368 17697 29377 17731
rect 29377 17697 29411 17731
rect 29411 17697 29420 17731
rect 29368 17688 29420 17697
rect 29920 17688 29972 17740
rect 30656 17756 30708 17808
rect 29644 17620 29696 17672
rect 29828 17620 29880 17672
rect 31208 17731 31260 17740
rect 31208 17697 31217 17731
rect 31217 17697 31251 17731
rect 31251 17697 31260 17731
rect 31208 17688 31260 17697
rect 33140 17688 33192 17740
rect 30656 17620 30708 17672
rect 28908 17552 28960 17604
rect 32128 17663 32180 17672
rect 32128 17629 32137 17663
rect 32137 17629 32171 17663
rect 32171 17629 32180 17663
rect 32128 17620 32180 17629
rect 29460 17484 29512 17536
rect 29552 17527 29604 17536
rect 29552 17493 29561 17527
rect 29561 17493 29595 17527
rect 29595 17493 29604 17527
rect 29552 17484 29604 17493
rect 30748 17484 30800 17536
rect 31024 17527 31076 17536
rect 31024 17493 31033 17527
rect 31033 17493 31067 17527
rect 31067 17493 31076 17527
rect 31024 17484 31076 17493
rect 6550 17382 6602 17434
rect 6614 17382 6666 17434
rect 6678 17382 6730 17434
rect 6742 17382 6794 17434
rect 6806 17382 6858 17434
rect 14439 17382 14491 17434
rect 14503 17382 14555 17434
rect 14567 17382 14619 17434
rect 14631 17382 14683 17434
rect 14695 17382 14747 17434
rect 22328 17382 22380 17434
rect 22392 17382 22444 17434
rect 22456 17382 22508 17434
rect 22520 17382 22572 17434
rect 22584 17382 22636 17434
rect 30217 17382 30269 17434
rect 30281 17382 30333 17434
rect 30345 17382 30397 17434
rect 30409 17382 30461 17434
rect 30473 17382 30525 17434
rect 3056 17280 3108 17332
rect 4344 17144 4396 17196
rect 5080 17187 5132 17196
rect 5080 17153 5089 17187
rect 5089 17153 5123 17187
rect 5123 17153 5132 17187
rect 5080 17144 5132 17153
rect 1308 17008 1360 17060
rect 6092 17280 6144 17332
rect 6368 17280 6420 17332
rect 9588 17323 9640 17332
rect 9588 17289 9597 17323
rect 9597 17289 9631 17323
rect 9631 17289 9640 17323
rect 9588 17280 9640 17289
rect 6460 17212 6512 17264
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 6368 17144 6420 17196
rect 8208 17212 8260 17264
rect 12164 17280 12216 17332
rect 12256 17280 12308 17332
rect 13452 17280 13504 17332
rect 5908 17076 5960 17128
rect 10876 17187 10928 17196
rect 10876 17153 10885 17187
rect 10885 17153 10919 17187
rect 10919 17153 10928 17187
rect 10876 17144 10928 17153
rect 13728 17212 13780 17264
rect 15016 17280 15068 17332
rect 18328 17280 18380 17332
rect 18788 17280 18840 17332
rect 20260 17280 20312 17332
rect 21548 17280 21600 17332
rect 12900 17144 12952 17196
rect 14188 17144 14240 17196
rect 15476 17212 15528 17264
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 6276 17008 6328 17060
rect 6828 17119 6880 17128
rect 6828 17085 6837 17119
rect 6837 17085 6871 17119
rect 6871 17085 6880 17119
rect 6828 17076 6880 17085
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 10416 17076 10468 17128
rect 14832 17119 14884 17128
rect 4804 16940 4856 16992
rect 7748 17008 7800 17060
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 9864 16940 9916 16992
rect 10232 16940 10284 16992
rect 12808 17051 12860 17060
rect 12808 17017 12817 17051
rect 12817 17017 12851 17051
rect 12851 17017 12860 17051
rect 12808 17008 12860 17017
rect 13820 17008 13872 17060
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 15568 17119 15620 17128
rect 15568 17085 15577 17119
rect 15577 17085 15611 17119
rect 15611 17085 15620 17119
rect 15568 17076 15620 17085
rect 16396 17144 16448 17196
rect 18144 17187 18196 17196
rect 18144 17153 18178 17187
rect 18178 17153 18196 17187
rect 22836 17280 22888 17332
rect 25228 17280 25280 17332
rect 26608 17280 26660 17332
rect 18144 17144 18196 17153
rect 17592 17076 17644 17128
rect 17868 17076 17920 17128
rect 18328 17076 18380 17128
rect 18696 17187 18748 17196
rect 18696 17153 18705 17187
rect 18705 17153 18739 17187
rect 18739 17153 18748 17187
rect 18696 17144 18748 17153
rect 19800 17144 19852 17196
rect 22284 17212 22336 17264
rect 22376 17212 22428 17264
rect 26976 17255 27028 17264
rect 26976 17221 26985 17255
rect 26985 17221 27019 17255
rect 27019 17221 27028 17255
rect 26976 17212 27028 17221
rect 29644 17280 29696 17332
rect 31024 17280 31076 17332
rect 32128 17280 32180 17332
rect 22560 17144 22612 17196
rect 23020 17144 23072 17196
rect 18512 17076 18564 17128
rect 18604 17076 18656 17128
rect 18788 17076 18840 17128
rect 21272 17076 21324 17128
rect 21364 17076 21416 17128
rect 22192 17076 22244 17128
rect 22284 17076 22336 17128
rect 28632 17144 28684 17196
rect 24308 17119 24360 17128
rect 24308 17085 24317 17119
rect 24317 17085 24351 17119
rect 24351 17085 24360 17119
rect 24308 17076 24360 17085
rect 24400 17076 24452 17128
rect 25136 17119 25188 17128
rect 25136 17085 25145 17119
rect 25145 17085 25179 17119
rect 25179 17085 25188 17119
rect 25136 17076 25188 17085
rect 25872 17119 25924 17128
rect 25872 17085 25881 17119
rect 25881 17085 25915 17119
rect 25915 17085 25924 17119
rect 25872 17076 25924 17085
rect 15660 17008 15712 17060
rect 16028 17051 16080 17060
rect 16028 17017 16037 17051
rect 16037 17017 16071 17051
rect 16071 17017 16080 17051
rect 16028 17008 16080 17017
rect 13912 16940 13964 16992
rect 14188 16983 14240 16992
rect 14188 16949 14197 16983
rect 14197 16949 14231 16983
rect 14231 16949 14240 16983
rect 14188 16940 14240 16949
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 18144 16940 18196 16992
rect 23756 16983 23808 16992
rect 23756 16949 23765 16983
rect 23765 16949 23799 16983
rect 23799 16949 23808 16983
rect 23756 16940 23808 16949
rect 23848 16940 23900 16992
rect 25596 16940 25648 16992
rect 26332 16940 26384 16992
rect 27620 16940 27672 16992
rect 29736 17076 29788 17128
rect 32956 17187 33008 17196
rect 32956 17153 32965 17187
rect 32965 17153 32999 17187
rect 32999 17153 33008 17187
rect 32956 17144 33008 17153
rect 33600 17187 33652 17196
rect 33600 17153 33609 17187
rect 33609 17153 33643 17187
rect 33643 17153 33652 17187
rect 33600 17144 33652 17153
rect 29000 17008 29052 17060
rect 28908 16940 28960 16992
rect 29460 16940 29512 16992
rect 30564 16983 30616 16992
rect 30564 16949 30573 16983
rect 30573 16949 30607 16983
rect 30607 16949 30616 16983
rect 30564 16940 30616 16949
rect 32036 17008 32088 17060
rect 31300 16940 31352 16992
rect 7210 16838 7262 16890
rect 7274 16838 7326 16890
rect 7338 16838 7390 16890
rect 7402 16838 7454 16890
rect 7466 16838 7518 16890
rect 15099 16838 15151 16890
rect 15163 16838 15215 16890
rect 15227 16838 15279 16890
rect 15291 16838 15343 16890
rect 15355 16838 15407 16890
rect 22988 16838 23040 16890
rect 23052 16838 23104 16890
rect 23116 16838 23168 16890
rect 23180 16838 23232 16890
rect 23244 16838 23296 16890
rect 30877 16838 30929 16890
rect 30941 16838 30993 16890
rect 31005 16838 31057 16890
rect 31069 16838 31121 16890
rect 31133 16838 31185 16890
rect 4528 16736 4580 16788
rect 4804 16736 4856 16788
rect 5264 16736 5316 16788
rect 5356 16736 5408 16788
rect 6460 16736 6512 16788
rect 7748 16779 7800 16788
rect 7748 16745 7757 16779
rect 7757 16745 7791 16779
rect 7791 16745 7800 16779
rect 7748 16736 7800 16745
rect 9312 16736 9364 16788
rect 11152 16736 11204 16788
rect 4252 16643 4304 16652
rect 4252 16609 4261 16643
rect 4261 16609 4295 16643
rect 4295 16609 4304 16643
rect 4252 16600 4304 16609
rect 15844 16736 15896 16788
rect 15936 16779 15988 16788
rect 15936 16745 15945 16779
rect 15945 16745 15979 16779
rect 15979 16745 15988 16779
rect 15936 16736 15988 16745
rect 16120 16736 16172 16788
rect 16580 16736 16632 16788
rect 11060 16668 11112 16720
rect 11980 16668 12032 16720
rect 12164 16668 12216 16720
rect 14004 16668 14056 16720
rect 6092 16600 6144 16652
rect 8208 16600 8260 16652
rect 8484 16643 8536 16652
rect 8484 16609 8493 16643
rect 8493 16609 8527 16643
rect 8527 16609 8536 16643
rect 8484 16600 8536 16609
rect 4344 16575 4396 16584
rect 4344 16541 4353 16575
rect 4353 16541 4387 16575
rect 4387 16541 4396 16575
rect 4344 16532 4396 16541
rect 4528 16575 4580 16584
rect 4528 16541 4537 16575
rect 4537 16541 4571 16575
rect 4571 16541 4580 16575
rect 4528 16532 4580 16541
rect 8300 16575 8352 16584
rect 8300 16541 8309 16575
rect 8309 16541 8343 16575
rect 8343 16541 8352 16575
rect 8300 16532 8352 16541
rect 8668 16600 8720 16652
rect 9128 16532 9180 16584
rect 13084 16600 13136 16652
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 13544 16532 13596 16584
rect 15568 16668 15620 16720
rect 16488 16668 16540 16720
rect 18604 16736 18656 16788
rect 21640 16736 21692 16788
rect 22376 16779 22428 16788
rect 22376 16745 22385 16779
rect 22385 16745 22419 16779
rect 22419 16745 22428 16779
rect 22376 16736 22428 16745
rect 22836 16779 22888 16788
rect 22836 16745 22845 16779
rect 22845 16745 22879 16779
rect 22879 16745 22888 16779
rect 22836 16736 22888 16745
rect 23848 16736 23900 16788
rect 24216 16736 24268 16788
rect 24308 16736 24360 16788
rect 25872 16736 25924 16788
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 17592 16643 17644 16652
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 17592 16600 17644 16609
rect 19340 16600 19392 16652
rect 20812 16668 20864 16720
rect 22008 16600 22060 16652
rect 25044 16668 25096 16720
rect 15660 16575 15712 16584
rect 15660 16541 15669 16575
rect 15669 16541 15703 16575
rect 15703 16541 15712 16575
rect 15660 16532 15712 16541
rect 16764 16532 16816 16584
rect 13176 16464 13228 16516
rect 3240 16396 3292 16448
rect 7932 16396 7984 16448
rect 14924 16439 14976 16448
rect 14924 16405 14933 16439
rect 14933 16405 14967 16439
rect 14967 16405 14976 16439
rect 14924 16396 14976 16405
rect 16488 16396 16540 16448
rect 18144 16396 18196 16448
rect 18420 16396 18472 16448
rect 18788 16396 18840 16448
rect 20352 16439 20404 16448
rect 20352 16405 20361 16439
rect 20361 16405 20395 16439
rect 20395 16405 20404 16439
rect 20352 16396 20404 16405
rect 20720 16396 20772 16448
rect 22560 16396 22612 16448
rect 22836 16396 22888 16448
rect 23480 16600 23532 16652
rect 23848 16643 23900 16652
rect 23848 16609 23857 16643
rect 23857 16609 23891 16643
rect 23891 16609 23900 16643
rect 23848 16600 23900 16609
rect 23388 16532 23440 16584
rect 24400 16600 24452 16652
rect 25596 16643 25648 16652
rect 25596 16609 25605 16643
rect 25605 16609 25639 16643
rect 25639 16609 25648 16643
rect 25596 16600 25648 16609
rect 26332 16643 26384 16652
rect 26332 16609 26341 16643
rect 26341 16609 26375 16643
rect 26375 16609 26384 16643
rect 26332 16600 26384 16609
rect 26424 16643 26476 16652
rect 26424 16609 26433 16643
rect 26433 16609 26467 16643
rect 26467 16609 26476 16643
rect 26424 16600 26476 16609
rect 26516 16600 26568 16652
rect 26608 16643 26660 16652
rect 26608 16609 26617 16643
rect 26617 16609 26651 16643
rect 26651 16609 26660 16643
rect 26608 16600 26660 16609
rect 27528 16643 27580 16652
rect 27528 16609 27537 16643
rect 27537 16609 27571 16643
rect 27571 16609 27580 16643
rect 27528 16600 27580 16609
rect 27620 16600 27672 16652
rect 27712 16600 27764 16652
rect 28172 16736 28224 16788
rect 28356 16736 28408 16788
rect 29552 16736 29604 16788
rect 29736 16779 29788 16788
rect 29736 16745 29745 16779
rect 29745 16745 29779 16779
rect 29779 16745 29788 16779
rect 29736 16736 29788 16745
rect 29828 16779 29880 16788
rect 29828 16745 29837 16779
rect 29837 16745 29871 16779
rect 29871 16745 29880 16779
rect 29828 16736 29880 16745
rect 30104 16736 30156 16788
rect 30656 16736 30708 16788
rect 31300 16736 31352 16788
rect 23572 16464 23624 16516
rect 26332 16464 26384 16516
rect 28540 16532 28592 16584
rect 28724 16643 28776 16652
rect 28724 16609 28733 16643
rect 28733 16609 28767 16643
rect 28767 16609 28776 16643
rect 28724 16600 28776 16609
rect 30196 16668 30248 16720
rect 30564 16711 30616 16720
rect 30564 16677 30573 16711
rect 30573 16677 30607 16711
rect 30607 16677 30616 16711
rect 30564 16668 30616 16677
rect 29736 16600 29788 16652
rect 29920 16600 29972 16652
rect 30748 16600 30800 16652
rect 29184 16532 29236 16584
rect 27896 16464 27948 16516
rect 29644 16464 29696 16516
rect 30472 16532 30524 16584
rect 30196 16507 30248 16516
rect 30196 16473 30205 16507
rect 30205 16473 30239 16507
rect 30239 16473 30248 16507
rect 30196 16464 30248 16473
rect 33048 16575 33100 16584
rect 33048 16541 33057 16575
rect 33057 16541 33091 16575
rect 33091 16541 33100 16575
rect 33048 16532 33100 16541
rect 28724 16396 28776 16448
rect 29828 16396 29880 16448
rect 6550 16294 6602 16346
rect 6614 16294 6666 16346
rect 6678 16294 6730 16346
rect 6742 16294 6794 16346
rect 6806 16294 6858 16346
rect 14439 16294 14491 16346
rect 14503 16294 14555 16346
rect 14567 16294 14619 16346
rect 14631 16294 14683 16346
rect 14695 16294 14747 16346
rect 22328 16294 22380 16346
rect 22392 16294 22444 16346
rect 22456 16294 22508 16346
rect 22520 16294 22572 16346
rect 22584 16294 22636 16346
rect 30217 16294 30269 16346
rect 30281 16294 30333 16346
rect 30345 16294 30397 16346
rect 30409 16294 30461 16346
rect 30473 16294 30525 16346
rect 4344 16192 4396 16244
rect 6368 16192 6420 16244
rect 11060 16124 11112 16176
rect 13176 16235 13228 16244
rect 13176 16201 13185 16235
rect 13185 16201 13219 16235
rect 13219 16201 13228 16235
rect 13176 16192 13228 16201
rect 14004 16235 14056 16244
rect 14004 16201 14013 16235
rect 14013 16201 14047 16235
rect 14047 16201 14056 16235
rect 14004 16192 14056 16201
rect 16028 16235 16080 16244
rect 16028 16201 16037 16235
rect 16037 16201 16071 16235
rect 16071 16201 16080 16235
rect 16028 16192 16080 16201
rect 16764 16235 16816 16244
rect 16764 16201 16773 16235
rect 16773 16201 16807 16235
rect 16807 16201 16816 16235
rect 16764 16192 16816 16201
rect 17684 16192 17736 16244
rect 23572 16192 23624 16244
rect 24584 16192 24636 16244
rect 15660 16124 15712 16176
rect 20812 16124 20864 16176
rect 4068 16056 4120 16108
rect 3056 16031 3108 16040
rect 3056 15997 3065 16031
rect 3065 15997 3099 16031
rect 3099 15997 3108 16031
rect 3056 15988 3108 15997
rect 5264 16056 5316 16108
rect 6460 16056 6512 16108
rect 13084 16099 13136 16108
rect 13084 16065 13093 16099
rect 13093 16065 13127 16099
rect 13127 16065 13136 16099
rect 13084 16056 13136 16065
rect 13820 16099 13872 16108
rect 13820 16065 13829 16099
rect 13829 16065 13863 16099
rect 13863 16065 13872 16099
rect 13820 16056 13872 16065
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 3240 15920 3292 15972
rect 5908 15920 5960 15972
rect 6920 15963 6972 15972
rect 6920 15929 6929 15963
rect 6929 15929 6963 15963
rect 6963 15929 6972 15963
rect 6920 15920 6972 15929
rect 9680 15920 9732 15972
rect 10140 15963 10192 15972
rect 10140 15929 10149 15963
rect 10149 15929 10183 15963
rect 10183 15929 10192 15963
rect 10140 15920 10192 15929
rect 10508 15988 10560 16040
rect 11336 16031 11388 16040
rect 11336 15997 11345 16031
rect 11345 15997 11379 16031
rect 11379 15997 11388 16031
rect 11336 15988 11388 15997
rect 13912 16031 13964 16040
rect 13912 15997 13921 16031
rect 13921 15997 13955 16031
rect 13955 15997 13964 16031
rect 13912 15988 13964 15997
rect 5448 15895 5500 15904
rect 5448 15861 5457 15895
rect 5457 15861 5491 15895
rect 5491 15861 5500 15895
rect 5448 15852 5500 15861
rect 5632 15852 5684 15904
rect 6276 15852 6328 15904
rect 9772 15852 9824 15904
rect 10232 15852 10284 15904
rect 10600 15895 10652 15904
rect 10600 15861 10609 15895
rect 10609 15861 10643 15895
rect 10643 15861 10652 15895
rect 10600 15852 10652 15861
rect 13176 15920 13228 15972
rect 12992 15852 13044 15904
rect 16580 16099 16632 16108
rect 16580 16065 16589 16099
rect 16589 16065 16623 16099
rect 16623 16065 16632 16099
rect 16580 16056 16632 16065
rect 17500 16056 17552 16108
rect 18420 16056 18472 16108
rect 21916 16056 21968 16108
rect 23756 16056 23808 16108
rect 25044 16192 25096 16244
rect 28908 16192 28960 16244
rect 29920 16192 29972 16244
rect 32036 16235 32088 16244
rect 32036 16201 32045 16235
rect 32045 16201 32079 16235
rect 32079 16201 32088 16235
rect 32036 16192 32088 16201
rect 26056 16124 26108 16176
rect 28448 16124 28500 16176
rect 29644 16099 29696 16108
rect 17040 15988 17092 16040
rect 19248 15988 19300 16040
rect 19800 15988 19852 16040
rect 20352 15988 20404 16040
rect 20444 15988 20496 16040
rect 16764 15920 16816 15972
rect 15476 15852 15528 15904
rect 16212 15852 16264 15904
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 19892 15852 19944 15904
rect 20904 16031 20956 16040
rect 20904 15997 20913 16031
rect 20913 15997 20947 16031
rect 20947 15997 20956 16031
rect 20904 15988 20956 15997
rect 24952 15988 25004 16040
rect 26700 16031 26752 16040
rect 23756 15920 23808 15972
rect 24400 15920 24452 15972
rect 26700 15997 26709 16031
rect 26709 15997 26743 16031
rect 26743 15997 26752 16031
rect 26700 15988 26752 15997
rect 26332 15920 26384 15972
rect 29644 16065 29653 16099
rect 29653 16065 29687 16099
rect 29687 16065 29696 16099
rect 29644 16056 29696 16065
rect 29920 16056 29972 16108
rect 27344 16031 27396 16040
rect 27344 15997 27353 16031
rect 27353 15997 27387 16031
rect 27387 15997 27396 16031
rect 27344 15988 27396 15997
rect 28724 15988 28776 16040
rect 28816 15988 28868 16040
rect 21180 15852 21232 15904
rect 21456 15852 21508 15904
rect 21640 15852 21692 15904
rect 24032 15852 24084 15904
rect 25136 15852 25188 15904
rect 26148 15852 26200 15904
rect 28816 15852 28868 15904
rect 31944 15988 31996 16040
rect 32036 15988 32088 16040
rect 33140 16056 33192 16108
rect 33600 15988 33652 16040
rect 29368 15852 29420 15904
rect 30564 15852 30616 15904
rect 34888 15920 34940 15972
rect 32404 15895 32456 15904
rect 32404 15861 32413 15895
rect 32413 15861 32447 15895
rect 32447 15861 32456 15895
rect 32404 15852 32456 15861
rect 7210 15750 7262 15802
rect 7274 15750 7326 15802
rect 7338 15750 7390 15802
rect 7402 15750 7454 15802
rect 7466 15750 7518 15802
rect 15099 15750 15151 15802
rect 15163 15750 15215 15802
rect 15227 15750 15279 15802
rect 15291 15750 15343 15802
rect 15355 15750 15407 15802
rect 22988 15750 23040 15802
rect 23052 15750 23104 15802
rect 23116 15750 23168 15802
rect 23180 15750 23232 15802
rect 23244 15750 23296 15802
rect 30877 15750 30929 15802
rect 30941 15750 30993 15802
rect 31005 15750 31057 15802
rect 31069 15750 31121 15802
rect 31133 15750 31185 15802
rect 4252 15648 4304 15700
rect 1308 15580 1360 15632
rect 4712 15623 4764 15632
rect 4712 15589 4721 15623
rect 4721 15589 4755 15623
rect 4755 15589 4764 15623
rect 4712 15580 4764 15589
rect 4344 15555 4396 15564
rect 4344 15521 4353 15555
rect 4353 15521 4387 15555
rect 4387 15521 4396 15555
rect 4344 15512 4396 15521
rect 5448 15648 5500 15700
rect 6920 15648 6972 15700
rect 5816 15623 5868 15632
rect 5816 15589 5825 15623
rect 5825 15589 5859 15623
rect 5859 15589 5868 15623
rect 7564 15648 7616 15700
rect 7932 15648 7984 15700
rect 9128 15648 9180 15700
rect 9680 15648 9732 15700
rect 10140 15648 10192 15700
rect 11336 15648 11388 15700
rect 11980 15691 12032 15700
rect 11980 15657 11989 15691
rect 11989 15657 12023 15691
rect 12023 15657 12032 15691
rect 11980 15648 12032 15657
rect 5816 15580 5868 15589
rect 7748 15580 7800 15632
rect 11152 15580 11204 15632
rect 13636 15648 13688 15700
rect 15752 15648 15804 15700
rect 18144 15648 18196 15700
rect 19248 15648 19300 15700
rect 20536 15648 20588 15700
rect 20720 15648 20772 15700
rect 22008 15648 22060 15700
rect 23756 15648 23808 15700
rect 24032 15648 24084 15700
rect 27344 15648 27396 15700
rect 5632 15555 5684 15564
rect 5632 15521 5641 15555
rect 5641 15521 5675 15555
rect 5675 15521 5684 15555
rect 5632 15512 5684 15521
rect 6276 15512 6328 15564
rect 5724 15376 5776 15428
rect 9772 15512 9824 15564
rect 10324 15512 10376 15564
rect 8852 15487 8904 15496
rect 8852 15453 8861 15487
rect 8861 15453 8895 15487
rect 8895 15453 8904 15487
rect 8852 15444 8904 15453
rect 9036 15444 9088 15496
rect 10416 15444 10468 15496
rect 6368 15308 6420 15360
rect 7012 15308 7064 15360
rect 11520 15376 11572 15428
rect 13176 15580 13228 15632
rect 13728 15580 13780 15632
rect 14740 15580 14792 15632
rect 15476 15580 15528 15632
rect 13084 15512 13136 15564
rect 16120 15512 16172 15564
rect 17408 15580 17460 15632
rect 17684 15580 17736 15632
rect 12164 15444 12216 15496
rect 12808 15444 12860 15496
rect 13912 15444 13964 15496
rect 7380 15308 7432 15360
rect 8024 15308 8076 15360
rect 11060 15308 11112 15360
rect 11152 15351 11204 15360
rect 11152 15317 11161 15351
rect 11161 15317 11195 15351
rect 11195 15317 11204 15351
rect 13452 15376 13504 15428
rect 15844 15444 15896 15496
rect 18052 15512 18104 15564
rect 18880 15555 18932 15564
rect 18880 15521 18889 15555
rect 18889 15521 18923 15555
rect 18923 15521 18932 15555
rect 26700 15580 26752 15632
rect 18880 15512 18932 15521
rect 22192 15512 22244 15564
rect 23480 15512 23532 15564
rect 23756 15555 23808 15564
rect 23756 15521 23765 15555
rect 23765 15521 23799 15555
rect 23799 15521 23808 15555
rect 23756 15512 23808 15521
rect 27436 15555 27488 15564
rect 27436 15521 27445 15555
rect 27445 15521 27479 15555
rect 27479 15521 27488 15555
rect 27436 15512 27488 15521
rect 27988 15580 28040 15632
rect 29000 15580 29052 15632
rect 30564 15580 30616 15632
rect 31300 15580 31352 15632
rect 32404 15648 32456 15700
rect 32956 15648 33008 15700
rect 28632 15555 28684 15564
rect 28632 15521 28641 15555
rect 28641 15521 28675 15555
rect 28675 15521 28684 15555
rect 28632 15512 28684 15521
rect 17040 15444 17092 15496
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 17224 15444 17276 15453
rect 19340 15487 19392 15496
rect 19340 15453 19349 15487
rect 19349 15453 19383 15487
rect 19383 15453 19392 15487
rect 19340 15444 19392 15453
rect 19432 15444 19484 15496
rect 20168 15444 20220 15496
rect 20628 15444 20680 15496
rect 20904 15444 20956 15496
rect 27896 15444 27948 15496
rect 28908 15487 28960 15496
rect 28908 15453 28917 15487
rect 28917 15453 28951 15487
rect 28951 15453 28960 15487
rect 28908 15444 28960 15453
rect 11152 15308 11204 15317
rect 13176 15308 13228 15360
rect 14280 15308 14332 15360
rect 16488 15308 16540 15360
rect 16764 15308 16816 15360
rect 19892 15376 19944 15428
rect 26608 15376 26660 15428
rect 26976 15376 27028 15428
rect 29920 15512 29972 15564
rect 18880 15308 18932 15360
rect 19984 15351 20036 15360
rect 19984 15317 19993 15351
rect 19993 15317 20027 15351
rect 20027 15317 20036 15351
rect 19984 15308 20036 15317
rect 21824 15351 21876 15360
rect 21824 15317 21833 15351
rect 21833 15317 21867 15351
rect 21867 15317 21876 15351
rect 21824 15308 21876 15317
rect 23388 15308 23440 15360
rect 27160 15308 27212 15360
rect 28080 15308 28132 15360
rect 31944 15376 31996 15428
rect 31852 15308 31904 15360
rect 33140 15512 33192 15564
rect 33876 15351 33928 15360
rect 33876 15317 33885 15351
rect 33885 15317 33919 15351
rect 33919 15317 33928 15351
rect 33876 15308 33928 15317
rect 6550 15206 6602 15258
rect 6614 15206 6666 15258
rect 6678 15206 6730 15258
rect 6742 15206 6794 15258
rect 6806 15206 6858 15258
rect 14439 15206 14491 15258
rect 14503 15206 14555 15258
rect 14567 15206 14619 15258
rect 14631 15206 14683 15258
rect 14695 15206 14747 15258
rect 22328 15206 22380 15258
rect 22392 15206 22444 15258
rect 22456 15206 22508 15258
rect 22520 15206 22572 15258
rect 22584 15206 22636 15258
rect 30217 15206 30269 15258
rect 30281 15206 30333 15258
rect 30345 15206 30397 15258
rect 30409 15206 30461 15258
rect 30473 15206 30525 15258
rect 5264 15104 5316 15156
rect 5816 15104 5868 15156
rect 5908 15104 5960 15156
rect 6276 15104 6328 15156
rect 7012 15104 7064 15156
rect 5080 15036 5132 15088
rect 5724 15079 5776 15088
rect 5724 15045 5733 15079
rect 5733 15045 5767 15079
rect 5767 15045 5776 15079
rect 5724 15036 5776 15045
rect 4344 15011 4396 15020
rect 4344 14977 4353 15011
rect 4353 14977 4387 15011
rect 4387 14977 4396 15011
rect 4344 14968 4396 14977
rect 4436 14968 4488 15020
rect 5356 14968 5408 15020
rect 7840 15147 7892 15156
rect 7840 15113 7849 15147
rect 7849 15113 7883 15147
rect 7883 15113 7892 15147
rect 7840 15104 7892 15113
rect 8208 15104 8260 15156
rect 8300 15104 8352 15156
rect 10416 15104 10468 15156
rect 11060 15147 11112 15156
rect 11060 15113 11069 15147
rect 11069 15113 11103 15147
rect 11103 15113 11112 15147
rect 11060 15104 11112 15113
rect 14832 15147 14884 15156
rect 14832 15113 14841 15147
rect 14841 15113 14875 15147
rect 14875 15113 14884 15147
rect 14832 15104 14884 15113
rect 7748 15036 7800 15088
rect 11336 15036 11388 15088
rect 5172 14900 5224 14952
rect 6276 14900 6328 14952
rect 4160 14807 4212 14816
rect 4160 14773 4169 14807
rect 4169 14773 4203 14807
rect 4203 14773 4212 14807
rect 4160 14764 4212 14773
rect 6920 14807 6972 14816
rect 6920 14773 6929 14807
rect 6929 14773 6963 14807
rect 6963 14773 6972 14807
rect 6920 14764 6972 14773
rect 7564 14832 7616 14884
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 8760 14832 8812 14884
rect 9956 14968 10008 15020
rect 11152 14968 11204 15020
rect 13268 14968 13320 15020
rect 13912 15011 13964 15020
rect 13912 14977 13921 15011
rect 13921 14977 13955 15011
rect 13955 14977 13964 15011
rect 13912 14968 13964 14977
rect 16764 15036 16816 15088
rect 10140 14900 10192 14952
rect 10968 14943 11020 14952
rect 10968 14909 10977 14943
rect 10977 14909 11011 14943
rect 11011 14909 11020 14943
rect 10968 14900 11020 14909
rect 7380 14764 7432 14816
rect 9036 14807 9088 14816
rect 9036 14773 9045 14807
rect 9045 14773 9079 14807
rect 9079 14773 9088 14807
rect 9036 14764 9088 14773
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 10508 14764 10560 14816
rect 12072 14832 12124 14884
rect 12164 14832 12216 14884
rect 13176 14832 13228 14884
rect 13636 14875 13688 14884
rect 13636 14841 13645 14875
rect 13645 14841 13679 14875
rect 13679 14841 13688 14875
rect 13636 14832 13688 14841
rect 14188 14900 14240 14952
rect 14740 14943 14792 14952
rect 14740 14909 14749 14943
rect 14749 14909 14783 14943
rect 14783 14909 14792 14943
rect 14740 14900 14792 14909
rect 15844 14943 15896 14952
rect 15844 14909 15853 14943
rect 15853 14909 15887 14943
rect 15887 14909 15896 14943
rect 15844 14900 15896 14909
rect 16488 14968 16540 15020
rect 17868 15104 17920 15156
rect 17960 15104 18012 15156
rect 18420 15104 18472 15156
rect 18144 15036 18196 15088
rect 17132 14968 17184 15020
rect 19432 15104 19484 15156
rect 20444 15104 20496 15156
rect 18696 15036 18748 15088
rect 19892 15036 19944 15088
rect 16672 14900 16724 14952
rect 16948 14900 17000 14952
rect 17684 14900 17736 14952
rect 16212 14832 16264 14884
rect 11428 14764 11480 14816
rect 13820 14764 13872 14816
rect 13912 14764 13964 14816
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 14464 14764 14516 14773
rect 15476 14764 15528 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 16120 14764 16172 14816
rect 17316 14764 17368 14816
rect 17960 14900 18012 14952
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 21640 15036 21692 15088
rect 19984 14943 20036 14952
rect 19984 14909 19993 14943
rect 19993 14909 20027 14943
rect 20027 14909 20036 14943
rect 19984 14900 20036 14909
rect 18880 14875 18932 14884
rect 18880 14841 18889 14875
rect 18889 14841 18923 14875
rect 18923 14841 18932 14875
rect 18880 14832 18932 14841
rect 19248 14764 19300 14816
rect 19892 14764 19944 14816
rect 21824 14968 21876 15020
rect 23480 15104 23532 15156
rect 24400 15036 24452 15088
rect 27528 15104 27580 15156
rect 31300 15147 31352 15156
rect 31300 15113 31309 15147
rect 31309 15113 31343 15147
rect 31343 15113 31352 15147
rect 31300 15104 31352 15113
rect 33600 15147 33652 15156
rect 33600 15113 33609 15147
rect 33609 15113 33643 15147
rect 33643 15113 33652 15147
rect 33600 15104 33652 15113
rect 28724 14968 28776 15020
rect 31852 15011 31904 15020
rect 31852 14977 31861 15011
rect 31861 14977 31895 15011
rect 31895 14977 31904 15011
rect 31852 14968 31904 14977
rect 20904 14943 20956 14952
rect 20904 14909 20913 14943
rect 20913 14909 20947 14943
rect 20947 14909 20956 14943
rect 20904 14900 20956 14909
rect 20536 14875 20588 14884
rect 20536 14841 20545 14875
rect 20545 14841 20579 14875
rect 20579 14841 20588 14875
rect 20536 14832 20588 14841
rect 20720 14832 20772 14884
rect 20628 14764 20680 14816
rect 21548 14807 21600 14816
rect 21548 14773 21557 14807
rect 21557 14773 21591 14807
rect 21591 14773 21600 14807
rect 21548 14764 21600 14773
rect 22100 14832 22152 14884
rect 22468 14943 22520 14952
rect 22468 14909 22477 14943
rect 22477 14909 22511 14943
rect 22511 14909 22520 14943
rect 22468 14900 22520 14909
rect 26700 14943 26752 14952
rect 26700 14909 26709 14943
rect 26709 14909 26743 14943
rect 26743 14909 26752 14943
rect 26700 14900 26752 14909
rect 29828 14943 29880 14952
rect 29828 14909 29837 14943
rect 29837 14909 29871 14943
rect 29871 14909 29880 14943
rect 29828 14900 29880 14909
rect 30012 14943 30064 14952
rect 30012 14909 30021 14943
rect 30021 14909 30055 14943
rect 30055 14909 30064 14943
rect 30012 14900 30064 14909
rect 24676 14832 24728 14884
rect 27344 14875 27396 14884
rect 27344 14841 27353 14875
rect 27353 14841 27387 14875
rect 27387 14841 27396 14875
rect 27344 14832 27396 14841
rect 28080 14832 28132 14884
rect 28632 14832 28684 14884
rect 33876 14900 33928 14952
rect 32036 14832 32088 14884
rect 32128 14875 32180 14884
rect 32128 14841 32137 14875
rect 32137 14841 32171 14875
rect 32171 14841 32180 14875
rect 32128 14832 32180 14841
rect 22008 14807 22060 14816
rect 22008 14773 22017 14807
rect 22017 14773 22051 14807
rect 22051 14773 22060 14807
rect 22008 14764 22060 14773
rect 23388 14764 23440 14816
rect 29460 14764 29512 14816
rect 30656 14807 30708 14816
rect 30656 14773 30665 14807
rect 30665 14773 30699 14807
rect 30699 14773 30708 14807
rect 30656 14764 30708 14773
rect 31208 14764 31260 14816
rect 7210 14662 7262 14714
rect 7274 14662 7326 14714
rect 7338 14662 7390 14714
rect 7402 14662 7454 14714
rect 7466 14662 7518 14714
rect 15099 14662 15151 14714
rect 15163 14662 15215 14714
rect 15227 14662 15279 14714
rect 15291 14662 15343 14714
rect 15355 14662 15407 14714
rect 22988 14662 23040 14714
rect 23052 14662 23104 14714
rect 23116 14662 23168 14714
rect 23180 14662 23232 14714
rect 23244 14662 23296 14714
rect 30877 14662 30929 14714
rect 30941 14662 30993 14714
rect 31005 14662 31057 14714
rect 31069 14662 31121 14714
rect 31133 14662 31185 14714
rect 4160 14560 4212 14612
rect 4988 14492 5040 14544
rect 7104 14560 7156 14612
rect 7748 14603 7800 14612
rect 7748 14569 7757 14603
rect 7757 14569 7791 14603
rect 7791 14569 7800 14603
rect 7748 14560 7800 14569
rect 8852 14560 8904 14612
rect 10140 14560 10192 14612
rect 13636 14560 13688 14612
rect 14464 14560 14516 14612
rect 15200 14560 15252 14612
rect 15844 14560 15896 14612
rect 16396 14560 16448 14612
rect 17132 14560 17184 14612
rect 17316 14560 17368 14612
rect 17408 14560 17460 14612
rect 3056 14467 3108 14476
rect 3056 14433 3065 14467
rect 3065 14433 3099 14467
rect 3099 14433 3108 14467
rect 3056 14424 3108 14433
rect 5816 14467 5868 14476
rect 5816 14433 5825 14467
rect 5825 14433 5859 14467
rect 5859 14433 5868 14467
rect 5816 14424 5868 14433
rect 5448 14399 5500 14408
rect 5448 14365 5457 14399
rect 5457 14365 5491 14399
rect 5491 14365 5500 14399
rect 5448 14356 5500 14365
rect 4436 14288 4488 14340
rect 10048 14492 10100 14544
rect 6828 14424 6880 14476
rect 7472 14467 7524 14476
rect 7472 14433 7481 14467
rect 7481 14433 7515 14467
rect 7515 14433 7524 14467
rect 7472 14424 7524 14433
rect 8024 14424 8076 14476
rect 6368 14288 6420 14340
rect 6460 14288 6512 14340
rect 5632 14263 5684 14272
rect 5632 14229 5641 14263
rect 5641 14229 5675 14263
rect 5675 14229 5684 14263
rect 5632 14220 5684 14229
rect 5908 14220 5960 14272
rect 7472 14220 7524 14272
rect 8208 14220 8260 14272
rect 8300 14220 8352 14272
rect 9128 14356 9180 14408
rect 11428 14492 11480 14544
rect 13268 14467 13320 14476
rect 13268 14433 13277 14467
rect 13277 14433 13311 14467
rect 13311 14433 13320 14467
rect 13268 14424 13320 14433
rect 10232 14356 10284 14408
rect 10692 14399 10744 14408
rect 10692 14365 10701 14399
rect 10701 14365 10735 14399
rect 10735 14365 10744 14399
rect 10692 14356 10744 14365
rect 13912 14356 13964 14408
rect 16120 14492 16172 14544
rect 17960 14560 18012 14612
rect 19892 14560 19944 14612
rect 20352 14560 20404 14612
rect 22192 14560 22244 14612
rect 22468 14560 22520 14612
rect 24032 14603 24084 14612
rect 24032 14569 24041 14603
rect 24041 14569 24075 14603
rect 24075 14569 24084 14603
rect 24032 14560 24084 14569
rect 24676 14560 24728 14612
rect 26424 14560 26476 14612
rect 26700 14603 26752 14612
rect 26700 14569 26709 14603
rect 26709 14569 26743 14603
rect 26743 14569 26752 14603
rect 26700 14560 26752 14569
rect 27344 14560 27396 14612
rect 14924 14424 14976 14476
rect 15936 14424 15988 14476
rect 16488 14424 16540 14476
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 18696 14492 18748 14544
rect 18788 14492 18840 14544
rect 20076 14492 20128 14544
rect 17776 14467 17828 14476
rect 17776 14433 17785 14467
rect 17785 14433 17819 14467
rect 17819 14433 17828 14467
rect 17776 14424 17828 14433
rect 17868 14467 17920 14476
rect 17868 14433 17877 14467
rect 17877 14433 17911 14467
rect 17911 14433 17920 14467
rect 17868 14424 17920 14433
rect 20536 14467 20588 14476
rect 20536 14433 20545 14467
rect 20545 14433 20579 14467
rect 20579 14433 20588 14467
rect 20536 14424 20588 14433
rect 21180 14492 21232 14544
rect 26056 14492 26108 14544
rect 22468 14424 22520 14476
rect 22652 14424 22704 14476
rect 23756 14424 23808 14476
rect 24952 14424 25004 14476
rect 25780 14467 25832 14476
rect 25780 14433 25789 14467
rect 25789 14433 25823 14467
rect 25823 14433 25832 14467
rect 25780 14424 25832 14433
rect 25964 14467 26016 14476
rect 25964 14433 25973 14467
rect 25973 14433 26007 14467
rect 26007 14433 26016 14467
rect 25964 14424 26016 14433
rect 14740 14356 14792 14408
rect 16120 14356 16172 14408
rect 12808 14220 12860 14272
rect 14096 14220 14148 14272
rect 14924 14220 14976 14272
rect 15660 14263 15712 14272
rect 15660 14229 15669 14263
rect 15669 14229 15703 14263
rect 15703 14229 15712 14263
rect 15660 14220 15712 14229
rect 17224 14288 17276 14340
rect 18328 14288 18380 14340
rect 18052 14220 18104 14272
rect 18880 14288 18932 14340
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 21272 14356 21324 14408
rect 23204 14356 23256 14408
rect 23388 14356 23440 14408
rect 26424 14467 26476 14476
rect 26424 14433 26433 14467
rect 26433 14433 26467 14467
rect 26467 14433 26476 14467
rect 26424 14424 26476 14433
rect 27988 14492 28040 14544
rect 29000 14492 29052 14544
rect 29828 14603 29880 14612
rect 29828 14569 29837 14603
rect 29837 14569 29871 14603
rect 29871 14569 29880 14603
rect 29828 14560 29880 14569
rect 30012 14560 30064 14612
rect 30656 14560 30708 14612
rect 31208 14492 31260 14544
rect 26700 14424 26752 14476
rect 28632 14424 28684 14476
rect 29184 14467 29236 14476
rect 29184 14433 29193 14467
rect 29193 14433 29227 14467
rect 29227 14433 29236 14467
rect 29184 14424 29236 14433
rect 29460 14467 29512 14476
rect 29460 14433 29469 14467
rect 29469 14433 29503 14467
rect 29503 14433 29512 14467
rect 29460 14424 29512 14433
rect 29828 14424 29880 14476
rect 31852 14424 31904 14476
rect 32312 14424 32364 14476
rect 27068 14399 27120 14408
rect 27068 14365 27077 14399
rect 27077 14365 27111 14399
rect 27111 14365 27120 14399
rect 27068 14356 27120 14365
rect 32864 14399 32916 14408
rect 32864 14365 32873 14399
rect 32873 14365 32907 14399
rect 32907 14365 32916 14399
rect 32864 14356 32916 14365
rect 18696 14220 18748 14272
rect 20536 14220 20588 14272
rect 22284 14288 22336 14340
rect 24492 14288 24544 14340
rect 26884 14288 26936 14340
rect 28816 14288 28868 14340
rect 30012 14288 30064 14340
rect 33692 14356 33744 14408
rect 22192 14220 22244 14272
rect 22928 14220 22980 14272
rect 23388 14220 23440 14272
rect 26424 14220 26476 14272
rect 26792 14220 26844 14272
rect 28908 14220 28960 14272
rect 29000 14263 29052 14272
rect 29000 14229 29009 14263
rect 29009 14229 29043 14263
rect 29043 14229 29052 14263
rect 29000 14220 29052 14229
rect 32404 14263 32456 14272
rect 32404 14229 32413 14263
rect 32413 14229 32447 14263
rect 32447 14229 32456 14263
rect 32404 14220 32456 14229
rect 33508 14263 33560 14272
rect 33508 14229 33517 14263
rect 33517 14229 33551 14263
rect 33551 14229 33560 14263
rect 33508 14220 33560 14229
rect 6550 14118 6602 14170
rect 6614 14118 6666 14170
rect 6678 14118 6730 14170
rect 6742 14118 6794 14170
rect 6806 14118 6858 14170
rect 14439 14118 14491 14170
rect 14503 14118 14555 14170
rect 14567 14118 14619 14170
rect 14631 14118 14683 14170
rect 14695 14118 14747 14170
rect 22328 14118 22380 14170
rect 22392 14118 22444 14170
rect 22456 14118 22508 14170
rect 22520 14118 22572 14170
rect 22584 14118 22636 14170
rect 30217 14118 30269 14170
rect 30281 14118 30333 14170
rect 30345 14118 30397 14170
rect 30409 14118 30461 14170
rect 30473 14118 30525 14170
rect 4528 14016 4580 14068
rect 4712 14059 4764 14068
rect 4712 14025 4721 14059
rect 4721 14025 4755 14059
rect 4755 14025 4764 14059
rect 4712 14016 4764 14025
rect 4988 14059 5040 14068
rect 4988 14025 4997 14059
rect 4997 14025 5031 14059
rect 5031 14025 5040 14059
rect 4988 14016 5040 14025
rect 5632 14016 5684 14068
rect 5816 14016 5868 14068
rect 6184 14016 6236 14068
rect 1308 13880 1360 13932
rect 6920 13948 6972 14000
rect 8668 14059 8720 14068
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 9128 14059 9180 14068
rect 9128 14025 9137 14059
rect 9137 14025 9171 14059
rect 9171 14025 9180 14059
rect 9128 14016 9180 14025
rect 9772 14016 9824 14068
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 10692 14016 10744 14068
rect 12532 14016 12584 14068
rect 8944 13991 8996 14000
rect 8944 13957 8953 13991
rect 8953 13957 8987 13991
rect 8987 13957 8996 13991
rect 8944 13948 8996 13957
rect 12808 13948 12860 14000
rect 12900 13991 12952 14000
rect 12900 13957 12909 13991
rect 12909 13957 12943 13991
rect 12943 13957 12952 13991
rect 12900 13948 12952 13957
rect 13820 14016 13872 14068
rect 14280 14016 14332 14068
rect 13728 13948 13780 14000
rect 5172 13812 5224 13864
rect 6368 13812 6420 13864
rect 8208 13812 8260 13864
rect 8668 13812 8720 13864
rect 11704 13923 11756 13932
rect 11704 13889 11713 13923
rect 11713 13889 11747 13923
rect 11747 13889 11756 13923
rect 11704 13880 11756 13889
rect 12624 13880 12676 13932
rect 13176 13880 13228 13932
rect 14096 13880 14148 13932
rect 15568 14016 15620 14068
rect 16120 14016 16172 14068
rect 16028 13948 16080 14000
rect 16304 13948 16356 14000
rect 10048 13812 10100 13864
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 6460 13719 6512 13728
rect 6460 13685 6469 13719
rect 6469 13685 6503 13719
rect 6503 13685 6512 13719
rect 6460 13676 6512 13685
rect 8852 13744 8904 13796
rect 9956 13744 10008 13796
rect 10324 13812 10376 13864
rect 12348 13812 12400 13864
rect 13268 13812 13320 13864
rect 14280 13812 14332 13864
rect 14464 13855 14516 13864
rect 14464 13821 14473 13855
rect 14473 13821 14507 13855
rect 14507 13821 14516 13855
rect 14464 13812 14516 13821
rect 15568 13880 15620 13932
rect 10416 13744 10468 13796
rect 13084 13744 13136 13796
rect 15476 13812 15528 13864
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 16120 13880 16172 13932
rect 17040 14016 17092 14068
rect 17224 14016 17276 14068
rect 18420 14016 18472 14068
rect 18788 14059 18840 14068
rect 18788 14025 18797 14059
rect 18797 14025 18831 14059
rect 18831 14025 18840 14059
rect 18788 14016 18840 14025
rect 19064 14016 19116 14068
rect 20168 14016 20220 14068
rect 20352 14016 20404 14068
rect 20536 14016 20588 14068
rect 16764 13880 16816 13932
rect 16948 13880 17000 13932
rect 9864 13676 9916 13728
rect 13360 13719 13412 13728
rect 13360 13685 13369 13719
rect 13369 13685 13403 13719
rect 13403 13685 13412 13719
rect 13360 13676 13412 13685
rect 15016 13787 15068 13796
rect 15016 13753 15025 13787
rect 15025 13753 15059 13787
rect 15059 13753 15068 13787
rect 15016 13744 15068 13753
rect 15844 13744 15896 13796
rect 14464 13676 14516 13728
rect 16488 13676 16540 13728
rect 16856 13676 16908 13728
rect 17408 13948 17460 14000
rect 19248 13948 19300 14000
rect 21548 14016 21600 14068
rect 22100 13948 22152 14000
rect 22376 13948 22428 14000
rect 17592 13812 17644 13864
rect 18052 13744 18104 13796
rect 19340 13812 19392 13864
rect 20352 13812 20404 13864
rect 22284 13880 22336 13932
rect 22928 13923 22980 13932
rect 22928 13889 22937 13923
rect 22937 13889 22971 13923
rect 22971 13889 22980 13923
rect 22928 13880 22980 13889
rect 23388 13880 23440 13932
rect 23480 13923 23532 13932
rect 23480 13889 23489 13923
rect 23489 13889 23523 13923
rect 23523 13889 23532 13923
rect 23480 13880 23532 13889
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 18512 13744 18564 13796
rect 19064 13744 19116 13796
rect 20812 13744 20864 13796
rect 21640 13855 21692 13864
rect 21640 13821 21649 13855
rect 21649 13821 21683 13855
rect 21683 13821 21692 13855
rect 21640 13812 21692 13821
rect 17132 13719 17184 13728
rect 17132 13685 17141 13719
rect 17141 13685 17175 13719
rect 17175 13685 17184 13719
rect 17132 13676 17184 13685
rect 19156 13676 19208 13728
rect 20076 13719 20128 13728
rect 20076 13685 20085 13719
rect 20085 13685 20119 13719
rect 20119 13685 20128 13719
rect 20076 13676 20128 13685
rect 20444 13676 20496 13728
rect 22008 13812 22060 13864
rect 22008 13676 22060 13728
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 24216 13880 24268 13932
rect 24124 13855 24176 13864
rect 24124 13821 24133 13855
rect 24133 13821 24167 13855
rect 24167 13821 24176 13855
rect 24124 13812 24176 13821
rect 24492 14016 24544 14068
rect 25780 14016 25832 14068
rect 25964 14016 26016 14068
rect 26884 14016 26936 14068
rect 27068 14059 27120 14068
rect 27068 14025 27077 14059
rect 27077 14025 27111 14059
rect 27111 14025 27120 14059
rect 27068 14016 27120 14025
rect 25688 13991 25740 14000
rect 25688 13957 25697 13991
rect 25697 13957 25731 13991
rect 25731 13957 25740 13991
rect 25688 13948 25740 13957
rect 26608 13948 26660 14000
rect 27620 14016 27672 14068
rect 28908 14016 28960 14068
rect 29092 14016 29144 14068
rect 27528 13880 27580 13932
rect 24032 13676 24084 13728
rect 24216 13719 24268 13728
rect 24216 13685 24225 13719
rect 24225 13685 24259 13719
rect 24259 13685 24268 13719
rect 24216 13676 24268 13685
rect 26424 13855 26476 13864
rect 26424 13821 26433 13855
rect 26433 13821 26467 13855
rect 26467 13821 26476 13855
rect 26424 13812 26476 13821
rect 26608 13855 26660 13864
rect 26608 13821 26617 13855
rect 26617 13821 26651 13855
rect 26651 13821 26660 13855
rect 26608 13812 26660 13821
rect 26700 13855 26752 13864
rect 26700 13821 26709 13855
rect 26709 13821 26743 13855
rect 26743 13821 26752 13855
rect 26700 13812 26752 13821
rect 26792 13855 26844 13864
rect 26792 13821 26801 13855
rect 26801 13821 26835 13855
rect 26835 13821 26844 13855
rect 26792 13812 26844 13821
rect 27068 13855 27120 13864
rect 27068 13821 27077 13855
rect 27077 13821 27111 13855
rect 27111 13821 27120 13855
rect 27068 13812 27120 13821
rect 29000 13812 29052 13864
rect 29092 13855 29144 13864
rect 29092 13821 29101 13855
rect 29101 13821 29135 13855
rect 29135 13821 29144 13855
rect 29092 13812 29144 13821
rect 30012 13923 30064 13932
rect 30012 13889 30021 13923
rect 30021 13889 30055 13923
rect 30055 13889 30064 13923
rect 30012 13880 30064 13889
rect 29736 13812 29788 13864
rect 29828 13855 29880 13864
rect 29828 13821 29837 13855
rect 29837 13821 29871 13855
rect 29871 13821 29880 13855
rect 29828 13812 29880 13821
rect 29920 13812 29972 13864
rect 31208 13855 31260 13864
rect 31208 13821 31217 13855
rect 31217 13821 31251 13855
rect 31251 13821 31260 13855
rect 31208 13812 31260 13821
rect 32128 14016 32180 14068
rect 32404 14016 32456 14068
rect 32864 14016 32916 14068
rect 33600 13880 33652 13932
rect 31484 13855 31536 13864
rect 31484 13821 31493 13855
rect 31493 13821 31527 13855
rect 31527 13821 31536 13855
rect 31484 13812 31536 13821
rect 27436 13787 27488 13796
rect 27436 13753 27445 13787
rect 27445 13753 27479 13787
rect 27479 13753 27488 13787
rect 27436 13744 27488 13753
rect 30196 13787 30248 13796
rect 30196 13753 30205 13787
rect 30205 13753 30239 13787
rect 30239 13753 30248 13787
rect 30196 13744 30248 13753
rect 30564 13787 30616 13796
rect 30564 13753 30573 13787
rect 30573 13753 30607 13787
rect 30607 13753 30616 13787
rect 30564 13744 30616 13753
rect 27712 13676 27764 13728
rect 28908 13719 28960 13728
rect 28908 13685 28917 13719
rect 28917 13685 28951 13719
rect 28951 13685 28960 13719
rect 28908 13676 28960 13685
rect 29092 13676 29144 13728
rect 30472 13676 30524 13728
rect 31300 13676 31352 13728
rect 7210 13574 7262 13626
rect 7274 13574 7326 13626
rect 7338 13574 7390 13626
rect 7402 13574 7454 13626
rect 7466 13574 7518 13626
rect 15099 13574 15151 13626
rect 15163 13574 15215 13626
rect 15227 13574 15279 13626
rect 15291 13574 15343 13626
rect 15355 13574 15407 13626
rect 22988 13574 23040 13626
rect 23052 13574 23104 13626
rect 23116 13574 23168 13626
rect 23180 13574 23232 13626
rect 23244 13574 23296 13626
rect 30877 13574 30929 13626
rect 30941 13574 30993 13626
rect 31005 13574 31057 13626
rect 31069 13574 31121 13626
rect 31133 13574 31185 13626
rect 5448 13472 5500 13524
rect 6276 13472 6328 13524
rect 7932 13472 7984 13524
rect 9128 13472 9180 13524
rect 9864 13472 9916 13524
rect 10416 13515 10468 13524
rect 10416 13481 10425 13515
rect 10425 13481 10459 13515
rect 10459 13481 10468 13515
rect 10416 13472 10468 13481
rect 5540 13404 5592 13456
rect 6460 13404 6512 13456
rect 8484 13404 8536 13456
rect 10600 13404 10652 13456
rect 11704 13472 11756 13524
rect 12900 13472 12952 13524
rect 14464 13515 14516 13524
rect 14464 13481 14473 13515
rect 14473 13481 14507 13515
rect 14507 13481 14516 13515
rect 14464 13472 14516 13481
rect 15568 13472 15620 13524
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 12992 13404 13044 13456
rect 13084 13404 13136 13456
rect 13820 13404 13872 13456
rect 14556 13404 14608 13456
rect 4068 13336 4120 13388
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 6552 13336 6604 13388
rect 8208 13379 8260 13388
rect 8208 13345 8217 13379
rect 8217 13345 8251 13379
rect 8251 13345 8260 13379
rect 8208 13336 8260 13345
rect 10416 13336 10468 13388
rect 11612 13336 11664 13388
rect 13176 13379 13228 13388
rect 13176 13345 13185 13379
rect 13185 13345 13219 13379
rect 13219 13345 13228 13379
rect 13176 13336 13228 13345
rect 1308 13268 1360 13320
rect 8024 13268 8076 13320
rect 6276 13132 6328 13184
rect 6368 13132 6420 13184
rect 8116 13132 8168 13184
rect 12072 13268 12124 13320
rect 13360 13268 13412 13320
rect 14740 13336 14792 13388
rect 14188 13311 14240 13320
rect 14188 13277 14197 13311
rect 14197 13277 14231 13311
rect 14231 13277 14240 13311
rect 14188 13268 14240 13277
rect 15568 13379 15620 13388
rect 15568 13345 15577 13379
rect 15577 13345 15611 13379
rect 15611 13345 15620 13379
rect 15568 13336 15620 13345
rect 16396 13404 16448 13456
rect 17500 13472 17552 13524
rect 17684 13472 17736 13524
rect 20720 13472 20772 13524
rect 20812 13472 20864 13524
rect 21180 13472 21232 13524
rect 18052 13404 18104 13456
rect 16488 13379 16540 13388
rect 16488 13345 16497 13379
rect 16497 13345 16531 13379
rect 16531 13345 16540 13379
rect 16488 13336 16540 13345
rect 16764 13336 16816 13388
rect 17408 13336 17460 13388
rect 17776 13379 17828 13388
rect 17776 13345 17785 13379
rect 17785 13345 17819 13379
rect 17819 13345 17828 13379
rect 17776 13336 17828 13345
rect 14648 13200 14700 13252
rect 15016 13200 15068 13252
rect 16856 13268 16908 13320
rect 9036 13132 9088 13184
rect 12440 13132 12492 13184
rect 12900 13132 12952 13184
rect 12992 13175 13044 13184
rect 12992 13141 13001 13175
rect 13001 13141 13035 13175
rect 13035 13141 13044 13175
rect 12992 13132 13044 13141
rect 15476 13132 15528 13184
rect 15936 13175 15988 13184
rect 15936 13141 15945 13175
rect 15945 13141 15979 13175
rect 15979 13141 15988 13175
rect 15936 13132 15988 13141
rect 16580 13175 16632 13184
rect 16580 13141 16589 13175
rect 16589 13141 16623 13175
rect 16623 13141 16632 13175
rect 16580 13132 16632 13141
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 17316 13268 17368 13320
rect 17684 13268 17736 13320
rect 18604 13336 18656 13388
rect 18788 13336 18840 13388
rect 19156 13379 19208 13388
rect 19156 13345 19166 13379
rect 19166 13345 19200 13379
rect 19200 13345 19208 13379
rect 19156 13336 19208 13345
rect 17868 13200 17920 13252
rect 20628 13336 20680 13388
rect 20904 13336 20956 13388
rect 23480 13472 23532 13524
rect 24216 13472 24268 13524
rect 25688 13472 25740 13524
rect 26516 13472 26568 13524
rect 27436 13515 27488 13524
rect 27436 13481 27445 13515
rect 27445 13481 27479 13515
rect 27479 13481 27488 13515
rect 27436 13472 27488 13481
rect 26148 13447 26200 13456
rect 26148 13413 26157 13447
rect 26157 13413 26191 13447
rect 26191 13413 26200 13447
rect 26148 13404 26200 13413
rect 22008 13311 22060 13320
rect 22008 13277 22017 13311
rect 22017 13277 22051 13311
rect 22051 13277 22060 13311
rect 22008 13268 22060 13277
rect 17316 13132 17368 13184
rect 19616 13200 19668 13252
rect 22652 13336 22704 13388
rect 23848 13268 23900 13320
rect 24032 13311 24084 13320
rect 24032 13277 24041 13311
rect 24041 13277 24075 13311
rect 24075 13277 24084 13311
rect 24032 13268 24084 13277
rect 24492 13311 24544 13320
rect 24492 13277 24501 13311
rect 24501 13277 24535 13311
rect 24535 13277 24544 13311
rect 24492 13268 24544 13277
rect 24676 13379 24728 13388
rect 24676 13345 24685 13379
rect 24685 13345 24719 13379
rect 24719 13345 24728 13379
rect 24676 13336 24728 13345
rect 26056 13379 26108 13388
rect 26056 13345 26065 13379
rect 26065 13345 26099 13379
rect 26099 13345 26108 13379
rect 26056 13336 26108 13345
rect 26240 13379 26292 13388
rect 26240 13345 26249 13379
rect 26249 13345 26283 13379
rect 26283 13345 26292 13379
rect 26240 13336 26292 13345
rect 26332 13379 26384 13388
rect 26332 13345 26367 13379
rect 26367 13345 26384 13379
rect 26332 13336 26384 13345
rect 27068 13379 27120 13388
rect 27068 13345 27077 13379
rect 27077 13345 27111 13379
rect 27111 13345 27120 13379
rect 27068 13336 27120 13345
rect 27896 13336 27948 13388
rect 25688 13311 25740 13320
rect 25688 13277 25697 13311
rect 25697 13277 25731 13311
rect 25731 13277 25740 13311
rect 25688 13268 25740 13277
rect 26608 13268 26660 13320
rect 19248 13175 19300 13184
rect 19248 13141 19257 13175
rect 19257 13141 19291 13175
rect 19291 13141 19300 13175
rect 19248 13132 19300 13141
rect 19340 13132 19392 13184
rect 21732 13132 21784 13184
rect 22100 13132 22152 13184
rect 22284 13132 22336 13184
rect 22376 13175 22428 13184
rect 22376 13141 22385 13175
rect 22385 13141 22419 13175
rect 22419 13141 22428 13175
rect 22376 13132 22428 13141
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 24124 13132 24176 13184
rect 25044 13175 25096 13184
rect 25044 13141 25053 13175
rect 25053 13141 25087 13175
rect 25087 13141 25096 13175
rect 25044 13132 25096 13141
rect 26976 13200 27028 13252
rect 28356 13379 28408 13388
rect 28356 13345 28365 13379
rect 28365 13345 28399 13379
rect 28399 13345 28408 13379
rect 28356 13336 28408 13345
rect 28816 13472 28868 13524
rect 29184 13472 29236 13524
rect 29460 13515 29512 13524
rect 29460 13481 29469 13515
rect 29469 13481 29503 13515
rect 29503 13481 29512 13515
rect 29460 13472 29512 13481
rect 30288 13472 30340 13524
rect 30380 13472 30432 13524
rect 28908 13336 28960 13388
rect 29092 13336 29144 13388
rect 30012 13336 30064 13388
rect 30196 13379 30248 13388
rect 30196 13345 30205 13379
rect 30205 13345 30239 13379
rect 30239 13345 30248 13379
rect 30196 13336 30248 13345
rect 30472 13447 30524 13456
rect 30472 13413 30481 13447
rect 30481 13413 30515 13447
rect 30515 13413 30524 13447
rect 31484 13472 31536 13524
rect 30472 13404 30524 13413
rect 32312 13404 32364 13456
rect 33048 13472 33100 13524
rect 35164 13472 35216 13524
rect 29920 13268 29972 13320
rect 32588 13379 32640 13388
rect 32588 13345 32597 13379
rect 32597 13345 32631 13379
rect 32631 13345 32640 13379
rect 32588 13336 32640 13345
rect 32312 13311 32364 13320
rect 32312 13277 32321 13311
rect 32321 13277 32355 13311
rect 32355 13277 32364 13311
rect 32312 13268 32364 13277
rect 29276 13200 29328 13252
rect 29920 13132 29972 13184
rect 6550 13030 6602 13082
rect 6614 13030 6666 13082
rect 6678 13030 6730 13082
rect 6742 13030 6794 13082
rect 6806 13030 6858 13082
rect 14439 13030 14491 13082
rect 14503 13030 14555 13082
rect 14567 13030 14619 13082
rect 14631 13030 14683 13082
rect 14695 13030 14747 13082
rect 22328 13030 22380 13082
rect 22392 13030 22444 13082
rect 22456 13030 22508 13082
rect 22520 13030 22572 13082
rect 22584 13030 22636 13082
rect 30217 13030 30269 13082
rect 30281 13030 30333 13082
rect 30345 13030 30397 13082
rect 30409 13030 30461 13082
rect 30473 13030 30525 13082
rect 3976 12928 4028 12980
rect 4344 12928 4396 12980
rect 6460 12928 6512 12980
rect 8576 12928 8628 12980
rect 8944 12928 8996 12980
rect 4344 12792 4396 12844
rect 3884 12767 3936 12776
rect 3884 12733 3893 12767
rect 3893 12733 3927 12767
rect 3927 12733 3936 12767
rect 3884 12724 3936 12733
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 5724 12767 5776 12776
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 5724 12724 5776 12733
rect 5908 12724 5960 12776
rect 5540 12656 5592 12708
rect 4528 12631 4580 12640
rect 4528 12597 4537 12631
rect 4537 12597 4571 12631
rect 4571 12597 4580 12631
rect 4528 12588 4580 12597
rect 5448 12588 5500 12640
rect 6184 12588 6236 12640
rect 6460 12631 6512 12640
rect 6460 12597 6469 12631
rect 6469 12597 6503 12631
rect 6503 12597 6512 12631
rect 6460 12588 6512 12597
rect 7840 12767 7892 12776
rect 7840 12733 7849 12767
rect 7849 12733 7883 12767
rect 7883 12733 7892 12767
rect 7840 12724 7892 12733
rect 8116 12724 8168 12776
rect 8576 12724 8628 12776
rect 12440 12928 12492 12980
rect 12716 12928 12768 12980
rect 12992 12928 13044 12980
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 16304 12928 16356 12980
rect 16764 12971 16816 12980
rect 16764 12937 16773 12971
rect 16773 12937 16807 12971
rect 16807 12937 16816 12971
rect 16764 12928 16816 12937
rect 16856 12971 16908 12980
rect 16856 12937 16865 12971
rect 16865 12937 16899 12971
rect 16899 12937 16908 12971
rect 16856 12928 16908 12937
rect 17316 12928 17368 12980
rect 18052 12928 18104 12980
rect 18144 12928 18196 12980
rect 18604 12928 18656 12980
rect 19248 12971 19300 12980
rect 19248 12937 19257 12971
rect 19257 12937 19291 12971
rect 19291 12937 19300 12971
rect 19248 12928 19300 12937
rect 20076 12928 20128 12980
rect 20168 12928 20220 12980
rect 22008 12928 22060 12980
rect 22100 12928 22152 12980
rect 22192 12928 22244 12980
rect 22836 12971 22888 12980
rect 22836 12937 22845 12971
rect 22845 12937 22879 12971
rect 22879 12937 22888 12971
rect 22836 12928 22888 12937
rect 23296 12928 23348 12980
rect 25688 12928 25740 12980
rect 15016 12860 15068 12912
rect 16028 12860 16080 12912
rect 11704 12792 11756 12844
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 8300 12656 8352 12708
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 8576 12631 8628 12640
rect 8576 12597 8585 12631
rect 8585 12597 8619 12631
rect 8619 12597 8628 12631
rect 8576 12588 8628 12597
rect 9036 12656 9088 12708
rect 12348 12792 12400 12844
rect 15200 12835 15252 12844
rect 15200 12801 15209 12835
rect 15209 12801 15243 12835
rect 15243 12801 15252 12835
rect 15200 12792 15252 12801
rect 15476 12835 15528 12844
rect 15476 12801 15485 12835
rect 15485 12801 15519 12835
rect 15519 12801 15528 12835
rect 15476 12792 15528 12801
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 15568 12724 15620 12776
rect 16028 12767 16080 12776
rect 16028 12733 16037 12767
rect 16037 12733 16071 12767
rect 16071 12733 16080 12767
rect 16028 12724 16080 12733
rect 16304 12724 16356 12776
rect 16580 12767 16632 12776
rect 16580 12733 16589 12767
rect 16589 12733 16623 12767
rect 16623 12733 16632 12767
rect 16580 12724 16632 12733
rect 16764 12767 16816 12776
rect 16764 12733 16773 12767
rect 16773 12733 16807 12767
rect 16807 12733 16816 12767
rect 16764 12724 16816 12733
rect 16948 12724 17000 12776
rect 17684 12860 17736 12912
rect 17592 12767 17644 12776
rect 17592 12733 17601 12767
rect 17601 12733 17635 12767
rect 17635 12733 17644 12767
rect 17592 12724 17644 12733
rect 18972 12767 19024 12776
rect 18972 12733 18981 12767
rect 18981 12733 19015 12767
rect 19015 12733 19024 12767
rect 18972 12724 19024 12733
rect 21640 12860 21692 12912
rect 19524 12724 19576 12776
rect 24676 12860 24728 12912
rect 27712 12971 27764 12980
rect 27712 12937 27721 12971
rect 27721 12937 27755 12971
rect 27755 12937 27764 12971
rect 27712 12928 27764 12937
rect 28816 12928 28868 12980
rect 32312 12928 32364 12980
rect 23756 12792 23808 12844
rect 12164 12656 12216 12708
rect 10600 12588 10652 12640
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 11428 12588 11480 12640
rect 11612 12588 11664 12640
rect 12900 12656 12952 12708
rect 14188 12656 14240 12708
rect 15936 12656 15988 12708
rect 17776 12656 17828 12708
rect 13176 12588 13228 12640
rect 14924 12588 14976 12640
rect 17040 12588 17092 12640
rect 17408 12588 17460 12640
rect 18512 12588 18564 12640
rect 22744 12724 22796 12776
rect 22928 12724 22980 12776
rect 25044 12792 25096 12844
rect 26240 12792 26292 12844
rect 28356 12792 28408 12844
rect 28816 12792 28868 12844
rect 31300 12835 31352 12844
rect 31300 12801 31309 12835
rect 31309 12801 31343 12835
rect 31343 12801 31352 12835
rect 31300 12792 31352 12801
rect 26148 12724 26200 12776
rect 27068 12724 27120 12776
rect 27988 12724 28040 12776
rect 29184 12767 29236 12776
rect 29184 12733 29193 12767
rect 29193 12733 29227 12767
rect 29227 12733 29236 12767
rect 29184 12724 29236 12733
rect 29552 12767 29604 12776
rect 29552 12733 29561 12767
rect 29561 12733 29595 12767
rect 29595 12733 29604 12767
rect 29552 12724 29604 12733
rect 30380 12767 30432 12776
rect 30380 12733 30389 12767
rect 30389 12733 30423 12767
rect 30423 12733 30432 12767
rect 30380 12724 30432 12733
rect 34428 12724 34480 12776
rect 19984 12699 20036 12708
rect 19984 12665 19993 12699
rect 19993 12665 20027 12699
rect 20027 12665 20036 12699
rect 19984 12656 20036 12665
rect 20444 12656 20496 12708
rect 21456 12656 21508 12708
rect 23756 12656 23808 12708
rect 23940 12656 23992 12708
rect 26516 12656 26568 12708
rect 27528 12656 27580 12708
rect 28080 12699 28132 12708
rect 28080 12665 28089 12699
rect 28089 12665 28123 12699
rect 28123 12665 28132 12699
rect 28080 12656 28132 12665
rect 19892 12588 19944 12640
rect 24308 12588 24360 12640
rect 26884 12631 26936 12640
rect 26884 12597 26893 12631
rect 26893 12597 26927 12631
rect 26927 12597 26936 12631
rect 26884 12588 26936 12597
rect 30012 12588 30064 12640
rect 31760 12588 31812 12640
rect 7210 12486 7262 12538
rect 7274 12486 7326 12538
rect 7338 12486 7390 12538
rect 7402 12486 7454 12538
rect 7466 12486 7518 12538
rect 15099 12486 15151 12538
rect 15163 12486 15215 12538
rect 15227 12486 15279 12538
rect 15291 12486 15343 12538
rect 15355 12486 15407 12538
rect 22988 12486 23040 12538
rect 23052 12486 23104 12538
rect 23116 12486 23168 12538
rect 23180 12486 23232 12538
rect 23244 12486 23296 12538
rect 30877 12486 30929 12538
rect 30941 12486 30993 12538
rect 31005 12486 31057 12538
rect 31069 12486 31121 12538
rect 31133 12486 31185 12538
rect 3884 12384 3936 12436
rect 5540 12384 5592 12436
rect 5816 12316 5868 12368
rect 6184 12384 6236 12436
rect 7840 12384 7892 12436
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 12164 12384 12216 12436
rect 12624 12384 12676 12436
rect 12900 12427 12952 12436
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 13176 12427 13228 12436
rect 13176 12393 13185 12427
rect 13185 12393 13219 12427
rect 13219 12393 13228 12427
rect 13176 12384 13228 12393
rect 13452 12384 13504 12436
rect 13820 12384 13872 12436
rect 14280 12384 14332 12436
rect 6552 12359 6604 12368
rect 6552 12325 6561 12359
rect 6561 12325 6595 12359
rect 6595 12325 6604 12359
rect 6552 12316 6604 12325
rect 8576 12316 8628 12368
rect 10784 12316 10836 12368
rect 3976 12180 4028 12232
rect 4068 12223 4120 12232
rect 4068 12189 4077 12223
rect 4077 12189 4111 12223
rect 4111 12189 4120 12223
rect 4068 12180 4120 12189
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 6368 12248 6420 12300
rect 5172 12180 5224 12232
rect 5264 12180 5316 12232
rect 8208 12291 8260 12300
rect 6828 12180 6880 12232
rect 8208 12257 8217 12291
rect 8217 12257 8251 12291
rect 8251 12257 8260 12291
rect 8208 12248 8260 12257
rect 9772 12248 9824 12300
rect 10232 12291 10284 12300
rect 10232 12257 10241 12291
rect 10241 12257 10275 12291
rect 10275 12257 10284 12291
rect 10232 12248 10284 12257
rect 11612 12248 11664 12300
rect 7012 12180 7064 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 7656 12180 7708 12232
rect 10600 12180 10652 12232
rect 13268 12248 13320 12300
rect 14648 12291 14700 12300
rect 14648 12257 14657 12291
rect 14657 12257 14691 12291
rect 14691 12257 14700 12291
rect 14648 12248 14700 12257
rect 16120 12316 16172 12368
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 15016 12248 15068 12300
rect 14832 12112 14884 12164
rect 16028 12248 16080 12300
rect 16580 12316 16632 12368
rect 16856 12359 16908 12368
rect 16856 12325 16865 12359
rect 16865 12325 16899 12359
rect 16899 12325 16908 12359
rect 16856 12316 16908 12325
rect 15476 12223 15528 12232
rect 15476 12189 15485 12223
rect 15485 12189 15519 12223
rect 15519 12189 15528 12223
rect 15476 12180 15528 12189
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 15844 12180 15896 12232
rect 15568 12112 15620 12164
rect 17132 12316 17184 12368
rect 17868 12316 17920 12368
rect 18972 12384 19024 12436
rect 19156 12384 19208 12436
rect 19524 12384 19576 12436
rect 19892 12384 19944 12436
rect 18604 12316 18656 12368
rect 19524 12248 19576 12300
rect 20720 12427 20772 12436
rect 20720 12393 20729 12427
rect 20729 12393 20763 12427
rect 20763 12393 20772 12427
rect 20720 12384 20772 12393
rect 20996 12384 21048 12436
rect 20904 12291 20956 12300
rect 20904 12257 20913 12291
rect 20913 12257 20947 12291
rect 20947 12257 20956 12291
rect 20904 12248 20956 12257
rect 20996 12248 21048 12300
rect 23940 12427 23992 12436
rect 23940 12393 23949 12427
rect 23949 12393 23983 12427
rect 23983 12393 23992 12427
rect 23940 12384 23992 12393
rect 23756 12316 23808 12368
rect 18052 12180 18104 12232
rect 17224 12112 17276 12164
rect 18880 12180 18932 12232
rect 20812 12180 20864 12232
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21272 12112 21324 12164
rect 3424 12087 3476 12096
rect 3424 12053 3433 12087
rect 3433 12053 3467 12087
rect 3467 12053 3476 12087
rect 3424 12044 3476 12053
rect 4436 12087 4488 12096
rect 4436 12053 4445 12087
rect 4445 12053 4479 12087
rect 4479 12053 4488 12087
rect 4436 12044 4488 12053
rect 5908 12044 5960 12096
rect 6552 12044 6604 12096
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 8392 12044 8444 12096
rect 10140 12087 10192 12096
rect 10140 12053 10149 12087
rect 10149 12053 10183 12087
rect 10183 12053 10192 12087
rect 10140 12044 10192 12053
rect 12716 12087 12768 12096
rect 12716 12053 12725 12087
rect 12725 12053 12759 12087
rect 12759 12053 12768 12087
rect 12716 12044 12768 12053
rect 12900 12044 12952 12096
rect 14924 12044 14976 12096
rect 15752 12044 15804 12096
rect 16304 12044 16356 12096
rect 17868 12044 17920 12096
rect 18788 12044 18840 12096
rect 19432 12087 19484 12096
rect 19432 12053 19441 12087
rect 19441 12053 19475 12087
rect 19475 12053 19484 12087
rect 19432 12044 19484 12053
rect 19984 12044 20036 12096
rect 21548 12044 21600 12096
rect 23572 12248 23624 12300
rect 22008 12180 22060 12232
rect 24124 12248 24176 12300
rect 25228 12384 25280 12436
rect 26424 12384 26476 12436
rect 26700 12384 26752 12436
rect 27896 12384 27948 12436
rect 28908 12384 28960 12436
rect 29276 12384 29328 12436
rect 29552 12384 29604 12436
rect 30104 12384 30156 12436
rect 33508 12427 33560 12436
rect 33508 12393 33517 12427
rect 33517 12393 33551 12427
rect 33551 12393 33560 12427
rect 33508 12384 33560 12393
rect 24584 12291 24636 12300
rect 24584 12257 24593 12291
rect 24593 12257 24627 12291
rect 24627 12257 24636 12291
rect 24584 12248 24636 12257
rect 24952 12180 25004 12232
rect 25320 12223 25372 12232
rect 25320 12189 25329 12223
rect 25329 12189 25363 12223
rect 25363 12189 25372 12223
rect 25320 12180 25372 12189
rect 25504 12180 25556 12232
rect 26424 12248 26476 12300
rect 26240 12180 26292 12232
rect 26976 12291 27028 12300
rect 26976 12257 26985 12291
rect 26985 12257 27019 12291
rect 27019 12257 27028 12291
rect 26976 12248 27028 12257
rect 29000 12291 29052 12300
rect 29000 12257 29009 12291
rect 29009 12257 29043 12291
rect 29043 12257 29052 12291
rect 29000 12248 29052 12257
rect 29736 12359 29788 12368
rect 29736 12325 29745 12359
rect 29745 12325 29779 12359
rect 29779 12325 29788 12359
rect 29736 12316 29788 12325
rect 30012 12316 30064 12368
rect 31300 12316 31352 12368
rect 31760 12359 31812 12368
rect 31760 12325 31769 12359
rect 31769 12325 31803 12359
rect 31803 12325 31812 12359
rect 31760 12316 31812 12325
rect 29276 12291 29328 12300
rect 29276 12257 29285 12291
rect 29285 12257 29319 12291
rect 29319 12257 29328 12291
rect 29276 12248 29328 12257
rect 27068 12180 27120 12232
rect 22744 12044 22796 12096
rect 23388 12044 23440 12096
rect 30380 12180 30432 12232
rect 32588 12248 32640 12300
rect 31208 12180 31260 12232
rect 32680 12223 32732 12232
rect 32680 12189 32689 12223
rect 32689 12189 32723 12223
rect 32723 12189 32732 12223
rect 32680 12180 32732 12189
rect 29920 12112 29972 12164
rect 27068 12087 27120 12096
rect 27068 12053 27077 12087
rect 27077 12053 27111 12087
rect 27111 12053 27120 12087
rect 27068 12044 27120 12053
rect 32128 12087 32180 12096
rect 32128 12053 32137 12087
rect 32137 12053 32171 12087
rect 32171 12053 32180 12087
rect 32128 12044 32180 12053
rect 33048 12087 33100 12096
rect 33048 12053 33057 12087
rect 33057 12053 33091 12087
rect 33091 12053 33100 12087
rect 33048 12044 33100 12053
rect 6550 11942 6602 11994
rect 6614 11942 6666 11994
rect 6678 11942 6730 11994
rect 6742 11942 6794 11994
rect 6806 11942 6858 11994
rect 14439 11942 14491 11994
rect 14503 11942 14555 11994
rect 14567 11942 14619 11994
rect 14631 11942 14683 11994
rect 14695 11942 14747 11994
rect 22328 11942 22380 11994
rect 22392 11942 22444 11994
rect 22456 11942 22508 11994
rect 22520 11942 22572 11994
rect 22584 11942 22636 11994
rect 30217 11942 30269 11994
rect 30281 11942 30333 11994
rect 30345 11942 30397 11994
rect 30409 11942 30461 11994
rect 30473 11942 30525 11994
rect 4068 11840 4120 11892
rect 5172 11840 5224 11892
rect 5264 11883 5316 11892
rect 5264 11849 5273 11883
rect 5273 11849 5307 11883
rect 5307 11849 5316 11883
rect 5264 11840 5316 11849
rect 5724 11840 5776 11892
rect 5816 11840 5868 11892
rect 7472 11840 7524 11892
rect 8392 11840 8444 11892
rect 8944 11840 8996 11892
rect 9772 11840 9824 11892
rect 12532 11840 12584 11892
rect 12716 11840 12768 11892
rect 13084 11840 13136 11892
rect 13360 11840 13412 11892
rect 14832 11840 14884 11892
rect 15200 11840 15252 11892
rect 15568 11840 15620 11892
rect 4528 11747 4580 11756
rect 4528 11713 4537 11747
rect 4537 11713 4571 11747
rect 4571 11713 4580 11747
rect 4528 11704 4580 11713
rect 5540 11704 5592 11756
rect 3424 11636 3476 11688
rect 6184 11636 6236 11688
rect 7012 11772 7064 11824
rect 10140 11772 10192 11824
rect 7656 11704 7708 11756
rect 10048 11636 10100 11688
rect 11152 11636 11204 11688
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 11612 11636 11664 11688
rect 12900 11636 12952 11688
rect 5448 11568 5500 11620
rect 6920 11568 6972 11620
rect 8116 11568 8168 11620
rect 8484 11568 8536 11620
rect 4620 11500 4672 11552
rect 5816 11543 5868 11552
rect 5816 11509 5825 11543
rect 5825 11509 5859 11543
rect 5859 11509 5868 11543
rect 5816 11500 5868 11509
rect 12164 11568 12216 11620
rect 10784 11500 10836 11552
rect 10968 11500 11020 11552
rect 12900 11500 12952 11552
rect 15844 11772 15896 11824
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 14188 11704 14240 11756
rect 15016 11704 15068 11756
rect 15200 11747 15252 11756
rect 15200 11713 15209 11747
rect 15209 11713 15243 11747
rect 15243 11713 15252 11747
rect 15200 11704 15252 11713
rect 15660 11704 15712 11756
rect 16028 11747 16080 11756
rect 16028 11713 16037 11747
rect 16037 11713 16071 11747
rect 16071 11713 16080 11747
rect 16028 11704 16080 11713
rect 16304 11772 16356 11824
rect 17408 11772 17460 11824
rect 18512 11883 18564 11892
rect 18512 11849 18521 11883
rect 18521 11849 18555 11883
rect 18555 11849 18564 11883
rect 18512 11840 18564 11849
rect 18696 11883 18748 11892
rect 18696 11849 18705 11883
rect 18705 11849 18739 11883
rect 18739 11849 18748 11883
rect 18696 11840 18748 11849
rect 19248 11840 19300 11892
rect 19340 11840 19392 11892
rect 20720 11840 20772 11892
rect 21916 11840 21968 11892
rect 22652 11883 22704 11892
rect 22652 11849 22661 11883
rect 22661 11849 22695 11883
rect 22695 11849 22704 11883
rect 22652 11840 22704 11849
rect 27068 11883 27120 11892
rect 27068 11849 27098 11883
rect 27098 11849 27120 11883
rect 27068 11840 27120 11849
rect 29276 11840 29328 11892
rect 31300 11883 31352 11892
rect 31300 11849 31309 11883
rect 31309 11849 31343 11883
rect 31343 11849 31352 11883
rect 31300 11840 31352 11849
rect 31944 11883 31996 11892
rect 31944 11849 31953 11883
rect 31953 11849 31987 11883
rect 31987 11849 31996 11883
rect 31944 11840 31996 11849
rect 32680 11840 32732 11892
rect 26056 11772 26108 11824
rect 26424 11772 26476 11824
rect 17040 11704 17092 11756
rect 19156 11704 19208 11756
rect 17224 11636 17276 11688
rect 18972 11636 19024 11688
rect 19432 11679 19484 11688
rect 19432 11645 19441 11679
rect 19441 11645 19475 11679
rect 19475 11645 19484 11679
rect 19432 11636 19484 11645
rect 19616 11679 19668 11688
rect 19616 11645 19625 11679
rect 19625 11645 19659 11679
rect 19659 11645 19668 11679
rect 19616 11636 19668 11645
rect 19340 11568 19392 11620
rect 17500 11500 17552 11552
rect 19156 11500 19208 11552
rect 22836 11704 22888 11756
rect 24216 11704 24268 11756
rect 19892 11636 19944 11688
rect 20904 11636 20956 11688
rect 21640 11679 21692 11688
rect 21640 11645 21649 11679
rect 21649 11645 21683 11679
rect 21683 11645 21692 11679
rect 21640 11636 21692 11645
rect 20536 11500 20588 11552
rect 20812 11500 20864 11552
rect 22100 11636 22152 11688
rect 24952 11679 25004 11688
rect 24952 11645 24961 11679
rect 24961 11645 24995 11679
rect 24995 11645 25004 11679
rect 24952 11636 25004 11645
rect 27804 11704 27856 11756
rect 28264 11704 28316 11756
rect 26608 11636 26660 11688
rect 28172 11636 28224 11688
rect 29184 11679 29236 11688
rect 29184 11645 29193 11679
rect 29193 11645 29227 11679
rect 29227 11645 29236 11679
rect 29184 11636 29236 11645
rect 30656 11636 30708 11688
rect 26148 11568 26200 11620
rect 28908 11568 28960 11620
rect 33508 11747 33560 11756
rect 33508 11713 33517 11747
rect 33517 11713 33551 11747
rect 33551 11713 33560 11747
rect 33508 11704 33560 11713
rect 33048 11679 33100 11688
rect 33048 11645 33057 11679
rect 33057 11645 33091 11679
rect 33091 11645 33100 11679
rect 33048 11636 33100 11645
rect 31944 11568 31996 11620
rect 29644 11500 29696 11552
rect 31208 11500 31260 11552
rect 32588 11543 32640 11552
rect 32588 11509 32597 11543
rect 32597 11509 32631 11543
rect 32631 11509 32640 11543
rect 32588 11500 32640 11509
rect 7210 11398 7262 11450
rect 7274 11398 7326 11450
rect 7338 11398 7390 11450
rect 7402 11398 7454 11450
rect 7466 11398 7518 11450
rect 15099 11398 15151 11450
rect 15163 11398 15215 11450
rect 15227 11398 15279 11450
rect 15291 11398 15343 11450
rect 15355 11398 15407 11450
rect 22988 11398 23040 11450
rect 23052 11398 23104 11450
rect 23116 11398 23168 11450
rect 23180 11398 23232 11450
rect 23244 11398 23296 11450
rect 30877 11398 30929 11450
rect 30941 11398 30993 11450
rect 31005 11398 31057 11450
rect 31069 11398 31121 11450
rect 31133 11398 31185 11450
rect 4896 11296 4948 11348
rect 1308 11228 1360 11280
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 8300 11296 8352 11348
rect 9956 11296 10008 11348
rect 10968 11296 11020 11348
rect 6092 11271 6144 11280
rect 6092 11237 6101 11271
rect 6101 11237 6135 11271
rect 6135 11237 6144 11271
rect 6092 11228 6144 11237
rect 6184 11228 6236 11280
rect 7380 11228 7432 11280
rect 7656 11271 7708 11280
rect 7656 11237 7665 11271
rect 7665 11237 7699 11271
rect 7699 11237 7708 11271
rect 7656 11228 7708 11237
rect 7748 11228 7800 11280
rect 9864 11228 9916 11280
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 3976 11024 4028 11076
rect 6920 11160 6972 11212
rect 10784 11203 10836 11212
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 13360 11296 13412 11348
rect 13728 11296 13780 11348
rect 15568 11339 15620 11348
rect 12624 11228 12676 11280
rect 12532 11203 12584 11212
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12532 11160 12584 11169
rect 13084 11160 13136 11212
rect 6276 11092 6328 11144
rect 10324 11135 10376 11144
rect 10324 11101 10333 11135
rect 10333 11101 10367 11135
rect 10367 11101 10376 11135
rect 10324 11092 10376 11101
rect 10600 11135 10652 11144
rect 10600 11101 10609 11135
rect 10609 11101 10643 11135
rect 10643 11101 10652 11135
rect 10600 11092 10652 11101
rect 11336 11092 11388 11144
rect 12900 11092 12952 11144
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 14188 11203 14240 11212
rect 14188 11169 14197 11203
rect 14197 11169 14231 11203
rect 14231 11169 14240 11203
rect 14188 11160 14240 11169
rect 14740 11203 14792 11212
rect 14740 11169 14749 11203
rect 14749 11169 14783 11203
rect 14783 11169 14792 11203
rect 15568 11305 15577 11339
rect 15577 11305 15611 11339
rect 15611 11305 15620 11339
rect 15568 11296 15620 11305
rect 15844 11296 15896 11348
rect 15936 11228 15988 11280
rect 16672 11271 16724 11280
rect 16672 11237 16681 11271
rect 16681 11237 16715 11271
rect 16715 11237 16724 11271
rect 16672 11228 16724 11237
rect 14740 11160 14792 11169
rect 17408 11160 17460 11212
rect 17500 11160 17552 11212
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 18328 11296 18380 11348
rect 19984 11339 20036 11348
rect 19984 11305 19993 11339
rect 19993 11305 20027 11339
rect 20027 11305 20036 11339
rect 19984 11296 20036 11305
rect 20996 11296 21048 11348
rect 22928 11296 22980 11348
rect 23388 11296 23440 11348
rect 26332 11296 26384 11348
rect 28172 11339 28224 11348
rect 28172 11305 28181 11339
rect 28181 11305 28215 11339
rect 28215 11305 28224 11339
rect 28172 11296 28224 11305
rect 29184 11296 29236 11348
rect 30656 11296 30708 11348
rect 30932 11296 30984 11348
rect 4712 10956 4764 11008
rect 5540 10956 5592 11008
rect 7656 10956 7708 11008
rect 8300 10956 8352 11008
rect 9680 10956 9732 11008
rect 11612 11024 11664 11076
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 11152 10999 11204 11008
rect 11152 10965 11161 10999
rect 11161 10965 11195 10999
rect 11195 10965 11204 10999
rect 11152 10956 11204 10965
rect 11520 10999 11572 11008
rect 11520 10965 11529 10999
rect 11529 10965 11563 10999
rect 11563 10965 11572 10999
rect 11520 10956 11572 10965
rect 12992 10956 13044 11008
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 13176 10956 13228 10965
rect 14004 10956 14056 11008
rect 15660 10956 15712 11008
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 17040 10999 17092 11008
rect 17040 10965 17049 10999
rect 17049 10965 17083 10999
rect 17083 10965 17092 10999
rect 17040 10956 17092 10965
rect 17224 10956 17276 11008
rect 18052 10999 18104 11008
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 18696 11024 18748 11076
rect 19432 11160 19484 11212
rect 19892 11203 19944 11212
rect 19892 11169 19901 11203
rect 19901 11169 19935 11203
rect 19935 11169 19944 11203
rect 19892 11160 19944 11169
rect 20076 11092 20128 11144
rect 27804 11228 27856 11280
rect 29644 11228 29696 11280
rect 32128 11271 32180 11280
rect 32128 11237 32137 11271
rect 32137 11237 32171 11271
rect 32171 11237 32180 11271
rect 32128 11228 32180 11237
rect 23020 11160 23072 11212
rect 23296 11160 23348 11212
rect 22652 11092 22704 11144
rect 23664 11160 23716 11212
rect 23480 11135 23532 11144
rect 23480 11101 23489 11135
rect 23489 11101 23523 11135
rect 23523 11101 23532 11135
rect 23480 11092 23532 11101
rect 24492 11092 24544 11144
rect 24860 11135 24912 11144
rect 24860 11101 24869 11135
rect 24869 11101 24903 11135
rect 24903 11101 24912 11135
rect 24860 11092 24912 11101
rect 26240 11092 26292 11144
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 28540 11160 28592 11212
rect 28724 11160 28776 11212
rect 28908 11160 28960 11212
rect 29092 11203 29144 11212
rect 29092 11169 29101 11203
rect 29101 11169 29135 11203
rect 29135 11169 29144 11203
rect 29092 11160 29144 11169
rect 26976 11092 27028 11144
rect 31208 11160 31260 11212
rect 31668 11092 31720 11144
rect 32588 11092 32640 11144
rect 19248 10956 19300 11008
rect 20996 10999 21048 11008
rect 20996 10965 21005 10999
rect 21005 10965 21039 10999
rect 21039 10965 21048 10999
rect 20996 10956 21048 10965
rect 21272 10999 21324 11008
rect 21272 10965 21281 10999
rect 21281 10965 21315 10999
rect 21315 10965 21324 10999
rect 21272 10956 21324 10965
rect 23940 10956 23992 11008
rect 24216 10999 24268 11008
rect 24216 10965 24225 10999
rect 24225 10965 24259 10999
rect 24259 10965 24268 10999
rect 24216 10956 24268 10965
rect 27344 10999 27396 11008
rect 27344 10965 27353 10999
rect 27353 10965 27387 10999
rect 27387 10965 27396 10999
rect 27344 10956 27396 10965
rect 6550 10854 6602 10906
rect 6614 10854 6666 10906
rect 6678 10854 6730 10906
rect 6742 10854 6794 10906
rect 6806 10854 6858 10906
rect 14439 10854 14491 10906
rect 14503 10854 14555 10906
rect 14567 10854 14619 10906
rect 14631 10854 14683 10906
rect 14695 10854 14747 10906
rect 22328 10854 22380 10906
rect 22392 10854 22444 10906
rect 22456 10854 22508 10906
rect 22520 10854 22572 10906
rect 22584 10854 22636 10906
rect 30217 10854 30269 10906
rect 30281 10854 30333 10906
rect 30345 10854 30397 10906
rect 30409 10854 30461 10906
rect 30473 10854 30525 10906
rect 6276 10752 6328 10804
rect 4160 10616 4212 10668
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 6644 10684 6696 10736
rect 5080 10591 5132 10600
rect 3516 10480 3568 10532
rect 4620 10480 4672 10532
rect 4160 10412 4212 10464
rect 4436 10412 4488 10464
rect 5080 10557 5081 10591
rect 5081 10557 5115 10591
rect 5115 10557 5132 10591
rect 5080 10548 5132 10557
rect 10324 10752 10376 10804
rect 11336 10795 11388 10804
rect 11336 10761 11345 10795
rect 11345 10761 11379 10795
rect 11379 10761 11388 10795
rect 11336 10752 11388 10761
rect 13176 10752 13228 10804
rect 16672 10752 16724 10804
rect 16948 10795 17000 10804
rect 16948 10761 16957 10795
rect 16957 10761 16991 10795
rect 16991 10761 17000 10795
rect 16948 10752 17000 10761
rect 18880 10795 18932 10804
rect 18880 10761 18889 10795
rect 18889 10761 18923 10795
rect 18923 10761 18932 10795
rect 18880 10752 18932 10761
rect 23480 10752 23532 10804
rect 25320 10752 25372 10804
rect 26976 10752 27028 10804
rect 28080 10752 28132 10804
rect 8116 10684 8168 10736
rect 7380 10616 7432 10668
rect 8392 10616 8444 10668
rect 8760 10548 8812 10600
rect 9128 10548 9180 10600
rect 9680 10616 9732 10668
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9864 10684 9916 10736
rect 11796 10616 11848 10668
rect 14280 10616 14332 10668
rect 14924 10684 14976 10736
rect 9588 10548 9640 10557
rect 10876 10548 10928 10600
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 5172 10455 5224 10464
rect 5172 10421 5181 10455
rect 5181 10421 5215 10455
rect 5215 10421 5224 10455
rect 5172 10412 5224 10421
rect 6092 10412 6144 10464
rect 6460 10412 6512 10464
rect 8208 10480 8260 10532
rect 8852 10480 8904 10532
rect 8484 10412 8536 10464
rect 13452 10548 13504 10600
rect 14188 10548 14240 10600
rect 16212 10616 16264 10668
rect 16488 10616 16540 10668
rect 15752 10591 15804 10600
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16304 10548 16356 10557
rect 11704 10480 11756 10532
rect 12992 10480 13044 10532
rect 13084 10480 13136 10532
rect 12532 10412 12584 10464
rect 17408 10548 17460 10600
rect 17776 10548 17828 10600
rect 18972 10548 19024 10600
rect 19156 10591 19208 10600
rect 19156 10557 19165 10591
rect 19165 10557 19199 10591
rect 19199 10557 19208 10591
rect 19156 10548 19208 10557
rect 19708 10616 19760 10668
rect 23020 10684 23072 10736
rect 20444 10548 20496 10600
rect 22836 10616 22888 10668
rect 24216 10616 24268 10668
rect 28816 10616 28868 10668
rect 34888 10616 34940 10668
rect 20996 10548 21048 10600
rect 15568 10412 15620 10464
rect 15752 10412 15804 10464
rect 15844 10455 15896 10464
rect 15844 10421 15853 10455
rect 15853 10421 15887 10455
rect 15887 10421 15896 10455
rect 15844 10412 15896 10421
rect 17592 10412 17644 10464
rect 19892 10480 19944 10532
rect 20628 10455 20680 10464
rect 20628 10421 20637 10455
rect 20637 10421 20671 10455
rect 20671 10421 20680 10455
rect 20628 10412 20680 10421
rect 22744 10548 22796 10600
rect 27804 10591 27856 10600
rect 27804 10557 27813 10591
rect 27813 10557 27847 10591
rect 27847 10557 27856 10591
rect 27804 10548 27856 10557
rect 29000 10548 29052 10600
rect 29368 10548 29420 10600
rect 29920 10591 29972 10600
rect 29920 10557 29929 10591
rect 29929 10557 29963 10591
rect 29963 10557 29972 10591
rect 29920 10548 29972 10557
rect 30012 10548 30064 10600
rect 21272 10480 21324 10532
rect 23940 10480 23992 10532
rect 25964 10480 26016 10532
rect 30932 10548 30984 10600
rect 32588 10591 32640 10600
rect 32588 10557 32597 10591
rect 32597 10557 32631 10591
rect 32631 10557 32640 10591
rect 32588 10548 32640 10557
rect 21180 10412 21232 10464
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 28908 10412 28960 10464
rect 30196 10412 30248 10464
rect 30656 10412 30708 10464
rect 7210 10310 7262 10362
rect 7274 10310 7326 10362
rect 7338 10310 7390 10362
rect 7402 10310 7454 10362
rect 7466 10310 7518 10362
rect 15099 10310 15151 10362
rect 15163 10310 15215 10362
rect 15227 10310 15279 10362
rect 15291 10310 15343 10362
rect 15355 10310 15407 10362
rect 22988 10310 23040 10362
rect 23052 10310 23104 10362
rect 23116 10310 23168 10362
rect 23180 10310 23232 10362
rect 23244 10310 23296 10362
rect 30877 10310 30929 10362
rect 30941 10310 30993 10362
rect 31005 10310 31057 10362
rect 31069 10310 31121 10362
rect 31133 10310 31185 10362
rect 3516 10208 3568 10260
rect 5356 10208 5408 10260
rect 5540 10208 5592 10260
rect 3976 10115 4028 10124
rect 3976 10081 3985 10115
rect 3985 10081 4019 10115
rect 4019 10081 4028 10115
rect 3976 10072 4028 10081
rect 4344 10115 4396 10124
rect 4344 10081 4353 10115
rect 4353 10081 4387 10115
rect 4387 10081 4396 10115
rect 4344 10072 4396 10081
rect 4620 10140 4672 10192
rect 4712 10183 4764 10192
rect 4712 10149 4721 10183
rect 4721 10149 4755 10183
rect 4755 10149 4764 10183
rect 4712 10140 4764 10149
rect 5172 10140 5224 10192
rect 6092 10208 6144 10260
rect 6368 10208 6420 10260
rect 8208 10208 8260 10260
rect 8300 10251 8352 10260
rect 8300 10217 8309 10251
rect 8309 10217 8343 10251
rect 8343 10217 8352 10251
rect 8300 10208 8352 10217
rect 8392 10208 8444 10260
rect 6552 10140 6604 10192
rect 8484 10140 8536 10192
rect 8760 10208 8812 10260
rect 10876 10208 10928 10260
rect 12532 10208 12584 10260
rect 13544 10208 13596 10260
rect 16304 10208 16356 10260
rect 17040 10251 17092 10260
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 18052 10208 18104 10260
rect 8668 10072 8720 10124
rect 9128 10140 9180 10192
rect 11520 10183 11572 10192
rect 11520 10149 11529 10183
rect 11529 10149 11563 10183
rect 11563 10149 11572 10183
rect 11520 10140 11572 10149
rect 13268 10140 13320 10192
rect 14832 10140 14884 10192
rect 15568 10140 15620 10192
rect 17224 10140 17276 10192
rect 20076 10251 20128 10260
rect 20076 10217 20085 10251
rect 20085 10217 20119 10251
rect 20119 10217 20128 10251
rect 20076 10208 20128 10217
rect 20628 10208 20680 10260
rect 22744 10208 22796 10260
rect 25044 10208 25096 10260
rect 25964 10251 26016 10260
rect 25964 10217 25973 10251
rect 25973 10217 26007 10251
rect 26007 10217 26016 10251
rect 25964 10208 26016 10217
rect 27344 10208 27396 10260
rect 29092 10208 29144 10260
rect 29736 10208 29788 10260
rect 19340 10140 19392 10192
rect 26424 10140 26476 10192
rect 30012 10140 30064 10192
rect 30196 10140 30248 10192
rect 9312 10072 9364 10124
rect 9588 10072 9640 10124
rect 10600 10072 10652 10124
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 4252 10004 4304 10056
rect 8208 10004 8260 10056
rect 8852 10004 8904 10056
rect 11152 10004 11204 10056
rect 12532 10004 12584 10056
rect 15752 10004 15804 10056
rect 16856 10004 16908 10056
rect 16948 10004 17000 10056
rect 17040 10004 17092 10056
rect 18328 10115 18380 10124
rect 18328 10081 18337 10115
rect 18337 10081 18371 10115
rect 18371 10081 18380 10115
rect 18328 10072 18380 10081
rect 22100 10072 22152 10124
rect 22744 10072 22796 10124
rect 17684 10004 17736 10056
rect 4436 9936 4488 9988
rect 7748 9936 7800 9988
rect 17408 9936 17460 9988
rect 5356 9868 5408 9920
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 9588 9868 9640 9920
rect 10876 9868 10928 9920
rect 19708 9936 19760 9988
rect 18328 9868 18380 9920
rect 20720 10047 20772 10056
rect 20720 10013 20729 10047
rect 20729 10013 20763 10047
rect 20763 10013 20772 10047
rect 20720 10004 20772 10013
rect 23940 10072 23992 10124
rect 26976 10072 27028 10124
rect 27436 10115 27488 10124
rect 27436 10081 27445 10115
rect 27445 10081 27479 10115
rect 27479 10081 27488 10115
rect 27436 10072 27488 10081
rect 28816 10072 28868 10124
rect 31208 10208 31260 10260
rect 31668 10208 31720 10260
rect 31392 10072 31444 10124
rect 23664 10047 23716 10056
rect 23664 10013 23673 10047
rect 23673 10013 23707 10047
rect 23707 10013 23716 10047
rect 23664 10004 23716 10013
rect 23756 10004 23808 10056
rect 25688 10047 25740 10056
rect 25688 10013 25697 10047
rect 25697 10013 25731 10047
rect 25731 10013 25740 10047
rect 25688 10004 25740 10013
rect 26240 10047 26292 10056
rect 26240 10013 26249 10047
rect 26249 10013 26283 10047
rect 26283 10013 26292 10047
rect 26240 10004 26292 10013
rect 26424 10047 26476 10056
rect 26424 10013 26433 10047
rect 26433 10013 26467 10047
rect 26467 10013 26476 10047
rect 26424 10004 26476 10013
rect 26516 10004 26568 10056
rect 21824 9936 21876 9988
rect 22100 9936 22152 9988
rect 23388 9936 23440 9988
rect 24860 9936 24912 9988
rect 21180 9868 21232 9920
rect 22652 9868 22704 9920
rect 22928 9911 22980 9920
rect 22928 9877 22937 9911
rect 22937 9877 22971 9911
rect 22971 9877 22980 9911
rect 22928 9868 22980 9877
rect 23296 9868 23348 9920
rect 29368 10004 29420 10056
rect 34428 10004 34480 10056
rect 25136 9911 25188 9920
rect 25136 9877 25145 9911
rect 25145 9877 25179 9911
rect 25179 9877 25188 9911
rect 25136 9868 25188 9877
rect 27160 9868 27212 9920
rect 29092 9868 29144 9920
rect 33784 9911 33836 9920
rect 33784 9877 33793 9911
rect 33793 9877 33827 9911
rect 33827 9877 33836 9911
rect 33784 9868 33836 9877
rect 6550 9766 6602 9818
rect 6614 9766 6666 9818
rect 6678 9766 6730 9818
rect 6742 9766 6794 9818
rect 6806 9766 6858 9818
rect 14439 9766 14491 9818
rect 14503 9766 14555 9818
rect 14567 9766 14619 9818
rect 14631 9766 14683 9818
rect 14695 9766 14747 9818
rect 22328 9766 22380 9818
rect 22392 9766 22444 9818
rect 22456 9766 22508 9818
rect 22520 9766 22572 9818
rect 22584 9766 22636 9818
rect 30217 9766 30269 9818
rect 30281 9766 30333 9818
rect 30345 9766 30397 9818
rect 30409 9766 30461 9818
rect 30473 9766 30525 9818
rect 3976 9664 4028 9716
rect 4712 9596 4764 9648
rect 11704 9707 11756 9716
rect 11704 9673 11713 9707
rect 11713 9673 11747 9707
rect 11747 9673 11756 9707
rect 11704 9664 11756 9673
rect 13268 9707 13320 9716
rect 13268 9673 13277 9707
rect 13277 9673 13311 9707
rect 13311 9673 13320 9707
rect 13268 9664 13320 9673
rect 14832 9707 14884 9716
rect 14832 9673 14841 9707
rect 14841 9673 14875 9707
rect 14875 9673 14884 9707
rect 14832 9664 14884 9673
rect 15752 9664 15804 9716
rect 17040 9707 17092 9716
rect 17040 9673 17049 9707
rect 17049 9673 17083 9707
rect 17083 9673 17092 9707
rect 17040 9664 17092 9673
rect 19340 9664 19392 9716
rect 1308 9528 1360 9580
rect 6092 9571 6144 9580
rect 6092 9537 6101 9571
rect 6101 9537 6135 9571
rect 6135 9537 6144 9571
rect 6092 9528 6144 9537
rect 6184 9528 6236 9580
rect 4160 9460 4212 9512
rect 5724 9503 5776 9512
rect 5724 9469 5733 9503
rect 5733 9469 5767 9503
rect 5767 9469 5776 9503
rect 5724 9460 5776 9469
rect 8576 9596 8628 9648
rect 14188 9596 14240 9648
rect 7656 9571 7708 9580
rect 7656 9537 7665 9571
rect 7665 9537 7699 9571
rect 7699 9537 7708 9571
rect 7656 9528 7708 9537
rect 8392 9528 8444 9580
rect 7564 9460 7616 9512
rect 8024 9460 8076 9512
rect 12072 9528 12124 9580
rect 3148 9324 3200 9376
rect 10692 9392 10744 9444
rect 13912 9460 13964 9512
rect 15384 9596 15436 9648
rect 17684 9596 17736 9648
rect 15844 9528 15896 9580
rect 16580 9571 16632 9580
rect 16580 9537 16589 9571
rect 16589 9537 16623 9571
rect 16623 9537 16632 9571
rect 16580 9528 16632 9537
rect 20812 9596 20864 9648
rect 20536 9528 20588 9580
rect 25136 9664 25188 9716
rect 22836 9528 22888 9580
rect 23112 9571 23164 9580
rect 23112 9537 23121 9571
rect 23121 9537 23155 9571
rect 23155 9537 23164 9571
rect 23112 9528 23164 9537
rect 28724 9664 28776 9716
rect 29000 9664 29052 9716
rect 29920 9664 29972 9716
rect 31392 9707 31444 9716
rect 31392 9673 31401 9707
rect 31401 9673 31435 9707
rect 31435 9673 31444 9707
rect 31392 9664 31444 9673
rect 25228 9596 25280 9648
rect 25504 9596 25556 9648
rect 26240 9596 26292 9648
rect 27804 9528 27856 9580
rect 17408 9460 17460 9512
rect 17592 9460 17644 9512
rect 6368 9367 6420 9376
rect 6368 9333 6377 9367
rect 6377 9333 6411 9367
rect 6411 9333 6420 9367
rect 6368 9324 6420 9333
rect 9956 9367 10008 9376
rect 9956 9333 9965 9367
rect 9965 9333 9999 9367
rect 9999 9333 10008 9367
rect 9956 9324 10008 9333
rect 10784 9324 10836 9376
rect 13084 9367 13136 9376
rect 13084 9333 13093 9367
rect 13093 9333 13127 9367
rect 13127 9333 13136 9367
rect 13084 9324 13136 9333
rect 13268 9324 13320 9376
rect 16764 9392 16816 9444
rect 18144 9392 18196 9444
rect 18604 9392 18656 9444
rect 19248 9460 19300 9512
rect 20352 9503 20404 9512
rect 20352 9469 20361 9503
rect 20361 9469 20395 9503
rect 20395 9469 20404 9503
rect 20352 9460 20404 9469
rect 15752 9324 15804 9376
rect 16672 9324 16724 9376
rect 17592 9324 17644 9376
rect 19340 9324 19392 9376
rect 20444 9324 20496 9376
rect 20904 9367 20956 9376
rect 20904 9333 20913 9367
rect 20913 9333 20947 9367
rect 20947 9333 20956 9367
rect 20904 9324 20956 9333
rect 22928 9460 22980 9512
rect 23756 9460 23808 9512
rect 23848 9503 23900 9512
rect 23848 9469 23857 9503
rect 23857 9469 23891 9503
rect 23891 9469 23900 9503
rect 23848 9460 23900 9469
rect 21732 9392 21784 9444
rect 22192 9392 22244 9444
rect 21824 9367 21876 9376
rect 21824 9333 21833 9367
rect 21833 9333 21867 9367
rect 21867 9333 21876 9367
rect 21824 9324 21876 9333
rect 22652 9324 22704 9376
rect 25412 9392 25464 9444
rect 27160 9392 27212 9444
rect 28540 9392 28592 9444
rect 26332 9324 26384 9376
rect 26792 9324 26844 9376
rect 33968 9596 34020 9648
rect 29000 9571 29052 9580
rect 29000 9537 29009 9571
rect 29009 9537 29043 9571
rect 29043 9537 29052 9571
rect 29000 9528 29052 9537
rect 29552 9528 29604 9580
rect 29092 9460 29144 9512
rect 28724 9367 28776 9376
rect 28724 9333 28733 9367
rect 28733 9333 28767 9367
rect 28767 9333 28776 9367
rect 28724 9324 28776 9333
rect 28816 9324 28868 9376
rect 7210 9222 7262 9274
rect 7274 9222 7326 9274
rect 7338 9222 7390 9274
rect 7402 9222 7454 9274
rect 7466 9222 7518 9274
rect 15099 9222 15151 9274
rect 15163 9222 15215 9274
rect 15227 9222 15279 9274
rect 15291 9222 15343 9274
rect 15355 9222 15407 9274
rect 22988 9222 23040 9274
rect 23052 9222 23104 9274
rect 23116 9222 23168 9274
rect 23180 9222 23232 9274
rect 23244 9222 23296 9274
rect 30877 9222 30929 9274
rect 30941 9222 30993 9274
rect 31005 9222 31057 9274
rect 31069 9222 31121 9274
rect 31133 9222 31185 9274
rect 4252 9120 4304 9172
rect 3240 9052 3292 9104
rect 6000 9052 6052 9104
rect 4436 8984 4488 9036
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 5356 9027 5408 9036
rect 5356 8993 5365 9027
rect 5365 8993 5399 9027
rect 5399 8993 5408 9027
rect 5356 8984 5408 8993
rect 7012 9120 7064 9172
rect 10232 9163 10284 9172
rect 10232 9129 10241 9163
rect 10241 9129 10275 9163
rect 10275 9129 10284 9163
rect 10232 9120 10284 9129
rect 10416 9120 10468 9172
rect 10692 9120 10744 9172
rect 13268 9120 13320 9172
rect 9772 9052 9824 9104
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 8484 8984 8536 9036
rect 11520 9052 11572 9104
rect 14188 9052 14240 9104
rect 14372 9052 14424 9104
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 9956 8916 10008 8968
rect 12256 8959 12308 8968
rect 12256 8925 12265 8959
rect 12265 8925 12299 8959
rect 12299 8925 12308 8959
rect 12256 8916 12308 8925
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 17592 8984 17644 9036
rect 18052 9120 18104 9172
rect 17868 9052 17920 9104
rect 20352 9120 20404 9172
rect 20720 9120 20772 9172
rect 25136 9120 25188 9172
rect 25688 9120 25740 9172
rect 26240 9120 26292 9172
rect 26332 9120 26384 9172
rect 27896 9120 27948 9172
rect 28724 9120 28776 9172
rect 29552 9163 29604 9172
rect 29552 9129 29561 9163
rect 29561 9129 29595 9163
rect 29595 9129 29604 9163
rect 29552 9120 29604 9129
rect 29736 9120 29788 9172
rect 18788 9027 18840 9036
rect 18788 8993 18797 9027
rect 18797 8993 18831 9027
rect 18831 8993 18840 9027
rect 18788 8984 18840 8993
rect 19616 9027 19668 9036
rect 19616 8993 19650 9027
rect 19650 8993 19668 9027
rect 19616 8984 19668 8993
rect 20904 8984 20956 9036
rect 14556 8916 14608 8968
rect 16948 8916 17000 8968
rect 16856 8848 16908 8900
rect 17132 8848 17184 8900
rect 18512 8916 18564 8968
rect 19156 8916 19208 8968
rect 19524 8959 19576 8968
rect 19524 8925 19533 8959
rect 19533 8925 19567 8959
rect 19567 8925 19576 8959
rect 19524 8916 19576 8925
rect 19340 8848 19392 8900
rect 3424 8780 3476 8832
rect 4436 8823 4488 8832
rect 4436 8789 4445 8823
rect 4445 8789 4479 8823
rect 4479 8789 4488 8823
rect 4436 8780 4488 8789
rect 5356 8780 5408 8832
rect 5908 8780 5960 8832
rect 8024 8780 8076 8832
rect 9312 8780 9364 8832
rect 9496 8823 9548 8832
rect 9496 8789 9505 8823
rect 9505 8789 9539 8823
rect 9539 8789 9548 8823
rect 9496 8780 9548 8789
rect 13912 8780 13964 8832
rect 14832 8780 14884 8832
rect 15936 8780 15988 8832
rect 16580 8780 16632 8832
rect 18144 8780 18196 8832
rect 18972 8780 19024 8832
rect 23572 8984 23624 9036
rect 21180 8916 21232 8968
rect 21824 8959 21876 8968
rect 21824 8925 21833 8959
rect 21833 8925 21867 8959
rect 21867 8925 21876 8959
rect 21824 8916 21876 8925
rect 24860 8984 24912 9036
rect 23940 8848 23992 8900
rect 22008 8780 22060 8832
rect 24952 8916 25004 8968
rect 25228 8984 25280 9036
rect 25412 9027 25464 9036
rect 25412 8993 25421 9027
rect 25421 8993 25455 9027
rect 25455 8993 25464 9027
rect 25412 8984 25464 8993
rect 26792 8984 26844 9036
rect 25688 8959 25740 8968
rect 25688 8925 25697 8959
rect 25697 8925 25731 8959
rect 25731 8925 25740 8959
rect 25688 8916 25740 8925
rect 25872 8959 25924 8968
rect 25872 8925 25881 8959
rect 25881 8925 25915 8959
rect 25915 8925 25924 8959
rect 25872 8916 25924 8925
rect 26608 8959 26660 8968
rect 26608 8925 26617 8959
rect 26617 8925 26651 8959
rect 26651 8925 26660 8959
rect 26608 8916 26660 8925
rect 26884 8959 26936 8968
rect 26884 8925 26893 8959
rect 26893 8925 26927 8959
rect 26927 8925 26936 8959
rect 26884 8916 26936 8925
rect 28448 8959 28500 8968
rect 28448 8925 28457 8959
rect 28457 8925 28491 8959
rect 28491 8925 28500 8959
rect 28448 8916 28500 8925
rect 28540 8916 28592 8968
rect 25320 8848 25372 8900
rect 27528 8823 27580 8832
rect 27528 8789 27537 8823
rect 27537 8789 27571 8823
rect 27571 8789 27580 8823
rect 27528 8780 27580 8789
rect 27620 8780 27672 8832
rect 29920 8959 29972 8968
rect 29920 8925 29929 8959
rect 29929 8925 29963 8959
rect 29963 8925 29972 8959
rect 29920 8916 29972 8925
rect 30656 8780 30708 8832
rect 32588 8959 32640 8968
rect 32588 8925 32597 8959
rect 32597 8925 32631 8959
rect 32631 8925 32640 8959
rect 32588 8916 32640 8925
rect 33416 8848 33468 8900
rect 32036 8823 32088 8832
rect 32036 8789 32045 8823
rect 32045 8789 32079 8823
rect 32079 8789 32088 8823
rect 32036 8780 32088 8789
rect 6550 8678 6602 8730
rect 6614 8678 6666 8730
rect 6678 8678 6730 8730
rect 6742 8678 6794 8730
rect 6806 8678 6858 8730
rect 14439 8678 14491 8730
rect 14503 8678 14555 8730
rect 14567 8678 14619 8730
rect 14631 8678 14683 8730
rect 14695 8678 14747 8730
rect 22328 8678 22380 8730
rect 22392 8678 22444 8730
rect 22456 8678 22508 8730
rect 22520 8678 22572 8730
rect 22584 8678 22636 8730
rect 30217 8678 30269 8730
rect 30281 8678 30333 8730
rect 30345 8678 30397 8730
rect 30409 8678 30461 8730
rect 30473 8678 30525 8730
rect 3424 8576 3476 8628
rect 5080 8619 5132 8628
rect 5080 8585 5089 8619
rect 5089 8585 5123 8619
rect 5123 8585 5132 8619
rect 5080 8576 5132 8585
rect 5264 8576 5316 8628
rect 5908 8576 5960 8628
rect 7104 8576 7156 8628
rect 8300 8576 8352 8628
rect 13084 8576 13136 8628
rect 13728 8576 13780 8628
rect 14188 8576 14240 8628
rect 14832 8576 14884 8628
rect 18880 8619 18932 8628
rect 4344 8440 4396 8492
rect 11520 8551 11572 8560
rect 11520 8517 11529 8551
rect 11529 8517 11563 8551
rect 11563 8517 11572 8551
rect 11520 8508 11572 8517
rect 11796 8508 11848 8560
rect 12164 8508 12216 8560
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 13820 8440 13872 8492
rect 14096 8440 14148 8492
rect 4436 8372 4488 8424
rect 5816 8372 5868 8424
rect 9680 8372 9732 8424
rect 12072 8372 12124 8424
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 18880 8585 18889 8619
rect 18889 8585 18923 8619
rect 18923 8585 18932 8619
rect 18880 8576 18932 8585
rect 19340 8576 19392 8628
rect 19616 8576 19668 8628
rect 15936 8483 15988 8492
rect 15936 8449 15945 8483
rect 15945 8449 15979 8483
rect 15979 8449 15988 8483
rect 15936 8440 15988 8449
rect 16672 8440 16724 8492
rect 16948 8508 17000 8560
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 17224 8415 17276 8424
rect 17224 8381 17258 8415
rect 17258 8381 17276 8415
rect 18972 8508 19024 8560
rect 17776 8440 17828 8492
rect 18144 8440 18196 8492
rect 19248 8483 19300 8492
rect 19248 8449 19257 8483
rect 19257 8449 19291 8483
rect 19291 8449 19300 8483
rect 19248 8440 19300 8449
rect 17224 8372 17276 8381
rect 17960 8415 18012 8424
rect 17960 8381 17969 8415
rect 17969 8381 18003 8415
rect 18003 8381 18012 8415
rect 17960 8372 18012 8381
rect 7656 8347 7708 8356
rect 7656 8313 7665 8347
rect 7665 8313 7699 8347
rect 7699 8313 7708 8347
rect 7656 8304 7708 8313
rect 9496 8304 9548 8356
rect 12532 8304 12584 8356
rect 13912 8304 13964 8356
rect 4804 8279 4856 8288
rect 4804 8245 4813 8279
rect 4813 8245 4847 8279
rect 4847 8245 4856 8279
rect 4804 8236 4856 8245
rect 6184 8236 6236 8288
rect 6552 8236 6604 8288
rect 9220 8279 9272 8288
rect 9220 8245 9229 8279
rect 9229 8245 9263 8279
rect 9263 8245 9272 8279
rect 9220 8236 9272 8245
rect 14924 8236 14976 8288
rect 16580 8304 16632 8356
rect 21732 8576 21784 8628
rect 22100 8576 22152 8628
rect 20812 8508 20864 8560
rect 22836 8576 22888 8628
rect 23388 8508 23440 8560
rect 23572 8619 23624 8628
rect 23572 8585 23581 8619
rect 23581 8585 23615 8619
rect 23615 8585 23624 8619
rect 23572 8576 23624 8585
rect 24216 8576 24268 8628
rect 25320 8619 25372 8628
rect 25320 8585 25329 8619
rect 25329 8585 25363 8619
rect 25363 8585 25372 8619
rect 25320 8576 25372 8585
rect 25688 8576 25740 8628
rect 26332 8576 26384 8628
rect 26700 8508 26752 8560
rect 26884 8508 26936 8560
rect 27436 8576 27488 8628
rect 28448 8576 28500 8628
rect 29000 8576 29052 8628
rect 29460 8576 29512 8628
rect 29920 8576 29972 8628
rect 33508 8576 33560 8628
rect 21640 8440 21692 8492
rect 21732 8483 21784 8492
rect 21732 8449 21741 8483
rect 21741 8449 21775 8483
rect 21775 8449 21784 8483
rect 21732 8440 21784 8449
rect 21824 8440 21876 8492
rect 19800 8415 19852 8424
rect 19800 8381 19809 8415
rect 19809 8381 19843 8415
rect 19843 8381 19852 8415
rect 19800 8372 19852 8381
rect 20536 8372 20588 8424
rect 21088 8415 21140 8424
rect 21088 8381 21097 8415
rect 21097 8381 21131 8415
rect 21131 8381 21140 8415
rect 21088 8372 21140 8381
rect 23112 8440 23164 8492
rect 22284 8415 22336 8424
rect 22284 8381 22293 8415
rect 22293 8381 22327 8415
rect 22327 8381 22336 8415
rect 22284 8372 22336 8381
rect 24860 8415 24912 8424
rect 24860 8381 24869 8415
rect 24869 8381 24903 8415
rect 24903 8381 24912 8415
rect 24860 8372 24912 8381
rect 25228 8372 25280 8424
rect 26332 8372 26384 8424
rect 26516 8372 26568 8424
rect 26884 8372 26936 8424
rect 27068 8415 27120 8424
rect 27068 8381 27077 8415
rect 27077 8381 27111 8415
rect 27111 8381 27120 8415
rect 27068 8372 27120 8381
rect 27436 8372 27488 8424
rect 27528 8415 27580 8424
rect 27528 8381 27537 8415
rect 27537 8381 27571 8415
rect 27571 8381 27580 8415
rect 27528 8372 27580 8381
rect 27896 8440 27948 8492
rect 33784 8551 33836 8560
rect 33784 8517 33793 8551
rect 33793 8517 33827 8551
rect 33827 8517 33836 8551
rect 33784 8508 33836 8517
rect 28172 8440 28224 8492
rect 15384 8279 15436 8288
rect 15384 8245 15409 8279
rect 15409 8245 15436 8279
rect 15384 8236 15436 8245
rect 15568 8279 15620 8288
rect 15568 8245 15577 8279
rect 15577 8245 15611 8279
rect 15611 8245 15620 8279
rect 15568 8236 15620 8245
rect 17408 8236 17460 8288
rect 17684 8236 17736 8288
rect 19432 8236 19484 8288
rect 20996 8236 21048 8288
rect 25688 8304 25740 8356
rect 27712 8304 27764 8356
rect 28724 8415 28776 8424
rect 28724 8381 28733 8415
rect 28733 8381 28767 8415
rect 28767 8381 28776 8415
rect 28724 8372 28776 8381
rect 29000 8415 29052 8424
rect 29000 8381 29009 8415
rect 29009 8381 29043 8415
rect 29043 8381 29052 8415
rect 29000 8372 29052 8381
rect 31208 8483 31260 8492
rect 31208 8449 31217 8483
rect 31217 8449 31251 8483
rect 31251 8449 31260 8483
rect 31208 8440 31260 8449
rect 24308 8279 24360 8288
rect 24308 8245 24317 8279
rect 24317 8245 24351 8279
rect 24351 8245 24360 8279
rect 24308 8236 24360 8245
rect 24492 8236 24544 8288
rect 26884 8236 26936 8288
rect 26976 8279 27028 8288
rect 26976 8245 26985 8279
rect 26985 8245 27019 8279
rect 27019 8245 27028 8279
rect 26976 8236 27028 8245
rect 28172 8236 28224 8288
rect 29092 8304 29144 8356
rect 29276 8347 29328 8356
rect 29276 8313 29285 8347
rect 29285 8313 29319 8347
rect 29319 8313 29328 8347
rect 29276 8304 29328 8313
rect 29460 8372 29512 8424
rect 31576 8415 31628 8424
rect 31576 8381 31585 8415
rect 31585 8381 31619 8415
rect 31619 8381 31628 8415
rect 31576 8372 31628 8381
rect 29828 8304 29880 8356
rect 34428 8304 34480 8356
rect 31852 8236 31904 8288
rect 7210 8134 7262 8186
rect 7274 8134 7326 8186
rect 7338 8134 7390 8186
rect 7402 8134 7454 8186
rect 7466 8134 7518 8186
rect 15099 8134 15151 8186
rect 15163 8134 15215 8186
rect 15227 8134 15279 8186
rect 15291 8134 15343 8186
rect 15355 8134 15407 8186
rect 22988 8134 23040 8186
rect 23052 8134 23104 8186
rect 23116 8134 23168 8186
rect 23180 8134 23232 8186
rect 23244 8134 23296 8186
rect 30877 8134 30929 8186
rect 30941 8134 30993 8186
rect 31005 8134 31057 8186
rect 31069 8134 31121 8186
rect 31133 8134 31185 8186
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 4160 8032 4212 8084
rect 4252 8032 4304 8084
rect 5816 8032 5868 8084
rect 6276 8032 6328 8084
rect 7656 8032 7708 8084
rect 8484 8075 8536 8084
rect 8484 8041 8493 8075
rect 8493 8041 8527 8075
rect 8527 8041 8536 8075
rect 8484 8032 8536 8041
rect 9220 8032 9272 8084
rect 9680 8032 9732 8084
rect 11704 8032 11756 8084
rect 11980 8032 12032 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 12532 8032 12584 8084
rect 1308 7896 1360 7948
rect 4068 7828 4120 7880
rect 4436 7828 4488 7880
rect 4804 7828 4856 7880
rect 5356 7828 5408 7880
rect 5724 7896 5776 7948
rect 14188 7964 14240 8016
rect 14924 8032 14976 8084
rect 6276 7939 6328 7948
rect 6276 7905 6285 7939
rect 6285 7905 6319 7939
rect 6319 7905 6328 7939
rect 6276 7896 6328 7905
rect 6460 7896 6512 7948
rect 8668 7896 8720 7948
rect 8852 7896 8904 7948
rect 9220 7939 9272 7948
rect 9220 7905 9229 7939
rect 9229 7905 9263 7939
rect 9263 7905 9272 7939
rect 9220 7896 9272 7905
rect 10048 7896 10100 7948
rect 10508 7896 10560 7948
rect 10784 7896 10836 7948
rect 11612 7939 11664 7948
rect 11612 7905 11621 7939
rect 11621 7905 11655 7939
rect 11655 7905 11664 7939
rect 11612 7896 11664 7905
rect 11796 7939 11848 7948
rect 11796 7905 11805 7939
rect 11805 7905 11839 7939
rect 11839 7905 11848 7939
rect 11796 7896 11848 7905
rect 11888 7939 11940 7948
rect 11888 7905 11897 7939
rect 11897 7905 11931 7939
rect 11931 7905 11940 7939
rect 11888 7896 11940 7905
rect 11980 7939 12032 7948
rect 11980 7905 11989 7939
rect 11989 7905 12023 7939
rect 12023 7905 12032 7939
rect 11980 7896 12032 7905
rect 15292 7964 15344 8016
rect 15752 8032 15804 8084
rect 16764 8032 16816 8084
rect 17132 8032 17184 8084
rect 17960 8032 18012 8084
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 9680 7828 9732 7880
rect 8208 7760 8260 7812
rect 9312 7760 9364 7812
rect 10232 7871 10284 7880
rect 10232 7837 10241 7871
rect 10241 7837 10275 7871
rect 10275 7837 10284 7871
rect 10232 7828 10284 7837
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 8576 7692 8628 7744
rect 9956 7692 10008 7744
rect 10416 7735 10468 7744
rect 10416 7701 10425 7735
rect 10425 7701 10459 7735
rect 10459 7701 10468 7735
rect 10416 7692 10468 7701
rect 11888 7760 11940 7812
rect 13636 7828 13688 7880
rect 14280 7828 14332 7880
rect 14740 7939 14792 7948
rect 14740 7905 14749 7939
rect 14749 7905 14783 7939
rect 14783 7905 14792 7939
rect 14740 7896 14792 7905
rect 16672 7896 16724 7948
rect 17684 7964 17736 8016
rect 17776 8007 17828 8016
rect 17776 7973 17785 8007
rect 17785 7973 17819 8007
rect 17819 7973 17828 8007
rect 17776 7964 17828 7973
rect 15752 7828 15804 7880
rect 17224 7828 17276 7880
rect 17316 7828 17368 7880
rect 18696 7896 18748 7948
rect 19984 8032 20036 8084
rect 19248 7964 19300 8016
rect 21456 7964 21508 8016
rect 21640 7964 21692 8016
rect 11612 7692 11664 7744
rect 12164 7735 12216 7744
rect 12164 7701 12173 7735
rect 12173 7701 12207 7735
rect 12207 7701 12216 7735
rect 12164 7692 12216 7701
rect 14004 7692 14056 7744
rect 18604 7760 18656 7812
rect 19156 7939 19208 7948
rect 19156 7905 19165 7939
rect 19165 7905 19199 7939
rect 19199 7905 19208 7939
rect 19156 7896 19208 7905
rect 22836 8032 22888 8084
rect 23388 8032 23440 8084
rect 24308 8032 24360 8084
rect 24952 8032 25004 8084
rect 26424 8032 26476 8084
rect 27896 8032 27948 8084
rect 29092 8032 29144 8084
rect 30196 8032 30248 8084
rect 32588 8032 32640 8084
rect 25412 7964 25464 8016
rect 28816 7964 28868 8016
rect 21732 7896 21784 7948
rect 22652 7896 22704 7948
rect 22744 7896 22796 7948
rect 25504 7896 25556 7948
rect 19708 7803 19760 7812
rect 19708 7769 19717 7803
rect 19717 7769 19751 7803
rect 19751 7769 19760 7803
rect 19708 7760 19760 7769
rect 23572 7828 23624 7880
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 24768 7828 24820 7880
rect 26424 7871 26476 7880
rect 26424 7837 26433 7871
rect 26433 7837 26467 7871
rect 26467 7837 26476 7871
rect 26424 7828 26476 7837
rect 27804 7828 27856 7880
rect 28908 7871 28960 7880
rect 28908 7837 28917 7871
rect 28917 7837 28951 7871
rect 28951 7837 28960 7871
rect 28908 7828 28960 7837
rect 30564 7896 30616 7948
rect 32588 7896 32640 7948
rect 33416 7939 33468 7948
rect 33416 7905 33425 7939
rect 33425 7905 33459 7939
rect 33459 7905 33468 7939
rect 33416 7896 33468 7905
rect 15200 7692 15252 7744
rect 16764 7692 16816 7744
rect 18420 7735 18472 7744
rect 18420 7701 18429 7735
rect 18429 7701 18463 7735
rect 18463 7701 18472 7735
rect 18420 7692 18472 7701
rect 19340 7692 19392 7744
rect 21180 7735 21232 7744
rect 21180 7701 21189 7735
rect 21189 7701 21223 7735
rect 21223 7701 21232 7735
rect 21180 7692 21232 7701
rect 21548 7692 21600 7744
rect 22008 7692 22060 7744
rect 22652 7692 22704 7744
rect 22744 7735 22796 7744
rect 22744 7701 22753 7735
rect 22753 7701 22787 7735
rect 22787 7701 22796 7735
rect 23756 7735 23808 7744
rect 22744 7692 22796 7701
rect 23756 7701 23765 7735
rect 23765 7701 23799 7735
rect 23799 7701 23808 7735
rect 23756 7692 23808 7701
rect 30748 7828 30800 7880
rect 32312 7828 32364 7880
rect 32680 7871 32732 7880
rect 32680 7837 32689 7871
rect 32689 7837 32723 7871
rect 32723 7837 32732 7871
rect 32680 7828 32732 7837
rect 33508 7828 33560 7880
rect 30012 7692 30064 7744
rect 6550 7590 6602 7642
rect 6614 7590 6666 7642
rect 6678 7590 6730 7642
rect 6742 7590 6794 7642
rect 6806 7590 6858 7642
rect 14439 7590 14491 7642
rect 14503 7590 14555 7642
rect 14567 7590 14619 7642
rect 14631 7590 14683 7642
rect 14695 7590 14747 7642
rect 22328 7590 22380 7642
rect 22392 7590 22444 7642
rect 22456 7590 22508 7642
rect 22520 7590 22572 7642
rect 22584 7590 22636 7642
rect 30217 7590 30269 7642
rect 30281 7590 30333 7642
rect 30345 7590 30397 7642
rect 30409 7590 30461 7642
rect 30473 7590 30525 7642
rect 3516 7395 3568 7404
rect 3516 7361 3525 7395
rect 3525 7361 3559 7395
rect 3559 7361 3568 7395
rect 3516 7352 3568 7361
rect 9036 7488 9088 7540
rect 10140 7531 10192 7540
rect 10140 7497 10149 7531
rect 10149 7497 10183 7531
rect 10183 7497 10192 7531
rect 10140 7488 10192 7497
rect 10600 7488 10652 7540
rect 12164 7531 12216 7540
rect 12164 7497 12194 7531
rect 12194 7497 12216 7531
rect 12164 7488 12216 7497
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 14096 7488 14148 7540
rect 15476 7488 15528 7540
rect 15752 7531 15804 7540
rect 15752 7497 15761 7531
rect 15761 7497 15795 7531
rect 15795 7497 15804 7531
rect 15752 7488 15804 7497
rect 16672 7531 16724 7540
rect 16672 7497 16681 7531
rect 16681 7497 16715 7531
rect 16715 7497 16724 7531
rect 16672 7488 16724 7497
rect 6092 7420 6144 7472
rect 3148 7327 3200 7336
rect 3148 7293 3157 7327
rect 3157 7293 3191 7327
rect 3191 7293 3200 7327
rect 3148 7284 3200 7293
rect 5448 7284 5500 7336
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 6460 7352 6512 7404
rect 9312 7352 9364 7404
rect 8300 7284 8352 7336
rect 10416 7420 10468 7472
rect 12256 7352 12308 7404
rect 14832 7420 14884 7472
rect 10784 7284 10836 7336
rect 13820 7284 13872 7336
rect 15568 7352 15620 7404
rect 15292 7284 15344 7336
rect 15476 7284 15528 7336
rect 15936 7284 15988 7336
rect 17316 7488 17368 7540
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 19708 7488 19760 7540
rect 22008 7488 22060 7540
rect 17408 7352 17460 7404
rect 21272 7420 21324 7472
rect 21916 7420 21968 7472
rect 16764 7327 16816 7336
rect 16764 7293 16773 7327
rect 16773 7293 16807 7327
rect 16807 7293 16816 7327
rect 16764 7284 16816 7293
rect 16948 7284 17000 7336
rect 18420 7284 18472 7336
rect 20260 7284 20312 7336
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 5264 7148 5316 7200
rect 15200 7216 15252 7268
rect 20352 7216 20404 7268
rect 21272 7284 21324 7336
rect 23388 7488 23440 7540
rect 24860 7488 24912 7540
rect 25412 7531 25464 7540
rect 25412 7497 25421 7531
rect 25421 7497 25455 7531
rect 25455 7497 25464 7531
rect 25412 7488 25464 7497
rect 26424 7488 26476 7540
rect 28816 7488 28868 7540
rect 28908 7488 28960 7540
rect 30012 7488 30064 7540
rect 30656 7488 30708 7540
rect 31852 7488 31904 7540
rect 24124 7420 24176 7472
rect 23848 7352 23900 7404
rect 24952 7395 25004 7404
rect 24952 7361 24961 7395
rect 24961 7361 24995 7395
rect 24995 7361 25004 7395
rect 24952 7352 25004 7361
rect 27804 7395 27856 7404
rect 27804 7361 27813 7395
rect 27813 7361 27847 7395
rect 27847 7361 27856 7395
rect 27804 7352 27856 7361
rect 30196 7352 30248 7404
rect 6552 7148 6604 7200
rect 8668 7148 8720 7200
rect 9036 7148 9088 7200
rect 9680 7148 9732 7200
rect 10232 7148 10284 7200
rect 10508 7148 10560 7200
rect 11428 7191 11480 7200
rect 11428 7157 11437 7191
rect 11437 7157 11471 7191
rect 11471 7157 11480 7191
rect 11428 7148 11480 7157
rect 11980 7148 12032 7200
rect 13544 7148 13596 7200
rect 14280 7148 14332 7200
rect 19432 7148 19484 7200
rect 19892 7148 19944 7200
rect 21732 7216 21784 7268
rect 22468 7284 22520 7336
rect 20720 7148 20772 7200
rect 20996 7148 21048 7200
rect 22100 7148 22152 7200
rect 25136 7216 25188 7268
rect 25228 7216 25280 7268
rect 26976 7216 27028 7268
rect 27620 7216 27672 7268
rect 23480 7148 23532 7200
rect 24308 7191 24360 7200
rect 24308 7157 24317 7191
rect 24317 7157 24351 7191
rect 24351 7157 24360 7191
rect 24308 7148 24360 7157
rect 24860 7191 24912 7200
rect 24860 7157 24869 7191
rect 24869 7157 24903 7191
rect 24903 7157 24912 7191
rect 24860 7148 24912 7157
rect 25780 7191 25832 7200
rect 25780 7157 25789 7191
rect 25789 7157 25823 7191
rect 25823 7157 25832 7191
rect 25780 7148 25832 7157
rect 27436 7148 27488 7200
rect 28172 7284 28224 7336
rect 31208 7352 31260 7404
rect 32036 7395 32088 7404
rect 32036 7361 32045 7395
rect 32045 7361 32079 7395
rect 32079 7361 32088 7395
rect 32036 7352 32088 7361
rect 32312 7216 32364 7268
rect 33692 7216 33744 7268
rect 31208 7148 31260 7200
rect 7210 7046 7262 7098
rect 7274 7046 7326 7098
rect 7338 7046 7390 7098
rect 7402 7046 7454 7098
rect 7466 7046 7518 7098
rect 15099 7046 15151 7098
rect 15163 7046 15215 7098
rect 15227 7046 15279 7098
rect 15291 7046 15343 7098
rect 15355 7046 15407 7098
rect 22988 7046 23040 7098
rect 23052 7046 23104 7098
rect 23116 7046 23168 7098
rect 23180 7046 23232 7098
rect 23244 7046 23296 7098
rect 30877 7046 30929 7098
rect 30941 7046 30993 7098
rect 31005 7046 31057 7098
rect 31069 7046 31121 7098
rect 31133 7046 31185 7098
rect 5264 6944 5316 6996
rect 6092 6987 6144 6996
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 12440 6944 12492 6996
rect 12900 6987 12952 6996
rect 12900 6953 12909 6987
rect 12909 6953 12943 6987
rect 12943 6953 12952 6987
rect 12900 6944 12952 6953
rect 14188 6944 14240 6996
rect 18696 6944 18748 6996
rect 19340 6944 19392 6996
rect 20352 6944 20404 6996
rect 3148 6876 3200 6928
rect 4620 6876 4672 6928
rect 6276 6876 6328 6928
rect 7104 6876 7156 6928
rect 15936 6876 15988 6928
rect 20720 6876 20772 6928
rect 23572 6944 23624 6996
rect 24860 6944 24912 6996
rect 26516 6987 26568 6996
rect 26516 6953 26525 6987
rect 26525 6953 26559 6987
rect 26559 6953 26568 6987
rect 26516 6944 26568 6953
rect 27620 6944 27672 6996
rect 30104 6944 30156 6996
rect 30748 6944 30800 6996
rect 3884 6740 3936 6792
rect 4252 6851 4304 6860
rect 4252 6817 4261 6851
rect 4261 6817 4295 6851
rect 4295 6817 4304 6851
rect 4252 6808 4304 6817
rect 8392 6808 8444 6860
rect 10508 6808 10560 6860
rect 11428 6808 11480 6860
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 16580 6808 16632 6860
rect 18052 6808 18104 6860
rect 20996 6808 21048 6860
rect 22100 6851 22152 6860
rect 22100 6817 22109 6851
rect 22109 6817 22143 6851
rect 22143 6817 22152 6851
rect 22100 6808 22152 6817
rect 22192 6808 22244 6860
rect 5264 6740 5316 6792
rect 7472 6740 7524 6792
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 5264 6604 5316 6656
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6000 6604 6052 6613
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 16948 6740 17000 6792
rect 18788 6740 18840 6792
rect 19064 6740 19116 6792
rect 23756 6808 23808 6860
rect 24124 6808 24176 6860
rect 25780 6876 25832 6928
rect 25412 6808 25464 6860
rect 25504 6851 25556 6860
rect 25504 6817 25513 6851
rect 25513 6817 25547 6851
rect 25547 6817 25556 6851
rect 25504 6808 25556 6817
rect 10140 6604 10192 6656
rect 10232 6604 10284 6656
rect 11704 6647 11756 6656
rect 11704 6613 11713 6647
rect 11713 6613 11747 6647
rect 11747 6613 11756 6647
rect 11704 6604 11756 6613
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 19340 6604 19392 6656
rect 19616 6647 19668 6656
rect 19616 6613 19625 6647
rect 19625 6613 19659 6647
rect 19659 6613 19668 6647
rect 19616 6604 19668 6613
rect 23020 6783 23072 6792
rect 23020 6749 23029 6783
rect 23029 6749 23063 6783
rect 23063 6749 23072 6783
rect 23020 6740 23072 6749
rect 25688 6783 25740 6792
rect 25688 6749 25697 6783
rect 25697 6749 25731 6783
rect 25731 6749 25740 6783
rect 25688 6740 25740 6749
rect 26332 6783 26384 6792
rect 26332 6749 26341 6783
rect 26341 6749 26375 6783
rect 26375 6749 26384 6783
rect 26332 6740 26384 6749
rect 27712 6808 27764 6860
rect 27988 6851 28040 6860
rect 27988 6817 27997 6851
rect 27997 6817 28031 6851
rect 28031 6817 28040 6851
rect 27988 6808 28040 6817
rect 28632 6851 28684 6860
rect 28632 6817 28641 6851
rect 28641 6817 28675 6851
rect 28675 6817 28684 6851
rect 28632 6808 28684 6817
rect 30564 6808 30616 6860
rect 32680 6944 32732 6996
rect 28448 6672 28500 6724
rect 29460 6672 29512 6724
rect 21180 6604 21232 6656
rect 21548 6647 21600 6656
rect 21548 6613 21557 6647
rect 21557 6613 21591 6647
rect 21591 6613 21600 6647
rect 21548 6604 21600 6613
rect 22468 6647 22520 6656
rect 22468 6613 22477 6647
rect 22477 6613 22511 6647
rect 22511 6613 22520 6647
rect 22468 6604 22520 6613
rect 22836 6604 22888 6656
rect 24768 6647 24820 6656
rect 24768 6613 24777 6647
rect 24777 6613 24811 6647
rect 24811 6613 24820 6647
rect 24768 6604 24820 6613
rect 24860 6604 24912 6656
rect 26240 6604 26292 6656
rect 30012 6604 30064 6656
rect 30196 6604 30248 6656
rect 30748 6604 30800 6656
rect 31208 6740 31260 6792
rect 32312 6851 32364 6860
rect 32312 6817 32321 6851
rect 32321 6817 32355 6851
rect 32355 6817 32364 6851
rect 32312 6808 32364 6817
rect 34704 6808 34756 6860
rect 31484 6647 31536 6656
rect 31484 6613 31493 6647
rect 31493 6613 31527 6647
rect 31527 6613 31536 6647
rect 32036 6672 32088 6724
rect 31484 6604 31536 6613
rect 6550 6502 6602 6554
rect 6614 6502 6666 6554
rect 6678 6502 6730 6554
rect 6742 6502 6794 6554
rect 6806 6502 6858 6554
rect 14439 6502 14491 6554
rect 14503 6502 14555 6554
rect 14567 6502 14619 6554
rect 14631 6502 14683 6554
rect 14695 6502 14747 6554
rect 22328 6502 22380 6554
rect 22392 6502 22444 6554
rect 22456 6502 22508 6554
rect 22520 6502 22572 6554
rect 22584 6502 22636 6554
rect 30217 6502 30269 6554
rect 30281 6502 30333 6554
rect 30345 6502 30397 6554
rect 30409 6502 30461 6554
rect 30473 6502 30525 6554
rect 4252 6400 4304 6452
rect 3056 6239 3108 6248
rect 3056 6205 3065 6239
rect 3065 6205 3099 6239
rect 3099 6205 3108 6239
rect 3056 6196 3108 6205
rect 8300 6400 8352 6452
rect 12440 6400 12492 6452
rect 13820 6400 13872 6452
rect 15476 6443 15528 6452
rect 15476 6409 15485 6443
rect 15485 6409 15519 6443
rect 15519 6409 15528 6443
rect 15476 6400 15528 6409
rect 19616 6400 19668 6452
rect 21548 6400 21600 6452
rect 23020 6400 23072 6452
rect 23480 6443 23532 6452
rect 23480 6409 23489 6443
rect 23489 6409 23523 6443
rect 23523 6409 23532 6443
rect 23480 6400 23532 6409
rect 25136 6443 25188 6452
rect 25136 6409 25145 6443
rect 25145 6409 25179 6443
rect 25179 6409 25188 6443
rect 25136 6400 25188 6409
rect 25320 6400 25372 6452
rect 30012 6443 30064 6452
rect 30012 6409 30021 6443
rect 30021 6409 30055 6443
rect 30055 6409 30064 6443
rect 30012 6400 30064 6409
rect 30564 6400 30616 6452
rect 31392 6400 31444 6452
rect 33692 6443 33744 6452
rect 33692 6409 33701 6443
rect 33701 6409 33735 6443
rect 33735 6409 33744 6443
rect 33692 6400 33744 6409
rect 6000 6332 6052 6384
rect 6460 6332 6512 6384
rect 7472 6375 7524 6384
rect 7472 6341 7481 6375
rect 7481 6341 7515 6375
rect 7515 6341 7524 6375
rect 7472 6332 7524 6341
rect 7840 6264 7892 6316
rect 9036 6264 9088 6316
rect 10416 6264 10468 6316
rect 11520 6264 11572 6316
rect 12256 6264 12308 6316
rect 9588 6239 9640 6248
rect 9588 6205 9597 6239
rect 9597 6205 9631 6239
rect 9631 6205 9640 6239
rect 9588 6196 9640 6205
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 13544 6264 13596 6316
rect 16580 6307 16632 6316
rect 16580 6273 16589 6307
rect 16589 6273 16623 6307
rect 16623 6273 16632 6307
rect 16580 6264 16632 6273
rect 16856 6264 16908 6316
rect 7932 6128 7984 6180
rect 10876 6171 10928 6180
rect 10876 6137 10885 6171
rect 10885 6137 10919 6171
rect 10919 6137 10928 6171
rect 10876 6128 10928 6137
rect 12164 6128 12216 6180
rect 4068 6060 4120 6112
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 9772 6060 9824 6112
rect 11796 6060 11848 6112
rect 12808 6171 12860 6180
rect 12808 6137 12817 6171
rect 12817 6137 12851 6171
rect 12851 6137 12860 6171
rect 12808 6128 12860 6137
rect 15660 6196 15712 6248
rect 16948 6239 17000 6248
rect 16948 6205 16957 6239
rect 16957 6205 16991 6239
rect 16991 6205 17000 6239
rect 16948 6196 17000 6205
rect 18696 6196 18748 6248
rect 18972 6196 19024 6248
rect 19432 6264 19484 6316
rect 19800 6307 19852 6316
rect 19800 6273 19809 6307
rect 19809 6273 19843 6307
rect 19843 6273 19852 6307
rect 19800 6264 19852 6273
rect 20260 6264 20312 6316
rect 23848 6264 23900 6316
rect 28816 6307 28868 6316
rect 28816 6273 28824 6307
rect 28824 6273 28858 6307
rect 28858 6273 28868 6307
rect 29184 6332 29236 6384
rect 29460 6332 29512 6384
rect 28816 6264 28868 6273
rect 30564 6264 30616 6316
rect 32036 6264 32088 6316
rect 14188 6128 14240 6180
rect 17960 6128 18012 6180
rect 19892 6239 19944 6248
rect 19892 6205 19901 6239
rect 19901 6205 19935 6239
rect 19935 6205 19944 6239
rect 19892 6196 19944 6205
rect 21732 6128 21784 6180
rect 13360 6060 13412 6112
rect 14464 6060 14516 6112
rect 18788 6060 18840 6112
rect 19616 6103 19668 6112
rect 19616 6069 19625 6103
rect 19625 6069 19659 6103
rect 19659 6069 19668 6103
rect 19616 6060 19668 6069
rect 22192 6060 22244 6112
rect 23572 6196 23624 6248
rect 23664 6239 23716 6248
rect 23664 6205 23673 6239
rect 23673 6205 23707 6239
rect 23707 6205 23716 6239
rect 23664 6196 23716 6205
rect 23756 6239 23808 6248
rect 23756 6205 23765 6239
rect 23765 6205 23799 6239
rect 23799 6205 23808 6239
rect 23756 6196 23808 6205
rect 24032 6239 24084 6248
rect 24032 6205 24041 6239
rect 24041 6205 24075 6239
rect 24075 6205 24084 6239
rect 24032 6196 24084 6205
rect 24308 6239 24360 6248
rect 24308 6205 24317 6239
rect 24317 6205 24351 6239
rect 24351 6205 24360 6239
rect 24308 6196 24360 6205
rect 25228 6239 25280 6248
rect 25228 6205 25237 6239
rect 25237 6205 25271 6239
rect 25271 6205 25280 6239
rect 25228 6196 25280 6205
rect 26424 6239 26476 6248
rect 26424 6205 26433 6239
rect 26433 6205 26467 6239
rect 26467 6205 26476 6239
rect 26424 6196 26476 6205
rect 26884 6196 26936 6248
rect 28448 6239 28500 6248
rect 28448 6205 28457 6239
rect 28457 6205 28491 6239
rect 28491 6205 28500 6239
rect 28448 6196 28500 6205
rect 28724 6239 28776 6248
rect 28724 6205 28732 6239
rect 28732 6205 28766 6239
rect 28766 6205 28776 6239
rect 28724 6196 28776 6205
rect 32588 6196 32640 6248
rect 25780 6128 25832 6180
rect 23388 6060 23440 6112
rect 23664 6060 23716 6112
rect 24492 6060 24544 6112
rect 24952 6103 25004 6112
rect 24952 6069 24961 6103
rect 24961 6069 24995 6103
rect 24995 6069 25004 6103
rect 24952 6060 25004 6069
rect 25688 6060 25740 6112
rect 26976 6128 27028 6180
rect 27252 6060 27304 6112
rect 27712 6103 27764 6112
rect 27712 6069 27721 6103
rect 27721 6069 27755 6103
rect 27755 6069 27764 6103
rect 27712 6060 27764 6069
rect 30656 6128 30708 6180
rect 28908 6060 28960 6112
rect 32312 6103 32364 6112
rect 32312 6069 32321 6103
rect 32321 6069 32355 6103
rect 32355 6069 32364 6103
rect 32312 6060 32364 6069
rect 32864 6103 32916 6112
rect 32864 6069 32873 6103
rect 32873 6069 32907 6103
rect 32907 6069 32916 6103
rect 32864 6060 32916 6069
rect 33784 6060 33836 6112
rect 7210 5958 7262 6010
rect 7274 5958 7326 6010
rect 7338 5958 7390 6010
rect 7402 5958 7454 6010
rect 7466 5958 7518 6010
rect 15099 5958 15151 6010
rect 15163 5958 15215 6010
rect 15227 5958 15279 6010
rect 15291 5958 15343 6010
rect 15355 5958 15407 6010
rect 22988 5958 23040 6010
rect 23052 5958 23104 6010
rect 23116 5958 23168 6010
rect 23180 5958 23232 6010
rect 23244 5958 23296 6010
rect 30877 5958 30929 6010
rect 30941 5958 30993 6010
rect 31005 5958 31057 6010
rect 31069 5958 31121 6010
rect 31133 5958 31185 6010
rect 3148 5856 3200 5908
rect 4252 5856 4304 5908
rect 5264 5856 5316 5908
rect 7104 5856 7156 5908
rect 7932 5856 7984 5908
rect 8392 5856 8444 5908
rect 9312 5856 9364 5908
rect 10048 5856 10100 5908
rect 10876 5856 10928 5908
rect 11704 5856 11756 5908
rect 12164 5899 12216 5908
rect 12164 5865 12173 5899
rect 12173 5865 12207 5899
rect 12207 5865 12216 5899
rect 12164 5856 12216 5865
rect 12808 5856 12860 5908
rect 3240 5788 3292 5840
rect 5080 5720 5132 5772
rect 6460 5788 6512 5840
rect 7656 5720 7708 5772
rect 8208 5788 8260 5840
rect 10784 5720 10836 5772
rect 11796 5831 11848 5840
rect 11796 5797 11805 5831
rect 11805 5797 11839 5831
rect 11839 5797 11848 5831
rect 11796 5788 11848 5797
rect 13360 5788 13412 5840
rect 16948 5856 17000 5908
rect 17960 5899 18012 5908
rect 17960 5865 17969 5899
rect 17969 5865 18003 5899
rect 18003 5865 18012 5899
rect 17960 5856 18012 5865
rect 20260 5856 20312 5908
rect 11612 5763 11664 5772
rect 11612 5729 11621 5763
rect 11621 5729 11655 5763
rect 11655 5729 11664 5763
rect 11612 5720 11664 5729
rect 4896 5652 4948 5704
rect 6920 5652 6972 5704
rect 8576 5695 8628 5704
rect 8576 5661 8585 5695
rect 8585 5661 8619 5695
rect 8619 5661 8628 5695
rect 8576 5652 8628 5661
rect 8668 5652 8720 5704
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 4988 5516 5040 5568
rect 7288 5559 7340 5568
rect 7288 5525 7297 5559
rect 7297 5525 7331 5559
rect 7331 5525 7340 5559
rect 7288 5516 7340 5525
rect 10048 5516 10100 5568
rect 11980 5763 12032 5772
rect 11980 5729 11989 5763
rect 11989 5729 12023 5763
rect 12023 5729 12032 5763
rect 11980 5720 12032 5729
rect 12072 5720 12124 5772
rect 14096 5720 14148 5772
rect 14464 5720 14516 5772
rect 21916 5856 21968 5908
rect 25504 5856 25556 5908
rect 27252 5856 27304 5908
rect 27988 5856 28040 5908
rect 23664 5788 23716 5840
rect 25320 5788 25372 5840
rect 29276 5856 29328 5908
rect 30564 5856 30616 5908
rect 30656 5856 30708 5908
rect 31760 5856 31812 5908
rect 16764 5720 16816 5772
rect 17868 5763 17920 5772
rect 17868 5729 17877 5763
rect 17877 5729 17911 5763
rect 17911 5729 17920 5763
rect 17868 5720 17920 5729
rect 22192 5720 22244 5772
rect 24216 5763 24268 5772
rect 24216 5729 24225 5763
rect 24225 5729 24259 5763
rect 24259 5729 24268 5763
rect 24216 5720 24268 5729
rect 11888 5652 11940 5704
rect 12164 5652 12216 5704
rect 12348 5695 12400 5704
rect 12348 5661 12357 5695
rect 12357 5661 12391 5695
rect 12391 5661 12400 5695
rect 12348 5652 12400 5661
rect 12256 5584 12308 5636
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 13728 5516 13780 5568
rect 16396 5516 16448 5568
rect 18328 5652 18380 5704
rect 19064 5695 19116 5704
rect 19064 5661 19073 5695
rect 19073 5661 19107 5695
rect 19107 5661 19116 5695
rect 19064 5652 19116 5661
rect 19340 5695 19392 5704
rect 19340 5661 19349 5695
rect 19349 5661 19383 5695
rect 19383 5661 19392 5695
rect 19340 5652 19392 5661
rect 24308 5652 24360 5704
rect 24492 5695 24544 5704
rect 24492 5661 24501 5695
rect 24501 5661 24535 5695
rect 24535 5661 24544 5695
rect 24492 5652 24544 5661
rect 24860 5652 24912 5704
rect 25228 5695 25280 5704
rect 25228 5661 25237 5695
rect 25237 5661 25271 5695
rect 25271 5661 25280 5695
rect 25228 5652 25280 5661
rect 25412 5695 25464 5704
rect 25412 5661 25421 5695
rect 25421 5661 25455 5695
rect 25455 5661 25464 5695
rect 25412 5652 25464 5661
rect 25688 5695 25740 5704
rect 25688 5661 25697 5695
rect 25697 5661 25731 5695
rect 25731 5661 25740 5695
rect 25688 5652 25740 5661
rect 26700 5763 26752 5772
rect 26700 5729 26709 5763
rect 26709 5729 26743 5763
rect 26743 5729 26752 5763
rect 26700 5720 26752 5729
rect 27436 5720 27488 5772
rect 29184 5788 29236 5840
rect 31944 5788 31996 5840
rect 32864 5856 32916 5908
rect 30012 5720 30064 5772
rect 30840 5720 30892 5772
rect 33784 5763 33836 5772
rect 33784 5729 33793 5763
rect 33793 5729 33827 5763
rect 33827 5729 33836 5763
rect 33784 5720 33836 5729
rect 22652 5584 22704 5636
rect 16580 5559 16632 5568
rect 16580 5525 16589 5559
rect 16589 5525 16623 5559
rect 16623 5525 16632 5559
rect 16580 5516 16632 5525
rect 18696 5559 18748 5568
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 20812 5559 20864 5568
rect 20812 5525 20821 5559
rect 20821 5525 20855 5559
rect 20855 5525 20864 5559
rect 20812 5516 20864 5525
rect 27620 5584 27672 5636
rect 27804 5695 27856 5704
rect 27804 5661 27813 5695
rect 27813 5661 27847 5695
rect 27847 5661 27856 5695
rect 27804 5652 27856 5661
rect 28172 5652 28224 5704
rect 29368 5652 29420 5704
rect 29552 5652 29604 5704
rect 31484 5695 31536 5704
rect 31484 5661 31493 5695
rect 31493 5661 31527 5695
rect 31527 5661 31536 5695
rect 31484 5652 31536 5661
rect 33140 5584 33192 5636
rect 27528 5559 27580 5568
rect 27528 5525 27537 5559
rect 27537 5525 27571 5559
rect 27571 5525 27580 5559
rect 27528 5516 27580 5525
rect 32404 5516 32456 5568
rect 6550 5414 6602 5466
rect 6614 5414 6666 5466
rect 6678 5414 6730 5466
rect 6742 5414 6794 5466
rect 6806 5414 6858 5466
rect 14439 5414 14491 5466
rect 14503 5414 14555 5466
rect 14567 5414 14619 5466
rect 14631 5414 14683 5466
rect 14695 5414 14747 5466
rect 22328 5414 22380 5466
rect 22392 5414 22444 5466
rect 22456 5414 22508 5466
rect 22520 5414 22572 5466
rect 22584 5414 22636 5466
rect 30217 5414 30269 5466
rect 30281 5414 30333 5466
rect 30345 5414 30397 5466
rect 30409 5414 30461 5466
rect 30473 5414 30525 5466
rect 8576 5312 8628 5364
rect 9772 5312 9824 5364
rect 4160 5176 4212 5228
rect 4988 5219 5040 5228
rect 4988 5185 4997 5219
rect 4997 5185 5031 5219
rect 5031 5185 5040 5219
rect 4988 5176 5040 5185
rect 5540 5176 5592 5228
rect 7840 5176 7892 5228
rect 7932 5176 7984 5228
rect 8300 5176 8352 5228
rect 8484 5176 8536 5228
rect 10140 5176 10192 5228
rect 11520 5312 11572 5364
rect 11888 5312 11940 5364
rect 14096 5355 14148 5364
rect 14096 5321 14105 5355
rect 14105 5321 14139 5355
rect 14139 5321 14148 5355
rect 14096 5312 14148 5321
rect 14188 5312 14240 5364
rect 15016 5312 15068 5364
rect 15660 5312 15712 5364
rect 16028 5312 16080 5364
rect 18604 5312 18656 5364
rect 19340 5312 19392 5364
rect 19800 5312 19852 5364
rect 21732 5355 21784 5364
rect 21732 5321 21741 5355
rect 21741 5321 21775 5355
rect 21775 5321 21784 5355
rect 21732 5312 21784 5321
rect 23572 5312 23624 5364
rect 23756 5312 23808 5364
rect 24216 5312 24268 5364
rect 27804 5312 27856 5364
rect 30012 5312 30064 5364
rect 26608 5244 26660 5296
rect 28908 5244 28960 5296
rect 31208 5244 31260 5296
rect 12348 5176 12400 5228
rect 13728 5176 13780 5228
rect 16304 5176 16356 5228
rect 16580 5176 16632 5228
rect 16856 5219 16908 5228
rect 16856 5185 16865 5219
rect 16865 5185 16899 5219
rect 16899 5185 16908 5219
rect 16856 5176 16908 5185
rect 7288 5108 7340 5160
rect 7656 5151 7708 5160
rect 7656 5117 7665 5151
rect 7665 5117 7699 5151
rect 7699 5117 7708 5151
rect 7656 5108 7708 5117
rect 3240 5083 3292 5092
rect 3240 5049 3249 5083
rect 3249 5049 3283 5083
rect 3283 5049 3292 5083
rect 3240 5040 3292 5049
rect 4528 5015 4580 5024
rect 4528 4981 4537 5015
rect 4537 4981 4571 5015
rect 4571 4981 4580 5015
rect 4528 4972 4580 4981
rect 5264 4972 5316 5024
rect 6460 5040 6512 5092
rect 8852 5108 8904 5160
rect 13268 5108 13320 5160
rect 14832 5108 14884 5160
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 8392 5040 8444 5092
rect 8576 5083 8628 5092
rect 8576 5049 8585 5083
rect 8585 5049 8619 5083
rect 8619 5049 8628 5083
rect 8576 5040 8628 5049
rect 5908 4972 5960 5024
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 8668 5015 8720 5024
rect 8668 4981 8677 5015
rect 8677 4981 8711 5015
rect 8711 4981 8720 5015
rect 8668 4972 8720 4981
rect 9680 5040 9732 5092
rect 10048 5040 10100 5092
rect 19156 5176 19208 5228
rect 19524 5176 19576 5228
rect 19616 5176 19668 5228
rect 20812 5176 20864 5228
rect 22836 5176 22888 5228
rect 18972 5108 19024 5160
rect 20352 5108 20404 5160
rect 23388 5108 23440 5160
rect 24952 5176 25004 5228
rect 25964 5176 26016 5228
rect 26700 5176 26752 5228
rect 27712 5176 27764 5228
rect 28448 5219 28500 5228
rect 28448 5185 28457 5219
rect 28457 5185 28491 5219
rect 28491 5185 28500 5219
rect 28448 5176 28500 5185
rect 29184 5176 29236 5228
rect 30748 5176 30800 5228
rect 31760 5219 31812 5228
rect 31760 5185 31769 5219
rect 31769 5185 31803 5219
rect 31803 5185 31812 5219
rect 31760 5176 31812 5185
rect 28632 5108 28684 5160
rect 29828 5151 29880 5160
rect 29828 5117 29837 5151
rect 29837 5117 29871 5151
rect 29871 5117 29880 5151
rect 29828 5108 29880 5117
rect 30012 5108 30064 5160
rect 34888 5176 34940 5228
rect 20076 5040 20128 5092
rect 13268 5015 13320 5024
rect 13268 4981 13277 5015
rect 13277 4981 13311 5015
rect 13311 4981 13320 5015
rect 13268 4972 13320 4981
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 17960 4972 18012 5024
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 23848 4972 23900 5024
rect 25412 5015 25464 5024
rect 25412 4981 25421 5015
rect 25421 4981 25455 5015
rect 25455 4981 25464 5015
rect 25412 4972 25464 4981
rect 27528 5040 27580 5092
rect 33140 5040 33192 5092
rect 28540 5015 28592 5024
rect 28540 4981 28549 5015
rect 28549 4981 28583 5015
rect 28583 4981 28592 5015
rect 28540 4972 28592 4981
rect 29092 4972 29144 5024
rect 31208 5015 31260 5024
rect 31208 4981 31217 5015
rect 31217 4981 31251 5015
rect 31251 4981 31260 5015
rect 31208 4972 31260 4981
rect 32036 5015 32088 5024
rect 32036 4981 32045 5015
rect 32045 4981 32079 5015
rect 32079 4981 32088 5015
rect 32036 4972 32088 4981
rect 32220 4972 32272 5024
rect 7210 4870 7262 4922
rect 7274 4870 7326 4922
rect 7338 4870 7390 4922
rect 7402 4870 7454 4922
rect 7466 4870 7518 4922
rect 15099 4870 15151 4922
rect 15163 4870 15215 4922
rect 15227 4870 15279 4922
rect 15291 4870 15343 4922
rect 15355 4870 15407 4922
rect 22988 4870 23040 4922
rect 23052 4870 23104 4922
rect 23116 4870 23168 4922
rect 23180 4870 23232 4922
rect 23244 4870 23296 4922
rect 30877 4870 30929 4922
rect 30941 4870 30993 4922
rect 31005 4870 31057 4922
rect 31069 4870 31121 4922
rect 31133 4870 31185 4922
rect 4896 4768 4948 4820
rect 5356 4768 5408 4820
rect 5448 4811 5500 4820
rect 5448 4777 5457 4811
rect 5457 4777 5491 4811
rect 5491 4777 5500 4811
rect 5448 4768 5500 4777
rect 1308 4632 1360 4684
rect 5908 4700 5960 4752
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 5816 4675 5868 4684
rect 5816 4641 5825 4675
rect 5825 4641 5859 4675
rect 5859 4641 5868 4675
rect 5816 4632 5868 4641
rect 6276 4768 6328 4820
rect 6368 4768 6420 4820
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 6092 4700 6144 4752
rect 7748 4700 7800 4752
rect 9680 4768 9732 4820
rect 11796 4768 11848 4820
rect 12256 4811 12308 4820
rect 12256 4777 12265 4811
rect 12265 4777 12299 4811
rect 12299 4777 12308 4811
rect 12256 4768 12308 4777
rect 15936 4768 15988 4820
rect 15292 4700 15344 4752
rect 4804 4607 4856 4616
rect 4804 4573 4813 4607
rect 4813 4573 4847 4607
rect 4847 4573 4856 4607
rect 4804 4564 4856 4573
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 5264 4564 5316 4616
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 10140 4632 10192 4684
rect 10784 4675 10836 4684
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 11796 4632 11848 4684
rect 16948 4768 17000 4820
rect 17868 4768 17920 4820
rect 16304 4743 16356 4752
rect 16304 4709 16313 4743
rect 16313 4709 16347 4743
rect 16347 4709 16356 4743
rect 16304 4700 16356 4709
rect 20076 4811 20128 4820
rect 20076 4777 20085 4811
rect 20085 4777 20119 4811
rect 20119 4777 20128 4811
rect 20076 4768 20128 4777
rect 23388 4768 23440 4820
rect 19156 4700 19208 4752
rect 18328 4675 18380 4684
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 6368 4564 6420 4573
rect 7932 4496 7984 4548
rect 8392 4496 8444 4548
rect 8300 4428 8352 4480
rect 9496 4607 9548 4616
rect 9496 4573 9505 4607
rect 9505 4573 9539 4607
rect 9539 4573 9548 4607
rect 9496 4564 9548 4573
rect 11888 4564 11940 4616
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 16764 4564 16816 4616
rect 18604 4607 18656 4616
rect 18604 4573 18613 4607
rect 18613 4573 18647 4607
rect 18647 4573 18656 4607
rect 18604 4564 18656 4573
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 24768 4768 24820 4820
rect 23848 4632 23900 4684
rect 25412 4768 25464 4820
rect 28172 4811 28224 4820
rect 28172 4777 28181 4811
rect 28181 4777 28215 4811
rect 28215 4777 28224 4811
rect 28172 4768 28224 4777
rect 28632 4811 28684 4820
rect 28632 4777 28641 4811
rect 28641 4777 28675 4811
rect 28675 4777 28684 4811
rect 28632 4768 28684 4777
rect 29000 4811 29052 4820
rect 29000 4777 29009 4811
rect 29009 4777 29043 4811
rect 29043 4777 29052 4811
rect 29000 4768 29052 4777
rect 29092 4811 29144 4820
rect 29092 4777 29101 4811
rect 29101 4777 29135 4811
rect 29135 4777 29144 4811
rect 29092 4768 29144 4777
rect 26884 4700 26936 4752
rect 24952 4607 25004 4616
rect 24952 4573 24961 4607
rect 24961 4573 24995 4607
rect 24995 4573 25004 4607
rect 24952 4564 25004 4573
rect 25596 4607 25648 4616
rect 25596 4573 25605 4607
rect 25605 4573 25639 4607
rect 25639 4573 25648 4607
rect 25596 4564 25648 4573
rect 25964 4564 26016 4616
rect 29552 4700 29604 4752
rect 31208 4768 31260 4820
rect 31944 4768 31996 4820
rect 32036 4700 32088 4752
rect 27436 4632 27488 4684
rect 30012 4632 30064 4684
rect 32220 4675 32272 4684
rect 32220 4641 32229 4675
rect 32229 4641 32263 4675
rect 32263 4641 32272 4675
rect 32220 4632 32272 4641
rect 28908 4564 28960 4616
rect 30748 4564 30800 4616
rect 34704 4564 34756 4616
rect 28724 4496 28776 4548
rect 15200 4471 15252 4480
rect 15200 4437 15209 4471
rect 15209 4437 15243 4471
rect 15243 4437 15252 4471
rect 15200 4428 15252 4437
rect 17960 4428 18012 4480
rect 19340 4428 19392 4480
rect 21180 4428 21232 4480
rect 23664 4428 23716 4480
rect 27068 4471 27120 4480
rect 27068 4437 27077 4471
rect 27077 4437 27111 4471
rect 27111 4437 27120 4471
rect 27068 4428 27120 4437
rect 29552 4471 29604 4480
rect 29552 4437 29561 4471
rect 29561 4437 29595 4471
rect 29595 4437 29604 4471
rect 29552 4428 29604 4437
rect 6550 4326 6602 4378
rect 6614 4326 6666 4378
rect 6678 4326 6730 4378
rect 6742 4326 6794 4378
rect 6806 4326 6858 4378
rect 14439 4326 14491 4378
rect 14503 4326 14555 4378
rect 14567 4326 14619 4378
rect 14631 4326 14683 4378
rect 14695 4326 14747 4378
rect 22328 4326 22380 4378
rect 22392 4326 22444 4378
rect 22456 4326 22508 4378
rect 22520 4326 22572 4378
rect 22584 4326 22636 4378
rect 30217 4326 30269 4378
rect 30281 4326 30333 4378
rect 30345 4326 30397 4378
rect 30409 4326 30461 4378
rect 30473 4326 30525 4378
rect 4804 4224 4856 4276
rect 5540 4224 5592 4276
rect 6092 4267 6144 4276
rect 6092 4233 6101 4267
rect 6101 4233 6135 4267
rect 6135 4233 6144 4267
rect 6092 4224 6144 4233
rect 6276 4224 6328 4276
rect 8484 4224 8536 4276
rect 9496 4224 9548 4276
rect 13636 4224 13688 4276
rect 15292 4267 15344 4276
rect 15292 4233 15301 4267
rect 15301 4233 15335 4267
rect 15335 4233 15344 4267
rect 15292 4224 15344 4233
rect 16856 4224 16908 4276
rect 18604 4224 18656 4276
rect 24952 4224 25004 4276
rect 25596 4224 25648 4276
rect 26884 4267 26936 4276
rect 26884 4233 26893 4267
rect 26893 4233 26927 4267
rect 26927 4233 26936 4267
rect 26884 4224 26936 4233
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 5632 4156 5684 4208
rect 6368 4088 6420 4140
rect 4436 4063 4488 4072
rect 4436 4029 4445 4063
rect 4445 4029 4479 4063
rect 4479 4029 4488 4063
rect 4436 4020 4488 4029
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 20 3952 72 4004
rect 8576 4020 8628 4072
rect 9036 4088 9088 4140
rect 12532 4088 12584 4140
rect 13728 4088 13780 4140
rect 14648 4088 14700 4140
rect 15200 4088 15252 4140
rect 18696 4088 18748 4140
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 21180 4131 21232 4140
rect 21180 4097 21189 4131
rect 21189 4097 21223 4131
rect 21223 4097 21232 4131
rect 21180 4088 21232 4097
rect 14004 4020 14056 4072
rect 14832 3952 14884 4004
rect 18236 4020 18288 4072
rect 21732 4020 21784 4072
rect 23756 4063 23808 4072
rect 23756 4029 23765 4063
rect 23765 4029 23799 4063
rect 23799 4029 23808 4063
rect 23756 4020 23808 4029
rect 22836 3884 22888 3936
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 25504 4131 25556 4140
rect 25504 4097 25513 4131
rect 25513 4097 25547 4131
rect 25547 4097 25556 4131
rect 25504 4088 25556 4097
rect 26608 4131 26660 4140
rect 26608 4097 26617 4131
rect 26617 4097 26651 4131
rect 26651 4097 26660 4131
rect 26608 4088 26660 4097
rect 28448 4224 28500 4276
rect 29828 4224 29880 4276
rect 28540 4088 28592 4140
rect 28724 4088 28776 4140
rect 27436 4020 27488 4072
rect 29552 4020 29604 4072
rect 28908 3884 28960 3936
rect 29000 3884 29052 3936
rect 33968 4063 34020 4072
rect 33968 4029 33977 4063
rect 33977 4029 34011 4063
rect 34011 4029 34020 4063
rect 33968 4020 34020 4029
rect 34428 4020 34480 4072
rect 7210 3782 7262 3834
rect 7274 3782 7326 3834
rect 7338 3782 7390 3834
rect 7402 3782 7454 3834
rect 7466 3782 7518 3834
rect 15099 3782 15151 3834
rect 15163 3782 15215 3834
rect 15227 3782 15279 3834
rect 15291 3782 15343 3834
rect 15355 3782 15407 3834
rect 22988 3782 23040 3834
rect 23052 3782 23104 3834
rect 23116 3782 23168 3834
rect 23180 3782 23232 3834
rect 23244 3782 23296 3834
rect 30877 3782 30929 3834
rect 30941 3782 30993 3834
rect 31005 3782 31057 3834
rect 31069 3782 31121 3834
rect 31133 3782 31185 3834
rect 9036 3723 9088 3732
rect 9036 3689 9045 3723
rect 9045 3689 9079 3723
rect 9079 3689 9088 3723
rect 9036 3680 9088 3689
rect 14648 3723 14700 3732
rect 14648 3689 14657 3723
rect 14657 3689 14691 3723
rect 14691 3689 14700 3723
rect 14648 3680 14700 3689
rect 25872 3680 25924 3732
rect 25964 3723 26016 3732
rect 25964 3689 25973 3723
rect 25973 3689 26007 3723
rect 26007 3689 26016 3723
rect 25964 3680 26016 3689
rect 26792 3680 26844 3732
rect 28724 3680 28776 3732
rect 28908 3723 28960 3732
rect 28908 3689 28917 3723
rect 28917 3689 28951 3723
rect 28951 3689 28960 3723
rect 28908 3680 28960 3689
rect 1308 3612 1360 3664
rect 3240 3612 3292 3664
rect 29000 3612 29052 3664
rect 4896 3544 4948 3596
rect 8668 3544 8720 3596
rect 16396 3587 16448 3596
rect 16396 3553 16405 3587
rect 16405 3553 16439 3587
rect 16439 3553 16448 3587
rect 16396 3544 16448 3553
rect 19340 3544 19392 3596
rect 32312 3587 32364 3596
rect 32312 3553 32321 3587
rect 32321 3553 32355 3587
rect 32355 3553 32364 3587
rect 32312 3544 32364 3553
rect 35440 3544 35492 3596
rect 1308 3476 1360 3528
rect 5172 3476 5224 3528
rect 16120 3476 16172 3528
rect 20628 3476 20680 3528
rect 21824 3476 21876 3528
rect 33048 3519 33100 3528
rect 33048 3485 33057 3519
rect 33057 3485 33091 3519
rect 33091 3485 33100 3519
rect 33048 3476 33100 3485
rect 13636 3408 13688 3460
rect 24400 3408 24452 3460
rect 9680 3340 9732 3392
rect 18512 3340 18564 3392
rect 6550 3238 6602 3290
rect 6614 3238 6666 3290
rect 6678 3238 6730 3290
rect 6742 3238 6794 3290
rect 6806 3238 6858 3290
rect 14439 3238 14491 3290
rect 14503 3238 14555 3290
rect 14567 3238 14619 3290
rect 14631 3238 14683 3290
rect 14695 3238 14747 3290
rect 22328 3238 22380 3290
rect 22392 3238 22444 3290
rect 22456 3238 22508 3290
rect 22520 3238 22572 3290
rect 22584 3238 22636 3290
rect 30217 3238 30269 3290
rect 30281 3238 30333 3290
rect 30345 3238 30397 3290
rect 30409 3238 30461 3290
rect 30473 3238 30525 3290
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 13636 3136 13688 3188
rect 24492 3136 24544 3188
rect 25228 3136 25280 3188
rect 27620 3136 27672 3188
rect 31576 3136 31628 3188
rect 2596 3000 2648 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 7748 3000 7800 3052
rect 3056 2975 3108 2984
rect 3056 2941 3065 2975
rect 3065 2941 3099 2975
rect 3099 2941 3108 2975
rect 3056 2932 3108 2941
rect 5264 2975 5316 2984
rect 5264 2941 5273 2975
rect 5273 2941 5307 2975
rect 5307 2941 5316 2975
rect 5264 2932 5316 2941
rect 4068 2907 4120 2916
rect 4068 2873 4077 2907
rect 4077 2873 4111 2907
rect 4111 2873 4120 2907
rect 4068 2864 4120 2873
rect 6644 2907 6696 2916
rect 6644 2873 6653 2907
rect 6653 2873 6687 2907
rect 6687 2873 6696 2907
rect 6644 2864 6696 2873
rect 8024 2975 8076 2984
rect 8024 2941 8033 2975
rect 8033 2941 8067 2975
rect 8067 2941 8076 2975
rect 8024 2932 8076 2941
rect 9036 2932 9088 2984
rect 9128 2864 9180 2916
rect 24308 3068 24360 3120
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 17408 3043 17460 3052
rect 17408 3009 17417 3043
rect 17417 3009 17451 3043
rect 17451 3009 17460 3043
rect 17408 3000 17460 3009
rect 18696 3000 18748 3052
rect 22008 3000 22060 3052
rect 24584 3000 24636 3052
rect 27160 3000 27212 3052
rect 29736 3000 29788 3052
rect 32864 3043 32916 3052
rect 32864 3009 32873 3043
rect 32873 3009 32907 3043
rect 32907 3009 32916 3043
rect 32864 3000 32916 3009
rect 10968 2932 11020 2984
rect 13268 2932 13320 2984
rect 13636 2975 13688 2984
rect 13636 2941 13645 2975
rect 13645 2941 13679 2975
rect 13679 2941 13688 2975
rect 13636 2932 13688 2941
rect 13912 2932 13964 2984
rect 16764 2975 16816 2984
rect 16764 2941 16773 2975
rect 16773 2941 16807 2975
rect 16807 2941 16816 2975
rect 16764 2932 16816 2941
rect 18788 2975 18840 2984
rect 18788 2941 18797 2975
rect 18797 2941 18831 2975
rect 18831 2941 18840 2975
rect 18788 2932 18840 2941
rect 21180 2932 21232 2984
rect 23388 2932 23440 2984
rect 23664 2932 23716 2984
rect 25780 2932 25832 2984
rect 27068 2975 27120 2984
rect 27068 2941 27077 2975
rect 27077 2941 27111 2975
rect 27111 2941 27120 2975
rect 27068 2932 27120 2941
rect 28356 2932 28408 2984
rect 29828 2975 29880 2984
rect 29828 2941 29837 2975
rect 29837 2941 29871 2975
rect 29871 2941 29880 2975
rect 29828 2932 29880 2941
rect 31576 2932 31628 2984
rect 31944 2932 31996 2984
rect 36728 2932 36780 2984
rect 21088 2864 21140 2916
rect 25688 2796 25740 2848
rect 7210 2694 7262 2746
rect 7274 2694 7326 2746
rect 7338 2694 7390 2746
rect 7402 2694 7454 2746
rect 7466 2694 7518 2746
rect 15099 2694 15151 2746
rect 15163 2694 15215 2746
rect 15227 2694 15279 2746
rect 15291 2694 15343 2746
rect 15355 2694 15407 2746
rect 22988 2694 23040 2746
rect 23052 2694 23104 2746
rect 23116 2694 23168 2746
rect 23180 2694 23232 2746
rect 23244 2694 23296 2746
rect 30877 2694 30929 2746
rect 30941 2694 30993 2746
rect 31005 2694 31057 2746
rect 31069 2694 31121 2746
rect 31133 2694 31185 2746
<< metal2 >>
rect 662 35678 718 36478
rect 1950 35678 2006 36478
rect 3238 35678 3294 36478
rect 3790 36136 3846 36145
rect 3790 36071 3846 36080
rect 676 32434 704 35678
rect 1964 33114 1992 35678
rect 3054 34776 3110 34785
rect 3054 34711 3110 34720
rect 3068 34066 3096 34711
rect 3056 34060 3108 34066
rect 3056 34002 3108 34008
rect 3252 33522 3280 35678
rect 3240 33516 3292 33522
rect 3240 33458 3292 33464
rect 3238 33416 3294 33425
rect 3238 33351 3294 33360
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 3252 33046 3280 33351
rect 3804 33046 3832 36071
rect 4526 35678 4582 36478
rect 5814 35678 5870 36478
rect 7746 35678 7802 36478
rect 9034 35678 9090 36478
rect 10322 35678 10378 36478
rect 11610 35678 11666 36478
rect 12898 35678 12954 36478
rect 14186 35678 14242 36478
rect 15474 35678 15530 36478
rect 17406 35678 17462 36478
rect 18694 35678 18750 36478
rect 19982 35678 20038 36478
rect 21270 35678 21326 36478
rect 22558 35678 22614 36478
rect 23846 35678 23902 36478
rect 25134 35678 25190 36478
rect 26422 35678 26478 36478
rect 28354 35678 28410 36478
rect 29642 35678 29698 36478
rect 30930 35678 30986 36478
rect 31036 35686 31340 35714
rect 4540 34134 4568 35678
rect 5828 34134 5856 35678
rect 7210 34300 7518 34309
rect 7210 34298 7216 34300
rect 7272 34298 7296 34300
rect 7352 34298 7376 34300
rect 7432 34298 7456 34300
rect 7512 34298 7518 34300
rect 7272 34246 7274 34298
rect 7454 34246 7456 34298
rect 7210 34244 7216 34246
rect 7272 34244 7296 34246
rect 7352 34244 7376 34246
rect 7432 34244 7456 34246
rect 7512 34244 7518 34246
rect 7210 34235 7518 34244
rect 7760 34202 7788 35678
rect 7748 34196 7800 34202
rect 7748 34138 7800 34144
rect 4528 34128 4580 34134
rect 4528 34070 4580 34076
rect 5816 34128 5868 34134
rect 5816 34070 5868 34076
rect 4712 34060 4764 34066
rect 4712 34002 4764 34008
rect 6000 34060 6052 34066
rect 9048 34048 9076 35678
rect 10336 34066 10364 35678
rect 9128 34060 9180 34066
rect 9048 34020 9128 34048
rect 6000 34002 6052 34008
rect 9128 34002 9180 34008
rect 10324 34060 10376 34066
rect 10324 34002 10376 34008
rect 3240 33040 3292 33046
rect 3240 32982 3292 32988
rect 3792 33040 3844 33046
rect 3792 32982 3844 32988
rect 664 32428 716 32434
rect 664 32370 716 32376
rect 4436 32360 4488 32366
rect 4434 32328 4436 32337
rect 4488 32328 4490 32337
rect 4434 32263 4490 32272
rect 4620 31884 4672 31890
rect 4620 31826 4672 31832
rect 3240 31816 3292 31822
rect 3240 31758 3292 31764
rect 3252 31385 3280 31758
rect 4632 31754 4660 31826
rect 4540 31726 4660 31754
rect 3238 31376 3294 31385
rect 3238 31311 3294 31320
rect 3332 31204 3384 31210
rect 3332 31146 3384 31152
rect 3344 30394 3372 31146
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 3332 30388 3384 30394
rect 3332 30330 3384 30336
rect 4172 30190 4200 30534
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 1308 30116 1360 30122
rect 1308 30058 1360 30064
rect 1320 30025 1348 30058
rect 3240 30048 3292 30054
rect 1306 30016 1362 30025
rect 3240 29990 3292 29996
rect 1306 29951 1362 29960
rect 1306 28656 1362 28665
rect 1306 28591 1308 28600
rect 1360 28591 1362 28600
rect 1308 28562 1360 28568
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 1320 26926 1348 27231
rect 1308 26920 1360 26926
rect 1308 26862 1360 26868
rect 3252 26466 3280 29990
rect 4540 29306 4568 31726
rect 4724 30954 4752 34002
rect 5540 33856 5592 33862
rect 5540 33798 5592 33804
rect 5448 33448 5500 33454
rect 5448 33390 5500 33396
rect 5172 33312 5224 33318
rect 5172 33254 5224 33260
rect 5080 32224 5132 32230
rect 5080 32166 5132 32172
rect 5092 31958 5120 32166
rect 5080 31952 5132 31958
rect 5080 31894 5132 31900
rect 4896 31884 4948 31890
rect 4896 31826 4948 31832
rect 4908 31346 4936 31826
rect 5080 31408 5132 31414
rect 5080 31350 5132 31356
rect 4896 31340 4948 31346
rect 4896 31282 4948 31288
rect 4896 31136 4948 31142
rect 4896 31078 4948 31084
rect 4632 30926 4752 30954
rect 4908 30938 4936 31078
rect 4896 30932 4948 30938
rect 4528 29300 4580 29306
rect 4528 29242 4580 29248
rect 4436 28620 4488 28626
rect 4436 28562 4488 28568
rect 3976 28008 4028 28014
rect 3976 27950 4028 27956
rect 3988 27130 4016 27950
rect 4448 27334 4476 28562
rect 4528 27872 4580 27878
rect 4528 27814 4580 27820
rect 4540 27606 4568 27814
rect 4528 27600 4580 27606
rect 4528 27542 4580 27548
rect 4436 27328 4488 27334
rect 4436 27270 4488 27276
rect 3976 27124 4028 27130
rect 3976 27066 4028 27072
rect 4448 26994 4476 27270
rect 4632 26994 4660 30926
rect 4896 30874 4948 30880
rect 4712 30864 4764 30870
rect 4712 30806 4764 30812
rect 4724 29714 4752 30806
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 4988 29572 5040 29578
rect 4988 29514 5040 29520
rect 5000 29102 5028 29514
rect 4988 29096 5040 29102
rect 4988 29038 5040 29044
rect 5000 27520 5028 29038
rect 5092 28914 5120 31350
rect 5184 29102 5212 33254
rect 5356 32836 5408 32842
rect 5356 32778 5408 32784
rect 5368 30870 5396 32778
rect 5460 31482 5488 33390
rect 5448 31476 5500 31482
rect 5448 31418 5500 31424
rect 5356 30864 5408 30870
rect 5356 30806 5408 30812
rect 5264 30728 5316 30734
rect 5264 30670 5316 30676
rect 5276 30394 5304 30670
rect 5264 30388 5316 30394
rect 5264 30330 5316 30336
rect 5460 30258 5488 31418
rect 5552 31278 5580 33798
rect 5908 33516 5960 33522
rect 5908 33458 5960 33464
rect 5920 33114 5948 33458
rect 5908 33108 5960 33114
rect 5908 33050 5960 33056
rect 5724 32972 5776 32978
rect 5724 32914 5776 32920
rect 5736 31754 5764 32914
rect 6012 32434 6040 34002
rect 9220 33992 9272 33998
rect 9220 33934 9272 33940
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 8208 33856 8260 33862
rect 8208 33798 8260 33804
rect 6550 33756 6858 33765
rect 6550 33754 6556 33756
rect 6612 33754 6636 33756
rect 6692 33754 6716 33756
rect 6772 33754 6796 33756
rect 6852 33754 6858 33756
rect 6612 33702 6614 33754
rect 6794 33702 6796 33754
rect 6550 33700 6556 33702
rect 6612 33700 6636 33702
rect 6692 33700 6716 33702
rect 6772 33700 6796 33702
rect 6852 33700 6858 33702
rect 6550 33691 6858 33700
rect 7932 33448 7984 33454
rect 7932 33390 7984 33396
rect 7210 33212 7518 33221
rect 7210 33210 7216 33212
rect 7272 33210 7296 33212
rect 7352 33210 7376 33212
rect 7432 33210 7456 33212
rect 7512 33210 7518 33212
rect 7272 33158 7274 33210
rect 7454 33158 7456 33210
rect 7210 33156 7216 33158
rect 7272 33156 7296 33158
rect 7352 33156 7376 33158
rect 7432 33156 7456 33158
rect 7512 33156 7518 33158
rect 7210 33147 7518 33156
rect 7288 32972 7340 32978
rect 7288 32914 7340 32920
rect 7300 32774 7328 32914
rect 7288 32768 7340 32774
rect 7288 32710 7340 32716
rect 6550 32668 6858 32677
rect 6550 32666 6556 32668
rect 6612 32666 6636 32668
rect 6692 32666 6716 32668
rect 6772 32666 6796 32668
rect 6852 32666 6858 32668
rect 6612 32614 6614 32666
rect 6794 32614 6796 32666
rect 6550 32612 6556 32614
rect 6612 32612 6636 32614
rect 6692 32612 6716 32614
rect 6772 32612 6796 32614
rect 6852 32612 6858 32614
rect 6550 32603 6858 32612
rect 7300 32502 7328 32710
rect 7288 32496 7340 32502
rect 7024 32444 7288 32450
rect 7024 32438 7340 32444
rect 6000 32428 6052 32434
rect 6000 32370 6052 32376
rect 6460 32428 6512 32434
rect 6460 32370 6512 32376
rect 7024 32422 7328 32438
rect 5908 32224 5960 32230
rect 5908 32166 5960 32172
rect 5644 31726 5764 31754
rect 5540 31272 5592 31278
rect 5540 31214 5592 31220
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 5644 29646 5672 31726
rect 5816 30592 5868 30598
rect 5816 30534 5868 30540
rect 5724 30116 5776 30122
rect 5724 30058 5776 30064
rect 5736 29850 5764 30058
rect 5828 29850 5856 30534
rect 5724 29844 5776 29850
rect 5724 29786 5776 29792
rect 5816 29844 5868 29850
rect 5816 29786 5868 29792
rect 5632 29640 5684 29646
rect 5632 29582 5684 29588
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5460 29238 5488 29446
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5448 29232 5500 29238
rect 5736 29186 5764 29242
rect 5448 29174 5500 29180
rect 5540 29164 5592 29170
rect 5540 29106 5592 29112
rect 5644 29158 5764 29186
rect 5172 29096 5224 29102
rect 5172 29038 5224 29044
rect 5552 29050 5580 29106
rect 5644 29050 5672 29158
rect 5552 29022 5672 29050
rect 5540 28960 5592 28966
rect 5092 28886 5212 28914
rect 5540 28902 5592 28908
rect 5080 27532 5132 27538
rect 5000 27492 5080 27520
rect 4436 26988 4488 26994
rect 4436 26930 4488 26936
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 3608 26784 3660 26790
rect 3608 26726 3660 26732
rect 3160 26438 3280 26466
rect 1308 24744 1360 24750
rect 1308 24686 1360 24692
rect 1320 24585 1348 24686
rect 1306 24576 1362 24585
rect 1306 24511 1362 24520
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 3068 22778 3096 23598
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 3068 22234 3096 22714
rect 3056 22228 3108 22234
rect 3056 22170 3108 22176
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 1320 21078 1348 21111
rect 1308 21072 1360 21078
rect 1308 21014 1360 21020
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18465 1348 18770
rect 1306 18456 1362 18465
rect 1306 18391 1362 18400
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 3068 17338 3096 17478
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 1306 17096 1362 17105
rect 1306 17031 1308 17040
rect 1360 17031 1362 17040
rect 1308 17002 1360 17008
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 1306 15736 1362 15745
rect 1306 15671 1362 15680
rect 1320 15638 1348 15671
rect 1308 15632 1360 15638
rect 1308 15574 1360 15580
rect 3068 14482 3096 15982
rect 3056 14476 3108 14482
rect 3056 14418 3108 14424
rect 1306 14376 1362 14385
rect 1306 14311 1362 14320
rect 1320 13938 1348 14311
rect 1308 13932 1360 13938
rect 1308 13874 1360 13880
rect 1308 13320 1360 13326
rect 1308 13262 1360 13268
rect 1320 13025 1348 13262
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1306 11656 1362 11665
rect 1306 11591 1362 11600
rect 1320 11286 1348 11591
rect 1308 11280 1360 11286
rect 1308 11222 1360 11228
rect 1306 9616 1362 9625
rect 1306 9551 1308 9560
rect 1360 9551 1362 9560
rect 1308 9522 1360 9528
rect 3160 9382 3188 26438
rect 3240 26376 3292 26382
rect 3240 26318 3292 26324
rect 3252 25945 3280 26318
rect 3238 25936 3294 25945
rect 3238 25871 3294 25880
rect 3516 23724 3568 23730
rect 3516 23666 3568 23672
rect 3528 23225 3556 23666
rect 3514 23216 3570 23225
rect 3514 23151 3570 23160
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3436 22234 3464 23054
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3252 21418 3280 21830
rect 3240 21412 3292 21418
rect 3240 21354 3292 21360
rect 3238 19816 3294 19825
rect 3238 19751 3294 19760
rect 3252 19310 3280 19751
rect 3240 19304 3292 19310
rect 3240 19246 3292 19252
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18426 3280 18566
rect 3620 18426 3648 26726
rect 4632 26586 4660 26930
rect 4896 26920 4948 26926
rect 4896 26862 4948 26868
rect 4908 26790 4936 26862
rect 4896 26784 4948 26790
rect 4896 26726 4948 26732
rect 4620 26580 4672 26586
rect 4620 26522 4672 26528
rect 4252 26444 4304 26450
rect 4252 26386 4304 26392
rect 3884 25696 3936 25702
rect 3884 25638 3936 25644
rect 3896 25430 3924 25638
rect 4264 25430 4292 26386
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 3884 25424 3936 25430
rect 3884 25366 3936 25372
rect 4252 25424 4304 25430
rect 4252 25366 4304 25372
rect 4264 24818 4292 25366
rect 4816 25362 4844 25774
rect 4804 25356 4856 25362
rect 4804 25298 4856 25304
rect 4342 24848 4398 24857
rect 4252 24812 4304 24818
rect 4342 24783 4398 24792
rect 4252 24754 4304 24760
rect 4356 24750 4384 24783
rect 4344 24744 4396 24750
rect 4344 24686 4396 24692
rect 4816 24070 4844 25298
rect 4908 24818 4936 26726
rect 5000 25906 5028 27492
rect 5080 27474 5132 27480
rect 4988 25900 5040 25906
rect 4988 25842 5040 25848
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4908 24614 4936 24754
rect 4896 24608 4948 24614
rect 4896 24550 4948 24556
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 4816 22982 4844 24006
rect 3792 22976 3844 22982
rect 3792 22918 3844 22924
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 3804 22166 3832 22918
rect 4080 22642 4108 22918
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 4816 22574 4844 22918
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4724 22234 4752 22374
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4816 22166 4844 22510
rect 3792 22160 3844 22166
rect 3792 22102 3844 22108
rect 4804 22160 4856 22166
rect 4804 22102 4856 22108
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4252 21888 4304 21894
rect 4252 21830 4304 21836
rect 4264 20466 4292 21830
rect 4540 21690 4568 21966
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 4816 21486 4844 22102
rect 4908 21894 4936 24550
rect 5000 23730 5028 25842
rect 5080 24336 5132 24342
rect 5080 24278 5132 24284
rect 5092 23866 5120 24278
rect 5080 23860 5132 23866
rect 5080 23802 5132 23808
rect 4988 23724 5040 23730
rect 5040 23684 5120 23712
rect 4988 23666 5040 23672
rect 5092 22574 5120 23684
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5092 22030 5120 22510
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 4896 21888 4948 21894
rect 4896 21830 4948 21836
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 4528 21412 4580 21418
rect 4528 21354 4580 21360
rect 4344 21344 4396 21350
rect 4344 21286 4396 21292
rect 4356 20466 4384 21286
rect 4540 21146 4568 21354
rect 4528 21140 4580 21146
rect 4528 21082 4580 21088
rect 4436 21004 4488 21010
rect 4436 20946 4488 20952
rect 4252 20460 4304 20466
rect 4252 20402 4304 20408
rect 4344 20460 4396 20466
rect 4344 20402 4396 20408
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 3712 18834 3740 20198
rect 4264 20074 4292 20402
rect 4264 20046 4384 20074
rect 3700 18828 3752 18834
rect 3700 18770 3752 18776
rect 3240 18420 3292 18426
rect 3240 18362 3292 18368
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3436 17746 3464 18022
rect 3424 17740 3476 17746
rect 3424 17682 3476 17688
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 4172 16538 4200 17478
rect 4356 17202 4384 20046
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4252 16652 4304 16658
rect 4252 16594 4304 16600
rect 4080 16510 4200 16538
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 3252 15978 3280 16390
rect 4080 16114 4108 16510
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 3240 15972 3292 15978
rect 3240 15914 3292 15920
rect 4264 15706 4292 16594
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 4356 16250 4384 16526
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4356 15570 4384 16186
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4448 15026 4476 20946
rect 4620 19984 4672 19990
rect 4620 19926 4672 19932
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 4540 18970 4568 19790
rect 4632 19310 4660 19926
rect 4816 19854 4844 21422
rect 5184 21162 5212 28886
rect 5552 28762 5580 28902
rect 5540 28756 5592 28762
rect 5540 28698 5592 28704
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5368 28218 5396 28494
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5552 27538 5580 28698
rect 5540 27532 5592 27538
rect 5540 27474 5592 27480
rect 5264 27464 5316 27470
rect 5264 27406 5316 27412
rect 5356 27464 5408 27470
rect 5356 27406 5408 27412
rect 5276 27130 5304 27406
rect 5264 27124 5316 27130
rect 5264 27066 5316 27072
rect 5368 22234 5396 27406
rect 5644 27062 5672 29022
rect 5920 28994 5948 32166
rect 6012 31940 6040 32370
rect 6012 31912 6224 31940
rect 6196 31822 6224 31912
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 6472 31754 6500 32370
rect 6920 31884 6972 31890
rect 6920 31826 6972 31832
rect 6380 31726 6500 31754
rect 6380 31210 6408 31726
rect 6550 31580 6858 31589
rect 6550 31578 6556 31580
rect 6612 31578 6636 31580
rect 6692 31578 6716 31580
rect 6772 31578 6796 31580
rect 6852 31578 6858 31580
rect 6612 31526 6614 31578
rect 6794 31526 6796 31578
rect 6550 31524 6556 31526
rect 6612 31524 6636 31526
rect 6692 31524 6716 31526
rect 6772 31524 6796 31526
rect 6852 31524 6858 31526
rect 6550 31515 6858 31524
rect 6932 31278 6960 31826
rect 7024 31414 7052 32422
rect 7210 32124 7518 32133
rect 7210 32122 7216 32124
rect 7272 32122 7296 32124
rect 7352 32122 7376 32124
rect 7432 32122 7456 32124
rect 7512 32122 7518 32124
rect 7272 32070 7274 32122
rect 7454 32070 7456 32122
rect 7210 32068 7216 32070
rect 7272 32068 7296 32070
rect 7352 32068 7376 32070
rect 7432 32068 7456 32070
rect 7512 32068 7518 32070
rect 7210 32059 7518 32068
rect 7944 31890 7972 33390
rect 7932 31884 7984 31890
rect 7932 31826 7984 31832
rect 7012 31408 7064 31414
rect 7012 31350 7064 31356
rect 6920 31272 6972 31278
rect 6920 31214 6972 31220
rect 7840 31272 7892 31278
rect 7840 31214 7892 31220
rect 6368 31204 6420 31210
rect 6368 31146 6420 31152
rect 6380 30938 6408 31146
rect 6368 30932 6420 30938
rect 6368 30874 6420 30880
rect 6380 30258 6408 30874
rect 6550 30492 6858 30501
rect 6550 30490 6556 30492
rect 6612 30490 6636 30492
rect 6692 30490 6716 30492
rect 6772 30490 6796 30492
rect 6852 30490 6858 30492
rect 6612 30438 6614 30490
rect 6794 30438 6796 30490
rect 6550 30436 6556 30438
rect 6612 30436 6636 30438
rect 6692 30436 6716 30438
rect 6772 30436 6796 30438
rect 6852 30436 6858 30438
rect 6550 30427 6858 30436
rect 6932 30410 6960 31214
rect 7210 31036 7518 31045
rect 7210 31034 7216 31036
rect 7272 31034 7296 31036
rect 7352 31034 7376 31036
rect 7432 31034 7456 31036
rect 7512 31034 7518 31036
rect 7272 30982 7274 31034
rect 7454 30982 7456 31034
rect 7210 30980 7216 30982
rect 7272 30980 7296 30982
rect 7352 30980 7376 30982
rect 7432 30980 7456 30982
rect 7512 30980 7518 30982
rect 7210 30971 7518 30980
rect 6932 30382 7236 30410
rect 6000 30252 6052 30258
rect 6000 30194 6052 30200
rect 6368 30252 6420 30258
rect 6368 30194 6420 30200
rect 7012 30252 7064 30258
rect 7012 30194 7064 30200
rect 6012 29186 6040 30194
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6840 29646 6868 30126
rect 6828 29640 6880 29646
rect 6828 29582 6880 29588
rect 6920 29640 6972 29646
rect 6920 29582 6972 29588
rect 6550 29404 6858 29413
rect 6550 29402 6556 29404
rect 6612 29402 6636 29404
rect 6692 29402 6716 29404
rect 6772 29402 6796 29404
rect 6852 29402 6858 29404
rect 6612 29350 6614 29402
rect 6794 29350 6796 29402
rect 6550 29348 6556 29350
rect 6612 29348 6636 29350
rect 6692 29348 6716 29350
rect 6772 29348 6796 29350
rect 6852 29348 6858 29350
rect 6550 29339 6858 29348
rect 6932 29306 6960 29582
rect 6920 29300 6972 29306
rect 6920 29242 6972 29248
rect 6012 29158 6500 29186
rect 6368 29028 6420 29034
rect 5920 28966 6040 28994
rect 6368 28970 6420 28976
rect 6012 27334 6040 28966
rect 5816 27328 5868 27334
rect 5816 27270 5868 27276
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 5632 27056 5684 27062
rect 5632 26998 5684 27004
rect 5540 26852 5592 26858
rect 5540 26794 5592 26800
rect 5724 26852 5776 26858
rect 5724 26794 5776 26800
rect 5552 24970 5580 26794
rect 5736 26586 5764 26794
rect 5828 26586 5856 27270
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5460 24942 5580 24970
rect 5644 24954 5672 25230
rect 5908 25152 5960 25158
rect 5908 25094 5960 25100
rect 5920 24993 5948 25094
rect 5906 24984 5962 24993
rect 5632 24948 5684 24954
rect 5460 24614 5488 24942
rect 5906 24919 5962 24928
rect 5632 24890 5684 24896
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5448 24608 5500 24614
rect 5448 24550 5500 24556
rect 5552 23254 5580 24754
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5540 23248 5592 23254
rect 5540 23190 5592 23196
rect 5448 23180 5500 23186
rect 5448 23122 5500 23128
rect 5460 22982 5488 23122
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5644 22778 5672 24550
rect 5816 24268 5868 24274
rect 5816 24210 5868 24216
rect 5828 23526 5856 24210
rect 6012 24018 6040 27270
rect 6380 27130 6408 28970
rect 6092 27124 6144 27130
rect 6092 27066 6144 27072
rect 6368 27124 6420 27130
rect 6368 27066 6420 27072
rect 6104 24138 6132 27066
rect 6184 26920 6236 26926
rect 6184 26862 6236 26868
rect 6276 26920 6328 26926
rect 6276 26862 6328 26868
rect 6196 26586 6224 26862
rect 6184 26580 6236 26586
rect 6184 26522 6236 26528
rect 6196 25430 6224 26522
rect 6184 25424 6236 25430
rect 6184 25366 6236 25372
rect 6184 24608 6236 24614
rect 6184 24550 6236 24556
rect 6196 24274 6224 24550
rect 6288 24410 6316 26862
rect 6368 26240 6420 26246
rect 6368 26182 6420 26188
rect 6380 25906 6408 26182
rect 6368 25900 6420 25906
rect 6368 25842 6420 25848
rect 6472 25344 6500 29158
rect 7024 28558 7052 30194
rect 7208 30190 7236 30382
rect 7196 30184 7248 30190
rect 7196 30126 7248 30132
rect 7210 29948 7518 29957
rect 7210 29946 7216 29948
rect 7272 29946 7296 29948
rect 7352 29946 7376 29948
rect 7432 29946 7456 29948
rect 7512 29946 7518 29948
rect 7272 29894 7274 29946
rect 7454 29894 7456 29946
rect 7210 29892 7216 29894
rect 7272 29892 7296 29894
rect 7352 29892 7376 29894
rect 7432 29892 7456 29894
rect 7512 29892 7518 29894
rect 7210 29883 7518 29892
rect 7564 29640 7616 29646
rect 7564 29582 7616 29588
rect 7576 29170 7604 29582
rect 7564 29164 7616 29170
rect 7564 29106 7616 29112
rect 7210 28860 7518 28869
rect 7210 28858 7216 28860
rect 7272 28858 7296 28860
rect 7352 28858 7376 28860
rect 7432 28858 7456 28860
rect 7512 28858 7518 28860
rect 7272 28806 7274 28858
rect 7454 28806 7456 28858
rect 7210 28804 7216 28806
rect 7272 28804 7296 28806
rect 7352 28804 7376 28806
rect 7432 28804 7456 28806
rect 7512 28804 7518 28806
rect 7210 28795 7518 28804
rect 7576 28694 7604 29106
rect 7564 28688 7616 28694
rect 7564 28630 7616 28636
rect 7012 28552 7064 28558
rect 7012 28494 7064 28500
rect 6550 28316 6858 28325
rect 6550 28314 6556 28316
rect 6612 28314 6636 28316
rect 6692 28314 6716 28316
rect 6772 28314 6796 28316
rect 6852 28314 6858 28316
rect 6612 28262 6614 28314
rect 6794 28262 6796 28314
rect 6550 28260 6556 28262
rect 6612 28260 6636 28262
rect 6692 28260 6716 28262
rect 6772 28260 6796 28262
rect 6852 28260 6858 28262
rect 6550 28251 6858 28260
rect 6736 27940 6788 27946
rect 6736 27882 6788 27888
rect 6748 27674 6776 27882
rect 6736 27668 6788 27674
rect 6736 27610 6788 27616
rect 7024 27606 7052 28494
rect 7576 27878 7604 28630
rect 7852 28082 7880 31214
rect 7944 31142 7972 31826
rect 8220 31754 8248 33798
rect 8944 33380 8996 33386
rect 8944 33322 8996 33328
rect 8956 33114 8984 33322
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 8944 32360 8996 32366
rect 8944 32302 8996 32308
rect 8392 32224 8444 32230
rect 8392 32166 8444 32172
rect 8404 31958 8432 32166
rect 8392 31952 8444 31958
rect 8392 31894 8444 31900
rect 8128 31726 8248 31754
rect 7932 31136 7984 31142
rect 7932 31078 7984 31084
rect 7944 30258 7972 31078
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 7944 29714 7972 29990
rect 7932 29708 7984 29714
rect 7932 29650 7984 29656
rect 7944 28762 7972 29650
rect 7932 28756 7984 28762
rect 7932 28698 7984 28704
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 7210 27772 7518 27781
rect 7210 27770 7216 27772
rect 7272 27770 7296 27772
rect 7352 27770 7376 27772
rect 7432 27770 7456 27772
rect 7512 27770 7518 27772
rect 7272 27718 7274 27770
rect 7454 27718 7456 27770
rect 7210 27716 7216 27718
rect 7272 27716 7296 27718
rect 7352 27716 7376 27718
rect 7432 27716 7456 27718
rect 7512 27716 7518 27718
rect 7210 27707 7518 27716
rect 7012 27600 7064 27606
rect 7012 27542 7064 27548
rect 7104 27532 7156 27538
rect 7104 27474 7156 27480
rect 7564 27532 7616 27538
rect 7564 27474 7616 27480
rect 6550 27228 6858 27237
rect 6550 27226 6556 27228
rect 6612 27226 6636 27228
rect 6692 27226 6716 27228
rect 6772 27226 6796 27228
rect 6852 27226 6858 27228
rect 6612 27174 6614 27226
rect 6794 27174 6796 27226
rect 6550 27172 6556 27174
rect 6612 27172 6636 27174
rect 6692 27172 6716 27174
rect 6772 27172 6796 27174
rect 6852 27172 6858 27174
rect 6550 27163 6858 27172
rect 7116 26772 7144 27474
rect 7196 26784 7248 26790
rect 7116 26744 7196 26772
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 6550 26140 6858 26149
rect 6550 26138 6556 26140
rect 6612 26138 6636 26140
rect 6692 26138 6716 26140
rect 6772 26138 6796 26140
rect 6852 26138 6858 26140
rect 6612 26086 6614 26138
rect 6794 26086 6796 26138
rect 6550 26084 6556 26086
rect 6612 26084 6636 26086
rect 6692 26084 6716 26086
rect 6772 26084 6796 26086
rect 6852 26084 6858 26086
rect 6550 26075 6858 26084
rect 6932 25498 6960 26318
rect 6920 25492 6972 25498
rect 6920 25434 6972 25440
rect 6380 25316 6500 25344
rect 6552 25356 6604 25362
rect 6380 24886 6408 25316
rect 6552 25298 6604 25304
rect 6460 25220 6512 25226
rect 6460 25162 6512 25168
rect 6368 24880 6420 24886
rect 6368 24822 6420 24828
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 6276 24404 6328 24410
rect 6276 24346 6328 24352
rect 6184 24268 6236 24274
rect 6184 24210 6236 24216
rect 6092 24132 6144 24138
rect 6092 24074 6144 24080
rect 6012 23990 6132 24018
rect 6000 23860 6052 23866
rect 6000 23802 6052 23808
rect 5908 23724 5960 23730
rect 5908 23666 5960 23672
rect 5816 23520 5868 23526
rect 5814 23488 5816 23497
rect 5868 23488 5870 23497
rect 5814 23423 5870 23432
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5264 22024 5316 22030
rect 5264 21966 5316 21972
rect 5092 21134 5212 21162
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4620 19304 4672 19310
rect 4620 19246 4672 19252
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4816 18902 4844 19790
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 5000 18766 5028 19654
rect 4988 18760 5040 18766
rect 4988 18702 5040 18708
rect 5092 18222 5120 21134
rect 5172 21072 5224 21078
rect 5172 21014 5224 21020
rect 5184 20602 5212 21014
rect 5172 20596 5224 20602
rect 5172 20538 5224 20544
rect 5276 19922 5304 21966
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 20058 5396 20198
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5184 19417 5212 19450
rect 5170 19408 5226 19417
rect 5276 19378 5304 19858
rect 5170 19343 5226 19352
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5276 18970 5304 19314
rect 5264 18964 5316 18970
rect 5264 18906 5316 18912
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4540 16794 4568 17614
rect 4528 16788 4580 16794
rect 4528 16730 4580 16736
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4344 15020 4396 15026
rect 4344 14962 4396 14968
rect 4436 15020 4488 15026
rect 4436 14962 4488 14968
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4172 14618 4200 14758
rect 4160 14612 4212 14618
rect 4160 14554 4212 14560
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3896 12442 3924 12718
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3988 12238 4016 12922
rect 4080 12238 4108 13330
rect 4356 12986 4384 14962
rect 4448 14346 4476 14962
rect 4436 14340 4488 14346
rect 4436 14282 4488 14288
rect 4540 14074 4568 16526
rect 4724 15638 4752 18158
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5080 17196 5132 17202
rect 5080 17138 5132 17144
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4816 16794 4844 16934
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4712 15632 4764 15638
rect 4712 15574 4764 15580
rect 4724 14498 4752 15574
rect 5092 15094 5120 17138
rect 5276 16794 5304 18090
rect 5460 17882 5488 22510
rect 5644 22094 5672 22714
rect 5644 22066 5764 22094
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5538 21040 5594 21049
rect 5538 20975 5540 20984
rect 5592 20975 5594 20984
rect 5540 20946 5592 20952
rect 5644 20890 5672 21286
rect 5552 20862 5672 20890
rect 5552 19854 5580 20862
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5552 19514 5580 19790
rect 5540 19508 5592 19514
rect 5540 19450 5592 19456
rect 5644 19446 5672 20402
rect 5736 20346 5764 22066
rect 5816 21684 5868 21690
rect 5816 21626 5868 21632
rect 5828 21010 5856 21626
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5920 20466 5948 23666
rect 6012 22438 6040 23802
rect 6000 22432 6052 22438
rect 6000 22374 6052 22380
rect 6000 21956 6052 21962
rect 6000 21898 6052 21904
rect 6012 21554 6040 21898
rect 6104 21554 6132 23990
rect 6196 23633 6224 24210
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6288 23866 6316 24006
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 6380 23730 6408 24550
rect 6472 24410 6500 25162
rect 6564 25140 6592 25298
rect 6920 25152 6972 25158
rect 6564 25112 6920 25140
rect 6920 25094 6972 25100
rect 6550 25052 6858 25061
rect 6550 25050 6556 25052
rect 6612 25050 6636 25052
rect 6692 25050 6716 25052
rect 6772 25050 6796 25052
rect 6852 25050 6858 25052
rect 6612 24998 6614 25050
rect 6794 24998 6796 25050
rect 6550 24996 6556 24998
rect 6612 24996 6636 24998
rect 6692 24996 6716 24998
rect 6772 24996 6796 24998
rect 6852 24996 6858 24998
rect 6550 24987 6858 24996
rect 6552 24880 6604 24886
rect 6552 24822 6604 24828
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 6564 24052 6592 24822
rect 6736 24744 6788 24750
rect 6736 24686 6788 24692
rect 6748 24410 6776 24686
rect 6932 24614 6960 25094
rect 6920 24608 6972 24614
rect 6920 24550 6972 24556
rect 7012 24608 7064 24614
rect 7012 24550 7064 24556
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6932 24206 6960 24550
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 6472 24024 6592 24052
rect 6472 23866 6500 24024
rect 6550 23964 6858 23973
rect 6550 23962 6556 23964
rect 6612 23962 6636 23964
rect 6692 23962 6716 23964
rect 6772 23962 6796 23964
rect 6852 23962 6858 23964
rect 6612 23910 6614 23962
rect 6794 23910 6796 23962
rect 6550 23908 6556 23910
rect 6612 23908 6636 23910
rect 6692 23908 6716 23910
rect 6772 23908 6796 23910
rect 6852 23908 6858 23910
rect 6550 23899 6858 23908
rect 6460 23860 6512 23866
rect 6460 23802 6512 23808
rect 6828 23860 6880 23866
rect 6828 23802 6880 23808
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 6182 23624 6238 23633
rect 6182 23559 6238 23568
rect 6840 22964 6868 23802
rect 6932 23100 6960 24142
rect 7024 24070 7052 24550
rect 7012 24064 7064 24070
rect 7012 24006 7064 24012
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 7024 23254 7052 23462
rect 7012 23248 7064 23254
rect 7012 23190 7064 23196
rect 6932 23072 7052 23100
rect 6840 22936 6960 22964
rect 6550 22876 6858 22885
rect 6550 22874 6556 22876
rect 6612 22874 6636 22876
rect 6692 22874 6716 22876
rect 6772 22874 6796 22876
rect 6852 22874 6858 22876
rect 6612 22822 6614 22874
rect 6794 22822 6796 22874
rect 6550 22820 6556 22822
rect 6612 22820 6636 22822
rect 6692 22820 6716 22822
rect 6772 22820 6796 22822
rect 6852 22820 6858 22822
rect 6550 22811 6858 22820
rect 6460 22432 6512 22438
rect 6460 22374 6512 22380
rect 6472 21570 6500 22374
rect 6550 21788 6858 21797
rect 6550 21786 6556 21788
rect 6612 21786 6636 21788
rect 6692 21786 6716 21788
rect 6772 21786 6796 21788
rect 6852 21786 6858 21788
rect 6612 21734 6614 21786
rect 6794 21734 6796 21786
rect 6550 21732 6556 21734
rect 6612 21732 6636 21734
rect 6692 21732 6716 21734
rect 6772 21732 6796 21734
rect 6852 21732 6858 21734
rect 6550 21723 6858 21732
rect 6932 21622 6960 22936
rect 6000 21548 6052 21554
rect 6000 21490 6052 21496
rect 6092 21548 6144 21554
rect 6092 21490 6144 21496
rect 6380 21542 6500 21570
rect 6920 21616 6972 21622
rect 6920 21558 6972 21564
rect 6092 21412 6144 21418
rect 6092 21354 6144 21360
rect 6104 21146 6132 21354
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6092 21140 6144 21146
rect 6092 21082 6144 21088
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5736 20318 5948 20346
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5814 20224 5870 20233
rect 5736 19786 5764 20198
rect 5814 20159 5870 20168
rect 5828 19922 5856 20159
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5724 19780 5776 19786
rect 5724 19722 5776 19728
rect 5632 19440 5684 19446
rect 5632 19382 5684 19388
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5552 18902 5580 19110
rect 5540 18896 5592 18902
rect 5540 18838 5592 18844
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5368 16794 5396 17682
rect 5264 16788 5316 16794
rect 5264 16730 5316 16736
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5276 16114 5304 16730
rect 5264 16108 5316 16114
rect 5316 16068 5396 16096
rect 5264 16050 5316 16056
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 4988 14544 5040 14550
rect 4724 14470 4844 14498
rect 4988 14486 5040 14492
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11694 3464 12038
rect 3424 11688 3476 11694
rect 3424 11630 3476 11636
rect 3988 11098 4016 12174
rect 4080 11898 4108 12174
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3896 11082 4016 11098
rect 3896 11076 4028 11082
rect 3896 11070 3976 11076
rect 3516 10532 3568 10538
rect 3516 10474 3568 10480
rect 3528 10266 3556 10474
rect 3516 10260 3568 10266
rect 3516 10202 3568 10208
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3240 9104 3292 9110
rect 3240 9046 3292 9052
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1320 7954 1348 8191
rect 3252 8090 3280 9046
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 8634 3464 8774
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 1308 7948 1360 7954
rect 1308 7890 1360 7896
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3160 6934 3188 7278
rect 3148 6928 3200 6934
rect 3528 6905 3556 7346
rect 3148 6870 3200 6876
rect 3514 6896 3570 6905
rect 3056 6248 3108 6254
rect 3056 6190 3108 6196
rect 3068 5545 3096 6190
rect 3160 5914 3188 6870
rect 3514 6831 3570 6840
rect 3896 6798 3924 11070
rect 3976 11018 4028 11024
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4172 10470 4200 10610
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 3976 10124 4028 10130
rect 3976 10066 4028 10072
rect 3988 9722 4016 10066
rect 3976 9716 4028 9722
rect 3976 9658 4028 9664
rect 4172 9518 4200 10406
rect 4356 10130 4384 12786
rect 4620 12776 4672 12782
rect 4448 12724 4620 12730
rect 4448 12718 4672 12724
rect 4448 12702 4660 12718
rect 4448 12102 4476 12702
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4436 12096 4488 12102
rect 4436 12038 4488 12044
rect 4448 11218 4476 12038
rect 4540 11762 4568 12582
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4632 10538 4660 11494
rect 4724 11014 4752 14010
rect 4816 11778 4844 14470
rect 5000 14074 5028 14486
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 5184 13870 5212 14894
rect 5172 13864 5224 13870
rect 5172 13806 5224 13812
rect 5184 12238 5212 13806
rect 5276 12238 5304 15098
rect 5368 15026 5396 16068
rect 5644 15994 5672 19382
rect 5736 19378 5764 19722
rect 5828 19718 5856 19858
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5724 19372 5776 19378
rect 5724 19314 5776 19320
rect 5816 18896 5868 18902
rect 5816 18838 5868 18844
rect 5722 18320 5778 18329
rect 5828 18290 5856 18838
rect 5722 18255 5724 18264
rect 5776 18255 5778 18264
rect 5816 18284 5868 18290
rect 5724 18226 5776 18232
rect 5816 18226 5868 18232
rect 5920 17134 5948 20318
rect 6196 19922 6224 21286
rect 6380 20262 6408 21542
rect 7024 21350 7052 23072
rect 7116 22094 7144 26744
rect 7196 26726 7248 26732
rect 7210 26684 7518 26693
rect 7210 26682 7216 26684
rect 7272 26682 7296 26684
rect 7352 26682 7376 26684
rect 7432 26682 7456 26684
rect 7512 26682 7518 26684
rect 7272 26630 7274 26682
rect 7454 26630 7456 26682
rect 7210 26628 7216 26630
rect 7272 26628 7296 26630
rect 7352 26628 7376 26630
rect 7432 26628 7456 26630
rect 7512 26628 7518 26630
rect 7210 26619 7518 26628
rect 7210 25596 7518 25605
rect 7210 25594 7216 25596
rect 7272 25594 7296 25596
rect 7352 25594 7376 25596
rect 7432 25594 7456 25596
rect 7512 25594 7518 25596
rect 7272 25542 7274 25594
rect 7454 25542 7456 25594
rect 7210 25540 7216 25542
rect 7272 25540 7296 25542
rect 7352 25540 7376 25542
rect 7432 25540 7456 25542
rect 7512 25540 7518 25542
rect 7210 25531 7518 25540
rect 7210 24508 7518 24517
rect 7210 24506 7216 24508
rect 7272 24506 7296 24508
rect 7352 24506 7376 24508
rect 7432 24506 7456 24508
rect 7512 24506 7518 24508
rect 7272 24454 7274 24506
rect 7454 24454 7456 24506
rect 7210 24452 7216 24454
rect 7272 24452 7296 24454
rect 7352 24452 7376 24454
rect 7432 24452 7456 24454
rect 7512 24452 7518 24454
rect 7210 24443 7518 24452
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7484 23526 7512 24074
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7210 23420 7518 23429
rect 7210 23418 7216 23420
rect 7272 23418 7296 23420
rect 7352 23418 7376 23420
rect 7432 23418 7456 23420
rect 7512 23418 7518 23420
rect 7272 23366 7274 23418
rect 7454 23366 7456 23418
rect 7210 23364 7216 23366
rect 7272 23364 7296 23366
rect 7352 23364 7376 23366
rect 7432 23364 7456 23366
rect 7512 23364 7518 23366
rect 7210 23355 7518 23364
rect 7210 22332 7518 22341
rect 7210 22330 7216 22332
rect 7272 22330 7296 22332
rect 7352 22330 7376 22332
rect 7432 22330 7456 22332
rect 7512 22330 7518 22332
rect 7272 22278 7274 22330
rect 7454 22278 7456 22330
rect 7210 22276 7216 22278
rect 7272 22276 7296 22278
rect 7352 22276 7376 22278
rect 7432 22276 7456 22278
rect 7512 22276 7518 22278
rect 7210 22267 7518 22276
rect 7116 22066 7512 22094
rect 7484 21434 7512 22066
rect 7576 21536 7604 27474
rect 7748 27328 7800 27334
rect 7748 27270 7800 27276
rect 7656 26376 7708 26382
rect 7656 26318 7708 26324
rect 7668 26042 7696 26318
rect 7656 26036 7708 26042
rect 7656 25978 7708 25984
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 7668 24750 7696 25842
rect 7760 25158 7788 27270
rect 7852 27130 7880 28018
rect 8024 27872 8076 27878
rect 8024 27814 8076 27820
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7748 25152 7800 25158
rect 7748 25094 7800 25100
rect 7852 24818 7880 27066
rect 8036 26926 8064 27814
rect 8024 26920 8076 26926
rect 8024 26862 8076 26868
rect 8036 26450 8064 26862
rect 8024 26444 8076 26450
rect 8024 26386 8076 26392
rect 8036 25362 8064 26386
rect 8024 25356 8076 25362
rect 8024 25298 8076 25304
rect 7840 24812 7892 24818
rect 7840 24754 7892 24760
rect 7656 24744 7708 24750
rect 8128 24721 8156 31726
rect 8956 30938 8984 32302
rect 9232 32026 9260 33934
rect 10600 33924 10652 33930
rect 10600 33866 10652 33872
rect 10048 32972 10100 32978
rect 10048 32914 10100 32920
rect 10060 32570 10088 32914
rect 10140 32904 10192 32910
rect 10140 32846 10192 32852
rect 10152 32586 10180 32846
rect 10612 32842 10640 33866
rect 10784 33448 10836 33454
rect 10784 33390 10836 33396
rect 10600 32836 10652 32842
rect 10600 32778 10652 32784
rect 10048 32564 10100 32570
rect 10152 32558 10364 32586
rect 10048 32506 10100 32512
rect 9312 32224 9364 32230
rect 9312 32166 9364 32172
rect 9220 32020 9272 32026
rect 9220 31962 9272 31968
rect 9232 30938 9260 31962
rect 9324 31958 9352 32166
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 9312 31952 9364 31958
rect 9312 31894 9364 31900
rect 10152 31278 10180 31962
rect 10336 31754 10364 32558
rect 10796 32434 10824 33390
rect 10888 33289 10916 33934
rect 11060 33312 11112 33318
rect 10874 33280 10930 33289
rect 11060 33254 11112 33260
rect 11426 33280 11482 33289
rect 10874 33215 10930 33224
rect 11072 32978 11100 33254
rect 11426 33215 11482 33224
rect 11440 33114 11468 33215
rect 11624 33153 11652 35678
rect 12912 34134 12940 35678
rect 12900 34128 12952 34134
rect 12900 34070 12952 34076
rect 14200 34066 14228 35678
rect 15099 34300 15407 34309
rect 15099 34298 15105 34300
rect 15161 34298 15185 34300
rect 15241 34298 15265 34300
rect 15321 34298 15345 34300
rect 15401 34298 15407 34300
rect 15161 34246 15163 34298
rect 15343 34246 15345 34298
rect 15099 34244 15105 34246
rect 15161 34244 15185 34246
rect 15241 34244 15265 34246
rect 15321 34244 15345 34246
rect 15401 34244 15407 34246
rect 15099 34235 15407 34244
rect 15488 34202 15516 35678
rect 15476 34196 15528 34202
rect 15476 34138 15528 34144
rect 12624 34060 12676 34066
rect 12624 34002 12676 34008
rect 13360 34060 13412 34066
rect 13360 34002 13412 34008
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 11704 33992 11756 33998
rect 11704 33934 11756 33940
rect 11610 33144 11666 33153
rect 11428 33108 11480 33114
rect 11716 33114 11744 33934
rect 12256 33856 12308 33862
rect 12256 33798 12308 33804
rect 12440 33856 12492 33862
rect 12440 33798 12492 33804
rect 12268 33522 12296 33798
rect 12256 33516 12308 33522
rect 12256 33458 12308 33464
rect 12452 33386 12480 33798
rect 12636 33658 12664 34002
rect 12624 33652 12676 33658
rect 12624 33594 12676 33600
rect 12440 33380 12492 33386
rect 12440 33322 12492 33328
rect 12532 33312 12584 33318
rect 12532 33254 12584 33260
rect 12544 33114 12572 33254
rect 11610 33079 11666 33088
rect 11704 33108 11756 33114
rect 11428 33050 11480 33056
rect 11704 33050 11756 33056
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 11888 33040 11940 33046
rect 12070 33008 12126 33017
rect 11888 32982 11940 32988
rect 10968 32972 11020 32978
rect 10968 32914 11020 32920
rect 11060 32972 11112 32978
rect 11112 32932 11192 32960
rect 11060 32914 11112 32920
rect 10980 32858 11008 32914
rect 11058 32872 11114 32881
rect 10980 32830 11058 32858
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10692 31884 10744 31890
rect 10692 31826 10744 31832
rect 10244 31726 10364 31754
rect 10140 31272 10192 31278
rect 10140 31214 10192 31220
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9784 30938 9812 31078
rect 8944 30932 8996 30938
rect 8944 30874 8996 30880
rect 9220 30932 9272 30938
rect 9220 30874 9272 30880
rect 9772 30932 9824 30938
rect 9772 30874 9824 30880
rect 8300 30796 8352 30802
rect 8300 30738 8352 30744
rect 9220 30796 9272 30802
rect 9220 30738 9272 30744
rect 8208 30592 8260 30598
rect 8208 30534 8260 30540
rect 8220 30122 8248 30534
rect 8208 30116 8260 30122
rect 8208 30058 8260 30064
rect 8312 29646 8340 30738
rect 9232 30258 9260 30738
rect 9600 30654 9812 30682
rect 9600 30598 9628 30654
rect 9588 30592 9640 30598
rect 9588 30534 9640 30540
rect 9680 30592 9732 30598
rect 9680 30534 9732 30540
rect 9692 30410 9720 30534
rect 9600 30382 9720 30410
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 8852 30116 8904 30122
rect 8852 30058 8904 30064
rect 8864 29850 8892 30058
rect 9600 29850 9628 30382
rect 9784 30054 9812 30654
rect 10244 30410 10272 31726
rect 10600 31680 10652 31686
rect 10600 31622 10652 31628
rect 10612 31346 10640 31622
rect 10600 31340 10652 31346
rect 10600 31282 10652 31288
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 10060 30382 10272 30410
rect 10336 30394 10364 31078
rect 10704 30666 10732 31826
rect 10796 30802 10824 32370
rect 10980 32042 11008 32830
rect 11058 32807 11114 32816
rect 11164 32774 11192 32932
rect 11704 32836 11756 32842
rect 11704 32778 11756 32784
rect 11060 32768 11112 32774
rect 11060 32710 11112 32716
rect 11152 32768 11204 32774
rect 11152 32710 11204 32716
rect 11072 32298 11100 32710
rect 11716 32366 11744 32778
rect 11900 32570 11928 32982
rect 11992 32978 12070 32994
rect 11980 32972 12070 32978
rect 12032 32966 12070 32972
rect 12070 32943 12126 32952
rect 12164 32972 12216 32978
rect 11980 32914 12032 32920
rect 12164 32914 12216 32920
rect 12070 32872 12126 32881
rect 12176 32858 12204 32914
rect 12126 32830 12204 32858
rect 12256 32904 12308 32910
rect 12256 32846 12308 32852
rect 12070 32807 12126 32816
rect 11888 32564 11940 32570
rect 11888 32506 11940 32512
rect 12268 32434 12296 32846
rect 12256 32428 12308 32434
rect 12256 32370 12308 32376
rect 11704 32360 11756 32366
rect 11704 32302 11756 32308
rect 12348 32360 12400 32366
rect 12348 32302 12400 32308
rect 12532 32360 12584 32366
rect 12532 32302 12584 32308
rect 11060 32292 11112 32298
rect 11060 32234 11112 32240
rect 10980 32014 11100 32042
rect 11072 31958 11100 32014
rect 11060 31952 11112 31958
rect 11060 31894 11112 31900
rect 10876 31884 10928 31890
rect 10876 31826 10928 31832
rect 10968 31884 11020 31890
rect 10968 31826 11020 31832
rect 10888 31686 10916 31826
rect 10876 31680 10928 31686
rect 10876 31622 10928 31628
rect 10980 31278 11008 31826
rect 10968 31272 11020 31278
rect 10968 31214 11020 31220
rect 10784 30796 10836 30802
rect 10784 30738 10836 30744
rect 10692 30660 10744 30666
rect 10692 30602 10744 30608
rect 10796 30598 10824 30738
rect 10784 30592 10836 30598
rect 10784 30534 10836 30540
rect 10324 30388 10376 30394
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9772 30048 9824 30054
rect 9772 29990 9824 29996
rect 8852 29844 8904 29850
rect 8852 29786 8904 29792
rect 9588 29844 9640 29850
rect 9588 29786 9640 29792
rect 9692 29782 9720 29990
rect 9680 29776 9732 29782
rect 9680 29718 9732 29724
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 9864 29640 9916 29646
rect 9916 29600 9996 29628
rect 9864 29582 9916 29588
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8312 28762 8340 28970
rect 8484 28960 8536 28966
rect 8484 28902 8536 28908
rect 8496 28762 8524 28902
rect 8300 28756 8352 28762
rect 8300 28698 8352 28704
rect 8484 28756 8536 28762
rect 8484 28698 8536 28704
rect 8208 28620 8260 28626
rect 8208 28562 8260 28568
rect 8220 27674 8248 28562
rect 9864 28552 9916 28558
rect 9864 28494 9916 28500
rect 9220 28416 9272 28422
rect 9220 28358 9272 28364
rect 9232 28218 9260 28358
rect 9876 28218 9904 28494
rect 9220 28212 9272 28218
rect 9220 28154 9272 28160
rect 9864 28212 9916 28218
rect 9864 28154 9916 28160
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 8404 27674 8432 27882
rect 8208 27668 8260 27674
rect 8208 27610 8260 27616
rect 8392 27668 8444 27674
rect 8392 27610 8444 27616
rect 8220 27130 8248 27610
rect 9968 27538 9996 29600
rect 10060 28694 10088 30382
rect 10324 30330 10376 30336
rect 10140 30048 10192 30054
rect 10140 29990 10192 29996
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10152 29170 10180 29990
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10232 29504 10284 29510
rect 10232 29446 10284 29452
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 10244 28762 10272 29446
rect 10336 28778 10364 29786
rect 10416 29708 10468 29714
rect 10416 29650 10468 29656
rect 10508 29708 10560 29714
rect 10508 29650 10560 29656
rect 10784 29708 10836 29714
rect 10784 29650 10836 29656
rect 10428 28966 10456 29650
rect 10416 28960 10468 28966
rect 10416 28902 10468 28908
rect 10232 28756 10284 28762
rect 10336 28750 10456 28778
rect 10232 28698 10284 28704
rect 10428 28694 10456 28750
rect 10048 28688 10100 28694
rect 10048 28630 10100 28636
rect 10324 28688 10376 28694
rect 10324 28630 10376 28636
rect 10416 28688 10468 28694
rect 10416 28630 10468 28636
rect 9956 27532 10008 27538
rect 9956 27474 10008 27480
rect 9588 27328 9640 27334
rect 9588 27270 9640 27276
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 9600 26858 9628 27270
rect 10060 27130 10088 28630
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 8852 26852 8904 26858
rect 8852 26794 8904 26800
rect 9588 26852 9640 26858
rect 9588 26794 9640 26800
rect 8864 26586 8892 26794
rect 8852 26580 8904 26586
rect 8852 26522 8904 26528
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9876 26042 9904 26318
rect 9864 26036 9916 26042
rect 9864 25978 9916 25984
rect 10336 25906 10364 28630
rect 10428 26858 10456 28630
rect 10520 28558 10548 29650
rect 10600 29028 10652 29034
rect 10600 28970 10652 28976
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10520 27946 10548 28494
rect 10612 28490 10640 28970
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10704 28626 10732 28902
rect 10796 28762 10824 29650
rect 10980 29646 11008 29990
rect 11072 29850 11100 31894
rect 11716 31890 11744 32302
rect 11888 32224 11940 32230
rect 11888 32166 11940 32172
rect 11900 31958 11928 32166
rect 11888 31952 11940 31958
rect 11888 31894 11940 31900
rect 12256 31952 12308 31958
rect 12360 31940 12388 32302
rect 12544 31958 12572 32302
rect 12308 31912 12388 31940
rect 12532 31952 12584 31958
rect 12256 31894 12308 31900
rect 12532 31894 12584 31900
rect 11704 31884 11756 31890
rect 11704 31826 11756 31832
rect 12164 31884 12216 31890
rect 12164 31826 12216 31832
rect 11336 31748 11388 31754
rect 11336 31690 11388 31696
rect 11348 31142 11376 31690
rect 11152 31136 11204 31142
rect 11152 31078 11204 31084
rect 11336 31136 11388 31142
rect 11336 31078 11388 31084
rect 11164 30598 11192 31078
rect 11716 30938 11744 31826
rect 11980 31680 12032 31686
rect 11980 31622 12032 31628
rect 11992 31346 12020 31622
rect 11980 31340 12032 31346
rect 11980 31282 12032 31288
rect 12176 31278 12204 31826
rect 12164 31272 12216 31278
rect 12164 31214 12216 31220
rect 11888 31204 11940 31210
rect 11888 31146 11940 31152
rect 11704 30932 11756 30938
rect 11704 30874 11756 30880
rect 11900 30870 11928 31146
rect 12268 31142 12296 31894
rect 12256 31136 12308 31142
rect 12256 31078 12308 31084
rect 12440 31136 12492 31142
rect 12440 31078 12492 31084
rect 11888 30864 11940 30870
rect 11888 30806 11940 30812
rect 12268 30802 12296 31078
rect 12452 30938 12480 31078
rect 12636 30938 12664 33594
rect 13372 33386 13400 34002
rect 17420 33998 17448 35678
rect 18420 34060 18472 34066
rect 18420 34002 18472 34008
rect 15200 33992 15252 33998
rect 15200 33934 15252 33940
rect 17408 33992 17460 33998
rect 17408 33934 17460 33940
rect 14188 33856 14240 33862
rect 14188 33798 14240 33804
rect 14200 33522 14228 33798
rect 14439 33756 14747 33765
rect 14439 33754 14445 33756
rect 14501 33754 14525 33756
rect 14581 33754 14605 33756
rect 14661 33754 14685 33756
rect 14741 33754 14747 33756
rect 14501 33702 14503 33754
rect 14683 33702 14685 33754
rect 14439 33700 14445 33702
rect 14501 33700 14525 33702
rect 14581 33700 14605 33702
rect 14661 33700 14685 33702
rect 14741 33700 14747 33702
rect 14439 33691 14747 33700
rect 14188 33516 14240 33522
rect 14188 33458 14240 33464
rect 13084 33380 13136 33386
rect 13084 33322 13136 33328
rect 13360 33380 13412 33386
rect 13360 33322 13412 33328
rect 14096 33380 14148 33386
rect 14096 33322 14148 33328
rect 13096 33289 13124 33322
rect 13082 33280 13138 33289
rect 13082 33215 13138 33224
rect 13268 32564 13320 32570
rect 13268 32506 13320 32512
rect 12808 32496 12860 32502
rect 13280 32473 13308 32506
rect 12808 32438 12860 32444
rect 13266 32464 13322 32473
rect 12820 32366 12848 32438
rect 13266 32399 13322 32408
rect 12808 32360 12860 32366
rect 12808 32302 12860 32308
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 13096 31754 13124 32166
rect 13372 31754 13400 33322
rect 14108 33130 14136 33322
rect 15212 33300 15240 33934
rect 15752 33856 15804 33862
rect 16948 33856 17000 33862
rect 15804 33816 16068 33844
rect 15752 33798 15804 33804
rect 15028 33272 15240 33300
rect 15384 33312 15436 33318
rect 13820 33108 13872 33114
rect 14108 33102 14228 33130
rect 15028 33114 15056 33272
rect 15436 33272 15516 33300
rect 15384 33254 15436 33260
rect 15099 33212 15407 33221
rect 15099 33210 15105 33212
rect 15161 33210 15185 33212
rect 15241 33210 15265 33212
rect 15321 33210 15345 33212
rect 15401 33210 15407 33212
rect 15161 33158 15163 33210
rect 15343 33158 15345 33210
rect 15099 33156 15105 33158
rect 15161 33156 15185 33158
rect 15241 33156 15265 33158
rect 15321 33156 15345 33158
rect 15401 33156 15407 33158
rect 15099 33147 15407 33156
rect 13820 33050 13872 33056
rect 13728 32768 13780 32774
rect 13728 32710 13780 32716
rect 13740 32570 13768 32710
rect 13728 32564 13780 32570
rect 13728 32506 13780 32512
rect 13832 32502 13860 33050
rect 14002 33008 14058 33017
rect 14002 32943 14004 32952
rect 14056 32943 14058 32952
rect 14096 32972 14148 32978
rect 14004 32914 14056 32920
rect 14096 32914 14148 32920
rect 13820 32496 13872 32502
rect 13820 32438 13872 32444
rect 13096 31726 13216 31754
rect 13372 31726 13492 31754
rect 12440 30932 12492 30938
rect 12440 30874 12492 30880
rect 12624 30932 12676 30938
rect 12624 30874 12676 30880
rect 12256 30796 12308 30802
rect 12256 30738 12308 30744
rect 12440 30796 12492 30802
rect 12440 30738 12492 30744
rect 12624 30796 12676 30802
rect 12624 30738 12676 30744
rect 11152 30592 11204 30598
rect 11152 30534 11204 30540
rect 11980 30592 12032 30598
rect 11980 30534 12032 30540
rect 12256 30592 12308 30598
rect 12256 30534 12308 30540
rect 11060 29844 11112 29850
rect 11060 29786 11112 29792
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 10980 28966 11008 29582
rect 11992 29306 12020 30534
rect 12268 30258 12296 30534
rect 12256 30252 12308 30258
rect 12256 30194 12308 30200
rect 12256 30048 12308 30054
rect 12256 29990 12308 29996
rect 12268 29714 12296 29990
rect 12256 29708 12308 29714
rect 12256 29650 12308 29656
rect 12072 29572 12124 29578
rect 12072 29514 12124 29520
rect 11980 29300 12032 29306
rect 11980 29242 12032 29248
rect 12084 29102 12112 29514
rect 12072 29096 12124 29102
rect 12072 29038 12124 29044
rect 10876 28960 10928 28966
rect 10876 28902 10928 28908
rect 10968 28960 11020 28966
rect 11152 28960 11204 28966
rect 10968 28902 11020 28908
rect 11072 28920 11152 28948
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10692 28620 10744 28626
rect 10692 28562 10744 28568
rect 10600 28484 10652 28490
rect 10600 28426 10652 28432
rect 10508 27940 10560 27946
rect 10508 27882 10560 27888
rect 10612 26926 10640 28426
rect 10888 28422 10916 28902
rect 10968 28756 11020 28762
rect 10968 28698 11020 28704
rect 10980 28626 11008 28698
rect 10968 28620 11020 28626
rect 10968 28562 11020 28568
rect 10876 28416 10928 28422
rect 10876 28358 10928 28364
rect 10888 28014 10916 28358
rect 10876 28008 10928 28014
rect 10876 27950 10928 27956
rect 10980 27606 11008 28562
rect 10968 27600 11020 27606
rect 10968 27542 11020 27548
rect 10784 27532 10836 27538
rect 10784 27474 10836 27480
rect 10600 26920 10652 26926
rect 10652 26880 10732 26908
rect 10600 26862 10652 26868
rect 10416 26852 10468 26858
rect 10416 26794 10468 26800
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10428 25702 10456 26794
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10612 25838 10640 26726
rect 10704 26586 10732 26880
rect 10692 26580 10744 26586
rect 10692 26522 10744 26528
rect 10704 26042 10732 26522
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10600 25832 10652 25838
rect 10600 25774 10652 25780
rect 10692 25832 10744 25838
rect 10796 25820 10824 27474
rect 10980 27470 11008 27542
rect 10968 27464 11020 27470
rect 10968 27406 11020 27412
rect 11072 27334 11100 28920
rect 11152 28902 11204 28908
rect 11336 28960 11388 28966
rect 11336 28902 11388 28908
rect 11348 28626 11376 28902
rect 11336 28620 11388 28626
rect 11336 28562 11388 28568
rect 11612 28416 11664 28422
rect 11612 28358 11664 28364
rect 11152 28076 11204 28082
rect 11152 28018 11204 28024
rect 11164 27674 11192 28018
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11428 28008 11480 28014
rect 11428 27950 11480 27956
rect 11256 27674 11284 27950
rect 11336 27940 11388 27946
rect 11336 27882 11388 27888
rect 11152 27668 11204 27674
rect 11152 27610 11204 27616
rect 11244 27668 11296 27674
rect 11244 27610 11296 27616
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11072 26994 11100 27270
rect 11348 27062 11376 27882
rect 11440 27130 11468 27950
rect 11624 27674 11652 28358
rect 12268 28150 12296 29650
rect 12452 29578 12480 30738
rect 12636 29850 12664 30738
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12624 29844 12676 29850
rect 12624 29786 12676 29792
rect 12728 29782 12756 30670
rect 12900 30048 12952 30054
rect 12900 29990 12952 29996
rect 12992 30048 13044 30054
rect 12992 29990 13044 29996
rect 12912 29782 12940 29990
rect 12716 29776 12768 29782
rect 12716 29718 12768 29724
rect 12900 29776 12952 29782
rect 12900 29718 12952 29724
rect 13004 29646 13032 29990
rect 12992 29640 13044 29646
rect 12992 29582 13044 29588
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 13084 29300 13136 29306
rect 13188 29288 13216 31726
rect 13360 31136 13412 31142
rect 13360 31078 13412 31084
rect 13372 30938 13400 31078
rect 13360 30932 13412 30938
rect 13360 30874 13412 30880
rect 13268 30592 13320 30598
rect 13268 30534 13320 30540
rect 13280 30190 13308 30534
rect 13268 30184 13320 30190
rect 13268 30126 13320 30132
rect 13188 29260 13308 29288
rect 13084 29242 13136 29248
rect 12900 29232 12952 29238
rect 13096 29209 13124 29242
rect 12900 29174 12952 29180
rect 13082 29200 13138 29209
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 12452 28218 12480 28494
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12440 28212 12492 28218
rect 12440 28154 12492 28160
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 12256 28144 12308 28150
rect 12256 28086 12308 28092
rect 11704 27872 11756 27878
rect 11704 27814 11756 27820
rect 11612 27668 11664 27674
rect 11612 27610 11664 27616
rect 11520 27328 11572 27334
rect 11520 27270 11572 27276
rect 11428 27124 11480 27130
rect 11428 27066 11480 27072
rect 11336 27056 11388 27062
rect 11336 26998 11388 27004
rect 11060 26988 11112 26994
rect 11060 26930 11112 26936
rect 10744 25792 10824 25820
rect 11060 25832 11112 25838
rect 10692 25774 10744 25780
rect 11060 25774 11112 25780
rect 10416 25696 10468 25702
rect 10416 25638 10468 25644
rect 10704 25498 10732 25774
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 8208 25424 8260 25430
rect 8208 25366 8260 25372
rect 8760 25424 8812 25430
rect 8760 25366 8812 25372
rect 7656 24686 7708 24692
rect 8114 24712 8170 24721
rect 7668 24138 7696 24686
rect 8114 24647 8170 24656
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7668 23662 7696 24074
rect 7656 23656 7708 23662
rect 7656 23598 7708 23604
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 7656 23520 7708 23526
rect 7656 23462 7708 23468
rect 7668 22114 7696 23462
rect 7852 23254 7880 23598
rect 7840 23248 7892 23254
rect 7840 23190 7892 23196
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 7748 22500 7800 22506
rect 7748 22442 7800 22448
rect 7760 22234 7788 22442
rect 7852 22234 7880 23054
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7668 22086 7788 22114
rect 7576 21508 7696 21536
rect 7484 21406 7604 21434
rect 7668 21418 7696 21508
rect 7012 21344 7064 21350
rect 7012 21286 7064 21292
rect 7210 21244 7518 21253
rect 7210 21242 7216 21244
rect 7272 21242 7296 21244
rect 7352 21242 7376 21244
rect 7432 21242 7456 21244
rect 7512 21242 7518 21244
rect 7272 21190 7274 21242
rect 7454 21190 7456 21242
rect 7210 21188 7216 21190
rect 7272 21188 7296 21190
rect 7352 21188 7376 21190
rect 7432 21188 7456 21190
rect 7512 21188 7518 21190
rect 7210 21179 7518 21188
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5644 15966 5764 15994
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5632 15904 5684 15910
rect 5632 15846 5684 15852
rect 5460 15706 5488 15846
rect 5448 15700 5500 15706
rect 5448 15642 5500 15648
rect 5644 15570 5672 15846
rect 5632 15564 5684 15570
rect 5632 15506 5684 15512
rect 5736 15434 5764 15966
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5816 15632 5868 15638
rect 5816 15574 5868 15580
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5722 15192 5778 15201
rect 5828 15162 5856 15574
rect 5920 15162 5948 15914
rect 5722 15127 5778 15136
rect 5816 15156 5868 15162
rect 5736 15094 5764 15127
rect 5816 15098 5868 15104
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 5448 14408 5500 14414
rect 5448 14350 5500 14356
rect 5460 13530 5488 14350
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5644 14074 5672 14214
rect 5828 14074 5856 14418
rect 5908 14272 5960 14278
rect 5908 14214 5960 14220
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5816 14068 5868 14074
rect 5816 14010 5868 14016
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5552 13462 5580 13670
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5920 12782 5948 14214
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5540 12708 5592 12714
rect 5540 12650 5592 12656
rect 5448 12640 5500 12646
rect 5448 12582 5500 12588
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5184 11898 5212 12174
rect 5276 11898 5304 12174
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 4816 11750 4936 11778
rect 4908 11354 4936 11750
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 5092 10606 5120 11086
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4436 10464 4488 10470
rect 4436 10406 4488 10412
rect 4344 10124 4396 10130
rect 4344 10066 4396 10072
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4264 9178 4292 9998
rect 4448 9994 4476 10406
rect 4632 10198 4660 10474
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5184 10198 5212 10406
rect 5276 10248 5304 11834
rect 5460 11626 5488 12582
rect 5552 12442 5580 12650
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5736 11898 5764 12718
rect 5816 12368 5868 12374
rect 5816 12310 5868 12316
rect 5828 11898 5856 12310
rect 5908 12096 5960 12102
rect 5908 12038 5960 12044
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5552 11014 5580 11698
rect 5816 11552 5868 11558
rect 5920 11540 5948 12038
rect 5868 11512 5948 11540
rect 5816 11494 5868 11500
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10674 5580 10950
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5552 10266 5580 10610
rect 5356 10260 5408 10266
rect 5276 10220 5356 10248
rect 4620 10192 4672 10198
rect 4620 10134 4672 10140
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 4436 9988 4488 9994
rect 4436 9930 4488 9936
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4172 8090 4200 8910
rect 4264 8090 4292 9114
rect 4448 9042 4476 9930
rect 4724 9654 4752 10134
rect 5276 9674 5304 10220
rect 5356 10202 5408 10208
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5356 9920 5408 9926
rect 5356 9862 5408 9868
rect 4712 9648 4764 9654
rect 4712 9590 4764 9596
rect 5092 9646 5304 9674
rect 4436 9036 4488 9042
rect 4436 8978 4488 8984
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 7880 4120 7886
rect 4066 7848 4068 7857
rect 4120 7848 4122 7857
rect 4066 7783 4122 7792
rect 4356 6882 4384 8434
rect 4448 8430 4476 8774
rect 5092 8634 5120 9646
rect 5368 9042 5396 9862
rect 5722 9616 5778 9625
rect 5722 9551 5778 9560
rect 5736 9518 5764 9551
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5276 8634 5304 8910
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 7886 4844 8230
rect 5368 7886 5396 8774
rect 5736 7954 5764 9454
rect 6012 9110 6040 18022
rect 6104 17338 6132 19790
rect 6380 19417 6408 20198
rect 6366 19408 6422 19417
rect 6366 19343 6422 19352
rect 6380 18902 6408 19343
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6196 17202 6224 18566
rect 6380 18086 6408 18838
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6368 17672 6420 17678
rect 6368 17614 6420 17620
rect 6472 17626 6500 20742
rect 6550 20700 6858 20709
rect 6550 20698 6556 20700
rect 6612 20698 6636 20700
rect 6692 20698 6716 20700
rect 6772 20698 6796 20700
rect 6852 20698 6858 20700
rect 6612 20646 6614 20698
rect 6794 20646 6796 20698
rect 6550 20644 6556 20646
rect 6612 20644 6636 20646
rect 6692 20644 6716 20646
rect 6772 20644 6796 20646
rect 6852 20644 6858 20646
rect 6550 20635 6858 20644
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6840 20262 6868 20538
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6550 19612 6858 19621
rect 6550 19610 6556 19612
rect 6612 19610 6636 19612
rect 6692 19610 6716 19612
rect 6772 19610 6796 19612
rect 6852 19610 6858 19612
rect 6612 19558 6614 19610
rect 6794 19558 6796 19610
rect 6550 19556 6556 19558
rect 6612 19556 6636 19558
rect 6692 19556 6716 19558
rect 6772 19556 6796 19558
rect 6852 19556 6858 19558
rect 6550 19547 6858 19556
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6748 19281 6776 19382
rect 6734 19272 6790 19281
rect 6734 19207 6790 19216
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6550 18524 6858 18533
rect 6550 18522 6556 18524
rect 6612 18522 6636 18524
rect 6692 18522 6716 18524
rect 6772 18522 6796 18524
rect 6852 18522 6858 18524
rect 6612 18470 6614 18522
rect 6794 18470 6796 18522
rect 6550 18468 6556 18470
rect 6612 18468 6636 18470
rect 6692 18468 6716 18470
rect 6772 18468 6796 18470
rect 6852 18468 6858 18470
rect 6550 18459 6858 18468
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6564 18290 6592 18362
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6932 17814 6960 19110
rect 7024 18970 7052 20198
rect 7116 19378 7144 20402
rect 7210 20156 7518 20165
rect 7210 20154 7216 20156
rect 7272 20154 7296 20156
rect 7352 20154 7376 20156
rect 7432 20154 7456 20156
rect 7512 20154 7518 20156
rect 7272 20102 7274 20154
rect 7454 20102 7456 20154
rect 7210 20100 7216 20102
rect 7272 20100 7296 20102
rect 7352 20100 7376 20102
rect 7432 20100 7456 20102
rect 7512 20100 7518 20102
rect 7210 20091 7518 20100
rect 7104 19372 7156 19378
rect 7104 19314 7156 19320
rect 7210 19068 7518 19077
rect 7210 19066 7216 19068
rect 7272 19066 7296 19068
rect 7352 19066 7376 19068
rect 7432 19066 7456 19068
rect 7512 19066 7518 19068
rect 7272 19014 7274 19066
rect 7454 19014 7456 19066
rect 7210 19012 7216 19014
rect 7272 19012 7296 19014
rect 7352 19012 7376 19014
rect 7432 19012 7456 19014
rect 7512 19012 7518 19014
rect 7210 19003 7518 19012
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7210 17980 7518 17989
rect 7210 17978 7216 17980
rect 7272 17978 7296 17980
rect 7352 17978 7376 17980
rect 7432 17978 7456 17980
rect 7512 17978 7518 17980
rect 7272 17926 7274 17978
rect 7454 17926 7456 17978
rect 7210 17924 7216 17926
rect 7272 17924 7296 17926
rect 7352 17924 7376 17926
rect 7432 17924 7456 17926
rect 7512 17924 7518 17926
rect 7210 17915 7518 17924
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6380 17338 6408 17614
rect 6472 17598 6960 17626
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6472 17270 6500 17478
rect 6550 17436 6858 17445
rect 6550 17434 6556 17436
rect 6612 17434 6636 17436
rect 6692 17434 6716 17436
rect 6772 17434 6796 17436
rect 6852 17434 6858 17436
rect 6612 17382 6614 17434
rect 6794 17382 6796 17434
rect 6550 17380 6556 17382
rect 6612 17380 6636 17382
rect 6692 17380 6716 17382
rect 6772 17380 6796 17382
rect 6852 17380 6858 17382
rect 6550 17371 6858 17380
rect 6460 17264 6512 17270
rect 6932 17252 6960 17598
rect 7104 17604 7156 17610
rect 7104 17546 7156 17552
rect 6460 17206 6512 17212
rect 6840 17224 6960 17252
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6276 17060 6328 17066
rect 6276 17002 6328 17008
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6104 11286 6132 16594
rect 6288 15910 6316 17002
rect 6380 16250 6408 17138
rect 6472 16794 6500 17206
rect 6840 17134 6868 17224
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6276 15904 6328 15910
rect 6276 15846 6328 15852
rect 6380 15586 6408 16186
rect 6472 16114 6500 16730
rect 6840 16538 6868 17070
rect 6840 16510 6960 16538
rect 6550 16348 6858 16357
rect 6550 16346 6556 16348
rect 6612 16346 6636 16348
rect 6692 16346 6716 16348
rect 6772 16346 6796 16348
rect 6852 16346 6858 16348
rect 6612 16294 6614 16346
rect 6794 16294 6796 16346
rect 6550 16292 6556 16294
rect 6612 16292 6636 16294
rect 6692 16292 6716 16294
rect 6772 16292 6796 16294
rect 6852 16292 6858 16294
rect 6550 16283 6858 16292
rect 6932 16130 6960 16510
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6840 16102 6960 16130
rect 6288 15570 6408 15586
rect 6276 15564 6408 15570
rect 6328 15558 6408 15564
rect 6276 15506 6328 15512
rect 6288 15162 6316 15506
rect 6840 15450 6868 16102
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 15706 6960 15914
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6840 15422 6960 15450
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6276 15156 6328 15162
rect 6276 15098 6328 15104
rect 6288 14958 6316 15098
rect 6276 14952 6328 14958
rect 6276 14894 6328 14900
rect 6288 14396 6316 14894
rect 6196 14368 6316 14396
rect 6196 14074 6224 14368
rect 6380 14346 6408 15302
rect 6550 15260 6858 15269
rect 6550 15258 6556 15260
rect 6612 15258 6636 15260
rect 6692 15258 6716 15260
rect 6772 15258 6796 15260
rect 6852 15258 6858 15260
rect 6612 15206 6614 15258
rect 6794 15206 6796 15258
rect 6550 15204 6556 15206
rect 6612 15204 6636 15206
rect 6692 15204 6716 15206
rect 6772 15204 6796 15206
rect 6852 15204 6858 15206
rect 6550 15195 6858 15204
rect 6932 15042 6960 15422
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 7024 15162 7052 15302
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 6840 15014 6960 15042
rect 6840 14482 6868 15014
rect 6920 14816 6972 14822
rect 6920 14758 6972 14764
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6368 14340 6420 14346
rect 6288 14300 6368 14328
rect 6184 14068 6236 14074
rect 6184 14010 6236 14016
rect 6288 13530 6316 14300
rect 6368 14282 6420 14288
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6368 13864 6420 13870
rect 6368 13806 6420 13812
rect 6472 13818 6500 14282
rect 6550 14172 6858 14181
rect 6550 14170 6556 14172
rect 6612 14170 6636 14172
rect 6692 14170 6716 14172
rect 6772 14170 6796 14172
rect 6852 14170 6858 14172
rect 6612 14118 6614 14170
rect 6794 14118 6796 14170
rect 6550 14116 6556 14118
rect 6612 14116 6636 14118
rect 6692 14116 6716 14118
rect 6772 14116 6796 14118
rect 6852 14116 6858 14118
rect 6550 14107 6858 14116
rect 6932 14006 6960 14758
rect 7116 14618 7144 17546
rect 7210 16892 7518 16901
rect 7210 16890 7216 16892
rect 7272 16890 7296 16892
rect 7352 16890 7376 16892
rect 7432 16890 7456 16892
rect 7512 16890 7518 16892
rect 7272 16838 7274 16890
rect 7454 16838 7456 16890
rect 7210 16836 7216 16838
rect 7272 16836 7296 16838
rect 7352 16836 7376 16838
rect 7432 16836 7456 16838
rect 7512 16836 7518 16838
rect 7210 16827 7518 16836
rect 7210 15804 7518 15813
rect 7210 15802 7216 15804
rect 7272 15802 7296 15804
rect 7352 15802 7376 15804
rect 7432 15802 7456 15804
rect 7512 15802 7518 15804
rect 7272 15750 7274 15802
rect 7454 15750 7456 15802
rect 7210 15748 7216 15750
rect 7272 15748 7296 15750
rect 7352 15748 7376 15750
rect 7432 15748 7456 15750
rect 7512 15748 7518 15750
rect 7210 15739 7518 15748
rect 7576 15706 7604 21406
rect 7656 21412 7708 21418
rect 7656 21354 7708 21360
rect 7656 20324 7708 20330
rect 7656 20266 7708 20272
rect 7668 20058 7696 20266
rect 7656 20052 7708 20058
rect 7656 19994 7708 20000
rect 7656 19780 7708 19786
rect 7656 19722 7708 19728
rect 7668 18970 7696 19722
rect 7760 19334 7788 22086
rect 8036 21690 8064 24142
rect 8116 22160 8168 22166
rect 8116 22102 8168 22108
rect 8024 21684 8076 21690
rect 8024 21626 8076 21632
rect 7840 21344 7892 21350
rect 7840 21286 7892 21292
rect 7852 20398 7880 21286
rect 8036 21078 8064 21626
rect 8128 21146 8156 22102
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8024 21072 8076 21078
rect 8024 21014 8076 21020
rect 8036 20466 8064 21014
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 7932 20324 7984 20330
rect 7932 20266 7984 20272
rect 7944 20058 7972 20266
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 8036 20058 8064 20198
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 8128 19446 8156 20334
rect 8116 19440 8168 19446
rect 8116 19382 8168 19388
rect 7760 19306 7972 19334
rect 7748 19236 7800 19242
rect 7748 19178 7800 19184
rect 7760 18970 7788 19178
rect 7656 18964 7708 18970
rect 7656 18906 7708 18912
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7668 17542 7696 18158
rect 7748 18080 7800 18086
rect 7748 18022 7800 18028
rect 7760 17785 7788 18022
rect 7746 17776 7802 17785
rect 7746 17711 7802 17720
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7748 17060 7800 17066
rect 7748 17002 7800 17008
rect 7760 16794 7788 17002
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7944 16454 7972 19306
rect 8024 18148 8076 18154
rect 8024 18090 8076 18096
rect 7932 16448 7984 16454
rect 7932 16390 7984 16396
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7944 15706 7972 15982
rect 7564 15700 7616 15706
rect 7564 15642 7616 15648
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7748 15632 7800 15638
rect 7748 15574 7800 15580
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7392 14822 7420 15302
rect 7760 15094 7788 15574
rect 8036 15366 8064 18090
rect 8220 17762 8248 25366
rect 8772 24954 8800 25366
rect 8852 25288 8904 25294
rect 8852 25230 8904 25236
rect 8864 24954 8892 25230
rect 8760 24948 8812 24954
rect 8760 24890 8812 24896
rect 8852 24948 8904 24954
rect 8852 24890 8904 24896
rect 9128 24812 9180 24818
rect 9128 24754 9180 24760
rect 8576 24608 8628 24614
rect 8576 24550 8628 24556
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 8312 23866 8340 24142
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8300 23860 8352 23866
rect 8300 23802 8352 23808
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8312 23322 8340 23598
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8496 23066 8524 24006
rect 8588 23730 8616 24550
rect 8576 23724 8628 23730
rect 8576 23666 8628 23672
rect 8588 23186 8616 23666
rect 8944 23520 8996 23526
rect 8944 23462 8996 23468
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 8496 23038 8616 23066
rect 8300 22092 8352 22098
rect 8300 22034 8352 22040
rect 8312 19718 8340 22034
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8496 20466 8524 20742
rect 8484 20460 8536 20466
rect 8484 20402 8536 20408
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8128 17734 8248 17762
rect 8024 15360 8076 15366
rect 8024 15302 8076 15308
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7748 15088 7800 15094
rect 7748 15030 7800 15036
rect 7564 14884 7616 14890
rect 7564 14826 7616 14832
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7210 14716 7518 14725
rect 7210 14714 7216 14716
rect 7272 14714 7296 14716
rect 7352 14714 7376 14716
rect 7432 14714 7456 14716
rect 7512 14714 7518 14716
rect 7272 14662 7274 14714
rect 7454 14662 7456 14714
rect 7210 14660 7216 14662
rect 7272 14660 7296 14662
rect 7352 14660 7376 14662
rect 7432 14660 7456 14662
rect 7512 14660 7518 14662
rect 7210 14651 7518 14660
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7484 14278 7512 14418
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6276 13524 6328 13530
rect 6276 13466 6328 13472
rect 6380 13394 6408 13806
rect 6472 13790 6592 13818
rect 6460 13728 6512 13734
rect 6460 13670 6512 13676
rect 6472 13462 6500 13670
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6564 13394 6592 13790
rect 7210 13628 7518 13637
rect 7210 13626 7216 13628
rect 7272 13626 7296 13628
rect 7352 13626 7376 13628
rect 7432 13626 7456 13628
rect 7512 13626 7518 13628
rect 7272 13574 7274 13626
rect 7454 13574 7456 13626
rect 7210 13572 7216 13574
rect 7272 13572 7296 13574
rect 7352 13572 7376 13574
rect 7432 13572 7456 13574
rect 7512 13572 7518 13574
rect 7210 13563 7518 13572
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6276 13184 6328 13190
rect 6276 13126 6328 13132
rect 6368 13184 6420 13190
rect 6564 13172 6592 13330
rect 6368 13126 6420 13132
rect 6472 13144 6592 13172
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 6196 12442 6224 12582
rect 6184 12436 6236 12442
rect 6184 12378 6236 12384
rect 6184 12300 6236 12306
rect 6288 12288 6316 13126
rect 6380 12306 6408 13126
rect 6472 12986 6500 13144
rect 6550 13084 6858 13093
rect 6550 13082 6556 13084
rect 6612 13082 6636 13084
rect 6692 13082 6716 13084
rect 6772 13082 6796 13084
rect 6852 13082 6858 13084
rect 6612 13030 6614 13082
rect 6794 13030 6796 13082
rect 6550 13028 6556 13030
rect 6612 13028 6636 13030
rect 6692 13028 6716 13030
rect 6772 13028 6796 13030
rect 6852 13028 6858 13030
rect 6550 13019 6858 13028
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6236 12260 6316 12288
rect 6368 12300 6420 12306
rect 6184 12242 6236 12248
rect 6368 12242 6420 12248
rect 6196 11694 6224 12242
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 6196 11286 6224 11630
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6184 11280 6236 11286
rect 6184 11222 6236 11228
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10810 6316 11086
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6472 10554 6500 12582
rect 7210 12540 7518 12549
rect 7210 12538 7216 12540
rect 7272 12538 7296 12540
rect 7352 12538 7376 12540
rect 7432 12538 7456 12540
rect 7512 12538 7518 12540
rect 7272 12486 7274 12538
rect 7454 12486 7456 12538
rect 7210 12484 7216 12486
rect 7272 12484 7296 12486
rect 7352 12484 7376 12486
rect 7432 12484 7456 12486
rect 7512 12484 7518 12486
rect 7210 12475 7518 12484
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6564 12102 6592 12310
rect 6828 12232 6880 12238
rect 7012 12232 7064 12238
rect 6880 12192 6960 12220
rect 6828 12174 6880 12180
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6550 11996 6858 12005
rect 6550 11994 6556 11996
rect 6612 11994 6636 11996
rect 6692 11994 6716 11996
rect 6772 11994 6796 11996
rect 6852 11994 6858 11996
rect 6612 11942 6614 11994
rect 6794 11942 6796 11994
rect 6550 11940 6556 11942
rect 6612 11940 6636 11942
rect 6692 11940 6716 11942
rect 6772 11940 6796 11942
rect 6852 11940 6858 11942
rect 6550 11931 6858 11940
rect 6932 11626 6960 12192
rect 7012 12174 7064 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7024 11830 7052 12174
rect 7484 11898 7512 12174
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 7210 11452 7518 11461
rect 7210 11450 7216 11452
rect 7272 11450 7296 11452
rect 7352 11450 7376 11452
rect 7432 11450 7456 11452
rect 7512 11450 7518 11452
rect 7272 11398 7274 11450
rect 7454 11398 7456 11450
rect 7210 11396 7216 11398
rect 7272 11396 7296 11398
rect 7352 11396 7376 11398
rect 7432 11396 7456 11398
rect 7512 11396 7518 11398
rect 7210 11387 7518 11396
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 6550 10908 6858 10917
rect 6550 10906 6556 10908
rect 6612 10906 6636 10908
rect 6692 10906 6716 10908
rect 6772 10906 6796 10908
rect 6852 10906 6858 10908
rect 6612 10854 6614 10906
rect 6794 10854 6796 10906
rect 6550 10852 6556 10854
rect 6612 10852 6636 10854
rect 6692 10852 6716 10854
rect 6772 10852 6796 10854
rect 6852 10852 6858 10854
rect 6550 10843 6858 10852
rect 6644 10736 6696 10742
rect 6932 10690 6960 11154
rect 6696 10684 6960 10690
rect 6644 10678 6960 10684
rect 6656 10662 6960 10678
rect 7392 10674 7420 11222
rect 7380 10668 7432 10674
rect 7024 10628 7380 10656
rect 6472 10526 6592 10554
rect 6092 10464 6144 10470
rect 6092 10406 6144 10412
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6104 10266 6132 10406
rect 6092 10260 6144 10266
rect 6368 10260 6420 10266
rect 6092 10202 6144 10208
rect 6288 10220 6368 10248
rect 6104 9586 6132 10202
rect 6092 9580 6144 9586
rect 6092 9522 6144 9528
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5920 8634 5948 8774
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 5828 8090 5856 8366
rect 6196 8294 6224 9522
rect 6184 8288 6236 8294
rect 6184 8230 6236 8236
rect 6288 8090 6316 10220
rect 6368 10202 6420 10208
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 8974 6408 9318
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 6276 8084 6328 8090
rect 6328 8044 6408 8072
rect 6276 8026 6328 8032
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 6276 7948 6328 7954
rect 6276 7890 6328 7896
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4804 7880 4856 7886
rect 4804 7822 4856 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 4264 6866 4384 6882
rect 4252 6860 4384 6866
rect 4304 6854 4384 6860
rect 4252 6802 4304 6808
rect 3884 6792 3936 6798
rect 3936 6752 4200 6780
rect 3884 6734 3936 6740
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3252 5846 3280 6598
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4080 6118 4108 6151
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3240 5840 3292 5846
rect 3240 5782 3292 5788
rect 3054 5536 3110 5545
rect 3054 5471 3110 5480
rect 4172 5234 4200 6752
rect 4264 6458 4292 6802
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4264 5914 4292 6394
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 1308 4684 1360 4690
rect 1308 4626 1360 4632
rect 1320 4185 1348 4626
rect 1306 4176 1362 4185
rect 1306 4111 1362 4120
rect 20 4004 72 4010
rect 20 3946 72 3952
rect 32 800 60 3946
rect 3252 3670 3280 5034
rect 4448 4078 4476 7822
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 4632 6934 4660 7142
rect 5276 7002 5304 7142
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 5264 6792 5316 6798
rect 5368 6780 5396 7822
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6104 7478 6132 7686
rect 6092 7472 6144 7478
rect 6092 7414 6144 7420
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 5316 6752 5396 6780
rect 5264 6734 5316 6740
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 5914 5304 6598
rect 5264 5908 5316 5914
rect 5264 5850 5316 5856
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 4896 5704 4948 5710
rect 4896 5646 4948 5652
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4540 4146 4568 4966
rect 4908 4826 4936 5646
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 5234 5028 5510
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4816 4282 4844 4558
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4436 4072 4488 4078
rect 4436 4014 4488 4020
rect 1308 3664 1360 3670
rect 1228 3612 1308 3618
rect 1228 3606 1360 3612
rect 3240 3664 3292 3670
rect 3240 3606 3292 3612
rect 1228 3590 1348 3606
rect 4908 3602 4936 4762
rect 5092 4622 5120 5714
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5276 4622 5304 4966
rect 5368 4826 5396 6752
rect 5460 4826 5488 7278
rect 6104 7002 6132 7278
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6012 6390 6040 6598
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 4896 3596 4948 3602
rect 1228 2530 1256 3590
rect 4896 3538 4948 3544
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 1320 2825 1348 3470
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 1306 2816 1362 2825
rect 1306 2751 1362 2760
rect 1228 2502 1348 2530
rect 1320 800 1348 2502
rect 2608 800 2636 2994
rect 3056 2984 3108 2990
rect 3056 2926 3108 2932
rect 3068 1465 3096 2926
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 3054 1456 3110 1465
rect 4080 1442 4108 2858
rect 3054 1391 3110 1400
rect 3896 1414 4108 1442
rect 3896 800 3924 1414
rect 5184 800 5212 3470
rect 5276 2990 5304 4558
rect 5552 4282 5580 5170
rect 5920 5030 5948 6054
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4758 5948 4966
rect 6196 4842 6224 7278
rect 6288 6934 6316 7890
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6196 4826 6316 4842
rect 6380 4826 6408 8044
rect 6472 7954 6500 10406
rect 6564 10198 6592 10526
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6550 9820 6858 9829
rect 6550 9818 6556 9820
rect 6612 9818 6636 9820
rect 6692 9818 6716 9820
rect 6772 9818 6796 9820
rect 6852 9818 6858 9820
rect 6612 9766 6614 9818
rect 6794 9766 6796 9818
rect 6550 9764 6556 9766
rect 6612 9764 6636 9766
rect 6692 9764 6716 9766
rect 6772 9764 6796 9766
rect 6852 9764 6858 9766
rect 6550 9755 6858 9764
rect 7024 9178 7052 10628
rect 7380 10610 7432 10616
rect 7210 10364 7518 10373
rect 7210 10362 7216 10364
rect 7272 10362 7296 10364
rect 7352 10362 7376 10364
rect 7432 10362 7456 10364
rect 7512 10362 7518 10364
rect 7272 10310 7274 10362
rect 7454 10310 7456 10362
rect 7210 10308 7216 10310
rect 7272 10308 7296 10310
rect 7352 10308 7376 10310
rect 7432 10308 7456 10310
rect 7512 10308 7518 10310
rect 7210 10299 7518 10308
rect 7576 9518 7604 14826
rect 7760 14618 7788 15030
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7852 14498 7880 15098
rect 7760 14470 7880 14498
rect 8036 14482 8064 15302
rect 8024 14476 8076 14482
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7668 11762 7696 12174
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7668 11286 7696 11698
rect 7760 11286 7788 14470
rect 8024 14418 8076 14424
rect 8036 13546 8064 14418
rect 8128 13682 8156 17734
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 8220 16658 8248 17206
rect 8208 16652 8260 16658
rect 8208 16594 8260 16600
rect 8220 15162 8248 16594
rect 8312 16590 8340 19654
rect 8404 18766 8432 19654
rect 8588 19242 8616 23038
rect 8956 22710 8984 23462
rect 9036 23248 9088 23254
rect 9036 23190 9088 23196
rect 9048 23118 9076 23190
rect 9036 23112 9088 23118
rect 9036 23054 9088 23060
rect 8944 22704 8996 22710
rect 8944 22646 8996 22652
rect 8956 22234 8984 22646
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8944 22228 8996 22234
rect 8944 22170 8996 22176
rect 9048 22030 9076 22374
rect 9036 22024 9088 22030
rect 9036 21966 9088 21972
rect 8852 20460 8904 20466
rect 8852 20402 8904 20408
rect 8576 19236 8628 19242
rect 8576 19178 8628 19184
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8496 18970 8524 19110
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8576 18828 8628 18834
rect 8576 18770 8628 18776
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8496 16658 8524 18702
rect 8588 18426 8616 18770
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8576 18420 8628 18426
rect 8576 18362 8628 18368
rect 8680 18329 8708 18634
rect 8666 18320 8722 18329
rect 8864 18290 8892 20402
rect 9048 20058 9076 21966
rect 9140 21418 9168 24754
rect 9692 24342 9720 25434
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10232 24744 10284 24750
rect 10232 24686 10284 24692
rect 9680 24336 9732 24342
rect 9680 24278 9732 24284
rect 9220 23656 9272 23662
rect 9220 23598 9272 23604
rect 9232 23526 9260 23598
rect 9220 23520 9272 23526
rect 9220 23462 9272 23468
rect 9232 23254 9260 23462
rect 9220 23248 9272 23254
rect 9692 23202 9720 24278
rect 10244 24018 10272 24686
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10152 23990 10272 24018
rect 9956 23860 10008 23866
rect 9956 23802 10008 23808
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9876 23322 9904 23598
rect 9968 23322 9996 23802
rect 10048 23656 10100 23662
rect 10046 23624 10048 23633
rect 10100 23624 10102 23633
rect 10152 23594 10180 23990
rect 10336 23866 10364 24210
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10232 23792 10284 23798
rect 10232 23734 10284 23740
rect 10046 23559 10102 23568
rect 10140 23588 10192 23594
rect 9864 23316 9916 23322
rect 9864 23258 9916 23264
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 9220 23190 9272 23196
rect 9508 23174 9720 23202
rect 9864 23180 9916 23186
rect 9508 23118 9536 23174
rect 9864 23122 9916 23128
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9588 23112 9640 23118
rect 9588 23054 9640 23060
rect 9220 22976 9272 22982
rect 9220 22918 9272 22924
rect 9496 22976 9548 22982
rect 9496 22918 9548 22924
rect 9232 22778 9260 22918
rect 9220 22772 9272 22778
rect 9220 22714 9272 22720
rect 9508 22574 9536 22918
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9508 22234 9536 22510
rect 9600 22506 9628 23054
rect 9772 23044 9824 23050
rect 9692 23004 9772 23032
rect 9588 22500 9640 22506
rect 9588 22442 9640 22448
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9128 21412 9180 21418
rect 9128 21354 9180 21360
rect 9508 20534 9536 21966
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9600 21146 9628 21830
rect 9692 21690 9720 23004
rect 9772 22986 9824 22992
rect 9876 22778 9904 23122
rect 9968 22930 9996 23258
rect 10060 23032 10088 23559
rect 10140 23530 10192 23536
rect 10152 23254 10180 23530
rect 10244 23254 10272 23734
rect 10428 23662 10456 25094
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 10520 24274 10548 24686
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10520 23730 10548 24210
rect 10508 23724 10560 23730
rect 10508 23666 10560 23672
rect 10416 23656 10468 23662
rect 10416 23598 10468 23604
rect 10140 23248 10192 23254
rect 10140 23190 10192 23196
rect 10232 23248 10284 23254
rect 10232 23190 10284 23196
rect 10060 23004 10272 23032
rect 9968 22902 10180 22930
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 9784 22234 9812 22510
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9772 22228 9824 22234
rect 9772 22170 9824 22176
rect 9680 21684 9732 21690
rect 9680 21626 9732 21632
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 9692 20806 9720 21626
rect 9862 21584 9918 21593
rect 9862 21519 9864 21528
rect 9916 21519 9918 21528
rect 9864 21490 9916 21496
rect 9772 21412 9824 21418
rect 9772 21354 9824 21360
rect 9680 20800 9732 20806
rect 9680 20742 9732 20748
rect 9692 20534 9720 20742
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9036 19848 9088 19854
rect 9034 19816 9036 19825
rect 9088 19816 9090 19825
rect 9034 19751 9090 19760
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 9140 18970 9168 19246
rect 9128 18964 9180 18970
rect 9128 18906 9180 18912
rect 9416 18766 9444 20198
rect 9508 19990 9536 20470
rect 9496 19984 9548 19990
rect 9496 19926 9548 19932
rect 9784 19378 9812 21354
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9876 20602 9904 20946
rect 9968 20942 9996 22374
rect 10152 21486 10180 22902
rect 10244 22166 10272 23004
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10232 22160 10284 22166
rect 10232 22102 10284 22108
rect 10336 22098 10364 22714
rect 10324 22092 10376 22098
rect 10324 22034 10376 22040
rect 10324 21888 10376 21894
rect 10324 21830 10376 21836
rect 10140 21480 10192 21486
rect 10140 21422 10192 21428
rect 10152 20942 10180 21422
rect 9956 20936 10008 20942
rect 10140 20936 10192 20942
rect 9956 20878 10008 20884
rect 10046 20904 10102 20913
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9968 20398 9996 20878
rect 10140 20878 10192 20884
rect 10232 20936 10284 20942
rect 10232 20878 10284 20884
rect 10046 20839 10102 20848
rect 10060 20466 10088 20839
rect 10244 20602 10272 20878
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 9956 20392 10008 20398
rect 9956 20334 10008 20340
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9968 19310 9996 20334
rect 10048 20324 10100 20330
rect 10048 20266 10100 20272
rect 10060 19786 10088 20266
rect 10336 19922 10364 21830
rect 10428 20330 10456 23598
rect 10612 23526 10640 24754
rect 11072 24410 11100 25774
rect 11348 25650 11376 26998
rect 11440 26586 11468 27066
rect 11532 27062 11560 27270
rect 11520 27056 11572 27062
rect 11520 26998 11572 27004
rect 11428 26580 11480 26586
rect 11428 26522 11480 26528
rect 11716 26450 11744 27814
rect 11992 27606 12020 28086
rect 12636 27674 12664 28358
rect 12912 27946 12940 29174
rect 13082 29135 13138 29144
rect 12992 28960 13044 28966
rect 12992 28902 13044 28908
rect 13004 28218 13032 28902
rect 13176 28416 13228 28422
rect 13176 28358 13228 28364
rect 13188 28218 13216 28358
rect 12992 28212 13044 28218
rect 12992 28154 13044 28160
rect 13176 28212 13228 28218
rect 13176 28154 13228 28160
rect 13280 28014 13308 29260
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13372 28082 13400 28358
rect 13360 28076 13412 28082
rect 13360 28018 13412 28024
rect 13268 28008 13320 28014
rect 13268 27950 13320 27956
rect 12900 27940 12952 27946
rect 12900 27882 12952 27888
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 11796 27532 11848 27538
rect 11796 27474 11848 27480
rect 12164 27532 12216 27538
rect 12164 27474 12216 27480
rect 11808 26994 11836 27474
rect 11796 26988 11848 26994
rect 11796 26930 11848 26936
rect 11704 26444 11756 26450
rect 11704 26386 11756 26392
rect 11348 25622 11468 25650
rect 11336 25492 11388 25498
rect 11336 25434 11388 25440
rect 11348 24750 11376 25434
rect 11440 25430 11468 25622
rect 11428 25424 11480 25430
rect 11428 25366 11480 25372
rect 11440 24954 11468 25366
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11624 24857 11652 25094
rect 11610 24848 11666 24857
rect 11610 24783 11666 24792
rect 11716 24750 11744 26386
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11520 24744 11572 24750
rect 11520 24686 11572 24692
rect 11704 24744 11756 24750
rect 11704 24686 11756 24692
rect 11428 24676 11480 24682
rect 11428 24618 11480 24624
rect 11060 24404 11112 24410
rect 11060 24346 11112 24352
rect 11440 24342 11468 24618
rect 11428 24336 11480 24342
rect 11428 24278 11480 24284
rect 11532 24274 11560 24686
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 11612 24064 11664 24070
rect 11612 24006 11664 24012
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10612 23186 10640 23462
rect 10600 23180 10652 23186
rect 10600 23122 10652 23128
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10520 21690 10548 21966
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10612 21554 10640 23122
rect 10888 22574 10916 24006
rect 11624 23866 11652 24006
rect 11060 23860 11112 23866
rect 11060 23802 11112 23808
rect 11612 23860 11664 23866
rect 11612 23802 11664 23808
rect 11072 23050 11100 23802
rect 11152 23792 11204 23798
rect 11152 23734 11204 23740
rect 10968 23044 11020 23050
rect 10968 22986 11020 22992
rect 11060 23044 11112 23050
rect 11060 22986 11112 22992
rect 10980 22710 11008 22986
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 10876 22568 10928 22574
rect 10876 22510 10928 22516
rect 11164 22250 11192 23734
rect 11716 23662 11744 24006
rect 11808 23662 11836 26930
rect 11888 26784 11940 26790
rect 11888 26726 11940 26732
rect 11980 26784 12032 26790
rect 11980 26726 12032 26732
rect 11900 26586 11928 26726
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11888 26308 11940 26314
rect 11888 26250 11940 26256
rect 11900 24342 11928 26250
rect 11992 25770 12020 26726
rect 11980 25764 12032 25770
rect 11980 25706 12032 25712
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 12084 25362 12112 25638
rect 12176 25498 12204 27474
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12452 26450 12480 26862
rect 12636 26450 12664 27066
rect 13096 26994 13124 27814
rect 13084 26988 13136 26994
rect 13084 26930 13136 26936
rect 13464 26874 13492 31726
rect 14016 30274 14044 32914
rect 14108 32230 14136 32914
rect 14200 32230 14228 33102
rect 15016 33108 15068 33114
rect 15016 33050 15068 33056
rect 15488 32978 15516 33272
rect 14832 32972 14884 32978
rect 14832 32914 14884 32920
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 15476 32972 15528 32978
rect 15476 32914 15528 32920
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 14280 32768 14332 32774
rect 14280 32710 14332 32716
rect 14292 32298 14320 32710
rect 14439 32668 14747 32677
rect 14439 32666 14445 32668
rect 14501 32666 14525 32668
rect 14581 32666 14605 32668
rect 14661 32666 14685 32668
rect 14741 32666 14747 32668
rect 14501 32614 14503 32666
rect 14683 32614 14685 32666
rect 14439 32612 14445 32614
rect 14501 32612 14525 32614
rect 14581 32612 14605 32614
rect 14661 32612 14685 32614
rect 14741 32612 14747 32614
rect 14439 32603 14747 32612
rect 14844 32502 14872 32914
rect 14924 32836 14976 32842
rect 14924 32778 14976 32784
rect 14832 32496 14884 32502
rect 14832 32438 14884 32444
rect 14936 32366 14964 32778
rect 15016 32768 15068 32774
rect 15016 32710 15068 32716
rect 15028 32473 15056 32710
rect 15014 32464 15070 32473
rect 15014 32399 15070 32408
rect 14372 32360 14424 32366
rect 14372 32302 14424 32308
rect 14832 32360 14884 32366
rect 14832 32302 14884 32308
rect 14924 32360 14976 32366
rect 15120 32348 15148 32914
rect 15580 32881 15608 32914
rect 15566 32872 15622 32881
rect 15566 32807 15622 32816
rect 15568 32496 15620 32502
rect 15568 32438 15620 32444
rect 14924 32302 14976 32308
rect 15028 32320 15148 32348
rect 14280 32292 14332 32298
rect 14280 32234 14332 32240
rect 14096 32224 14148 32230
rect 14096 32166 14148 32172
rect 14188 32224 14240 32230
rect 14188 32166 14240 32172
rect 14108 31958 14136 32166
rect 14096 31952 14148 31958
rect 14096 31894 14148 31900
rect 14200 30802 14228 32166
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14188 30796 14240 30802
rect 14188 30738 14240 30744
rect 14188 30592 14240 30598
rect 14188 30534 14240 30540
rect 14200 30394 14228 30534
rect 14188 30388 14240 30394
rect 14188 30330 14240 30336
rect 14016 30246 14228 30274
rect 14096 30116 14148 30122
rect 14096 30058 14148 30064
rect 14108 29850 14136 30058
rect 13544 29844 13596 29850
rect 13544 29786 13596 29792
rect 14096 29844 14148 29850
rect 14096 29786 14148 29792
rect 13556 28014 13584 29786
rect 13912 29708 13964 29714
rect 13912 29650 13964 29656
rect 13820 29572 13872 29578
rect 13820 29514 13872 29520
rect 13832 29288 13860 29514
rect 13740 29260 13860 29288
rect 13740 29186 13768 29260
rect 13648 29170 13768 29186
rect 13648 29164 13780 29170
rect 13648 29158 13728 29164
rect 13648 28762 13676 29158
rect 13728 29106 13780 29112
rect 13728 29028 13780 29034
rect 13728 28970 13780 28976
rect 13636 28756 13688 28762
rect 13636 28698 13688 28704
rect 13636 28620 13688 28626
rect 13636 28562 13688 28568
rect 13648 28082 13676 28562
rect 13636 28076 13688 28082
rect 13636 28018 13688 28024
rect 13544 28008 13596 28014
rect 13544 27950 13596 27956
rect 13188 26846 13492 26874
rect 13648 26858 13676 28018
rect 13636 26852 13688 26858
rect 12716 26784 12768 26790
rect 12716 26726 12768 26732
rect 12440 26444 12492 26450
rect 12440 26386 12492 26392
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12636 26042 12664 26386
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12164 25492 12216 25498
rect 12164 25434 12216 25440
rect 12256 25424 12308 25430
rect 12256 25366 12308 25372
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 12084 23662 12112 25298
rect 12268 25226 12296 25366
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 12440 25220 12492 25226
rect 12440 25162 12492 25168
rect 12348 24200 12400 24206
rect 12348 24142 12400 24148
rect 12164 24064 12216 24070
rect 12164 24006 12216 24012
rect 11704 23656 11756 23662
rect 11704 23598 11756 23604
rect 11796 23656 11848 23662
rect 11796 23598 11848 23604
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 12072 23656 12124 23662
rect 12072 23598 12124 23604
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11610 23216 11666 23225
rect 11336 23180 11388 23186
rect 11610 23151 11666 23160
rect 11336 23122 11388 23128
rect 11244 22568 11296 22574
rect 11244 22510 11296 22516
rect 10980 22222 11192 22250
rect 10600 21548 10652 21554
rect 10600 21490 10652 21496
rect 10980 21298 11008 22222
rect 11060 22160 11112 22166
rect 11060 22102 11112 22108
rect 11072 21876 11100 22102
rect 11152 21888 11204 21894
rect 11072 21848 11152 21876
rect 11152 21830 11204 21836
rect 10704 21270 11008 21298
rect 11060 21344 11112 21350
rect 11060 21286 11112 21292
rect 10704 20466 10732 21270
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10796 20602 10824 20878
rect 10784 20596 10836 20602
rect 10784 20538 10836 20544
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10506 20360 10562 20369
rect 10416 20324 10468 20330
rect 10796 20346 10824 20538
rect 10888 20466 10916 21082
rect 10980 21010 11008 21270
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10980 20534 11008 20810
rect 10968 20528 11020 20534
rect 10968 20470 11020 20476
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 10506 20295 10562 20304
rect 10612 20318 10824 20346
rect 10416 20266 10468 20272
rect 10428 20058 10456 20266
rect 10416 20052 10468 20058
rect 10416 19994 10468 20000
rect 10520 19922 10548 20295
rect 10612 20262 10640 20318
rect 10600 20256 10652 20262
rect 10876 20256 10928 20262
rect 10600 20198 10652 20204
rect 10796 20204 10876 20210
rect 10796 20198 10928 20204
rect 10796 20182 10916 20198
rect 10324 19916 10376 19922
rect 10324 19858 10376 19864
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 10796 19854 10824 20182
rect 10874 20088 10930 20097
rect 10874 20023 10930 20032
rect 10888 19922 10916 20023
rect 10980 19922 11008 20470
rect 11072 19961 11100 21286
rect 11058 19952 11114 19961
rect 10876 19916 10928 19922
rect 10876 19858 10928 19864
rect 10968 19916 11020 19922
rect 11058 19887 11114 19896
rect 10968 19858 11020 19864
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10048 19780 10100 19786
rect 10048 19722 10100 19728
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 10704 19553 10732 19654
rect 10690 19544 10746 19553
rect 10690 19479 10746 19488
rect 10796 19378 10824 19790
rect 10876 19780 10928 19786
rect 10876 19722 10928 19728
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9508 18970 9536 19178
rect 10784 19168 10836 19174
rect 10784 19110 10836 19116
rect 9954 19000 10010 19009
rect 9496 18964 9548 18970
rect 9954 18935 10010 18944
rect 9496 18906 9548 18912
rect 9968 18902 9996 18935
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9680 18624 9732 18630
rect 9680 18566 9732 18572
rect 10600 18624 10652 18630
rect 10600 18566 10652 18572
rect 8666 18255 8722 18264
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 16658 8708 16934
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8312 14278 8340 15098
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8220 13870 8248 14214
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8128 13654 8248 13682
rect 7944 13530 8064 13546
rect 7932 13524 8064 13530
rect 7984 13518 8064 13524
rect 7932 13466 7984 13472
rect 8220 13394 8248 13654
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8024 13320 8076 13326
rect 8312 13274 8340 14214
rect 8496 13462 8524 16594
rect 8864 15502 8892 18226
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9140 17882 9168 18022
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9588 17808 9640 17814
rect 9588 17750 9640 17756
rect 9600 17338 9628 17750
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9692 17134 9720 18566
rect 10612 18290 10640 18566
rect 10796 18290 10824 19110
rect 10888 18902 10916 19722
rect 10980 19514 11008 19858
rect 10968 19508 11020 19514
rect 10968 19450 11020 19456
rect 10876 18896 10928 18902
rect 10876 18838 10928 18844
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10784 18284 10836 18290
rect 10784 18226 10836 18232
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 10876 18080 10928 18086
rect 10876 18022 10928 18028
rect 9784 17542 9812 18022
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 9324 16794 9352 17070
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 9312 16788 9364 16794
rect 9312 16730 9364 16736
rect 9128 16584 9180 16590
rect 9128 16526 9180 16532
rect 9140 15706 9168 16526
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9692 15706 9720 15914
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9784 15570 9812 15846
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8680 14074 8708 14894
rect 8760 14884 8812 14890
rect 8760 14826 8812 14832
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8668 13864 8720 13870
rect 8668 13806 8720 13812
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8024 13262 8076 13268
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7852 12442 7880 12718
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 7656 11280 7708 11286
rect 7656 11222 7708 11228
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7656 11008 7708 11014
rect 7656 10950 7708 10956
rect 7668 9586 7696 10950
rect 7760 9994 7788 11222
rect 8036 10724 8064 13262
rect 8220 13246 8340 13274
rect 8116 13184 8168 13190
rect 8116 13126 8168 13132
rect 8128 12782 8156 13126
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 8220 12306 8248 13246
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8588 12782 8616 12922
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11626 8156 12038
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 8312 11354 8340 12650
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8576 12640 8628 12646
rect 8576 12582 8628 12588
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8404 11898 8432 12038
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8116 10736 8168 10742
rect 8036 10696 8116 10724
rect 8116 10678 8168 10684
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8220 10266 8248 10474
rect 8312 10266 8340 10950
rect 8404 10674 8432 11834
rect 8496 11626 8524 12582
rect 8588 12374 8616 12582
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8404 10266 8432 10610
rect 8484 10464 8536 10470
rect 8484 10406 8536 10412
rect 8208 10260 8260 10266
rect 8208 10202 8260 10208
rect 8300 10260 8352 10266
rect 8300 10202 8352 10208
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 7210 9276 7518 9285
rect 7210 9274 7216 9276
rect 7272 9274 7296 9276
rect 7352 9274 7376 9276
rect 7432 9274 7456 9276
rect 7512 9274 7518 9276
rect 7272 9222 7274 9274
rect 7454 9222 7456 9274
rect 7210 9220 7216 9222
rect 7272 9220 7296 9222
rect 7352 9220 7376 9222
rect 7432 9220 7456 9222
rect 7512 9220 7518 9222
rect 7210 9211 7518 9220
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6550 8732 6858 8741
rect 6550 8730 6556 8732
rect 6612 8730 6636 8732
rect 6692 8730 6716 8732
rect 6772 8730 6796 8732
rect 6852 8730 6858 8732
rect 6612 8678 6614 8730
rect 6794 8678 6796 8730
rect 6550 8676 6556 8678
rect 6612 8676 6636 8678
rect 6692 8676 6716 8678
rect 6772 8676 6796 8678
rect 6852 8676 6858 8678
rect 6550 8667 6858 8676
rect 7024 8650 7052 9114
rect 8036 8838 8064 9454
rect 8220 9042 8248 9998
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 7024 8634 7144 8650
rect 7024 8628 7156 8634
rect 7024 8622 7104 8628
rect 7104 8570 7156 8576
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6460 7948 6512 7954
rect 6460 7890 6512 7896
rect 6564 7834 6592 8230
rect 7210 8188 7518 8197
rect 7210 8186 7216 8188
rect 7272 8186 7296 8188
rect 7352 8186 7376 8188
rect 7432 8186 7456 8188
rect 7512 8186 7518 8188
rect 7272 8134 7274 8186
rect 7454 8134 7456 8186
rect 7210 8132 7216 8134
rect 7272 8132 7296 8134
rect 7352 8132 7376 8134
rect 7432 8132 7456 8134
rect 7512 8132 7518 8134
rect 7210 8123 7518 8132
rect 7668 8090 7696 8298
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 6472 7806 6592 7834
rect 6472 7410 6500 7806
rect 6550 7644 6858 7653
rect 6550 7642 6556 7644
rect 6612 7642 6636 7644
rect 6692 7642 6716 7644
rect 6772 7642 6796 7644
rect 6852 7642 6858 7644
rect 6612 7590 6614 7642
rect 6794 7590 6796 7642
rect 6550 7588 6556 7590
rect 6612 7588 6636 7590
rect 6692 7588 6716 7590
rect 6772 7588 6796 7590
rect 6852 7588 6858 7590
rect 6550 7579 6858 7588
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6552 7200 6604 7206
rect 6552 7142 6604 7148
rect 6564 6746 6592 7142
rect 7210 7100 7518 7109
rect 7210 7098 7216 7100
rect 7272 7098 7296 7100
rect 7352 7098 7376 7100
rect 7432 7098 7456 7100
rect 7512 7098 7518 7100
rect 7272 7046 7274 7098
rect 7454 7046 7456 7098
rect 7210 7044 7216 7046
rect 7272 7044 7296 7046
rect 7352 7044 7376 7046
rect 7432 7044 7456 7046
rect 7512 7044 7518 7046
rect 7210 7035 7518 7044
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 6472 6718 6592 6746
rect 6472 6390 6500 6718
rect 6550 6556 6858 6565
rect 6550 6554 6556 6556
rect 6612 6554 6636 6556
rect 6692 6554 6716 6556
rect 6772 6554 6796 6556
rect 6852 6554 6858 6556
rect 6612 6502 6614 6554
rect 6794 6502 6796 6554
rect 6550 6500 6556 6502
rect 6612 6500 6636 6502
rect 6692 6500 6716 6502
rect 6772 6500 6796 6502
rect 6852 6500 6858 6502
rect 6550 6491 6858 6500
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 7116 5914 7144 6870
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7484 6390 7512 6734
rect 7472 6384 7524 6390
rect 7472 6326 7524 6332
rect 7852 6322 7880 6734
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 7210 6012 7518 6021
rect 7210 6010 7216 6012
rect 7272 6010 7296 6012
rect 7352 6010 7376 6012
rect 7432 6010 7456 6012
rect 7512 6010 7518 6012
rect 7272 5958 7274 6010
rect 7454 5958 7456 6010
rect 7210 5956 7216 5958
rect 7272 5956 7296 5958
rect 7352 5956 7376 5958
rect 7432 5956 7456 5958
rect 7512 5956 7518 5958
rect 7210 5947 7518 5956
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6472 5098 6500 5782
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6550 5468 6858 5477
rect 6550 5466 6556 5468
rect 6612 5466 6636 5468
rect 6692 5466 6716 5468
rect 6772 5466 6796 5468
rect 6852 5466 6858 5468
rect 6612 5414 6614 5466
rect 6794 5414 6796 5466
rect 6550 5412 6556 5414
rect 6612 5412 6636 5414
rect 6692 5412 6716 5414
rect 6772 5412 6796 5414
rect 6852 5412 6858 5414
rect 6550 5403 6858 5412
rect 6460 5092 6512 5098
rect 6460 5034 6512 5040
rect 6932 4826 6960 5646
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5166 7328 5510
rect 7668 5166 7696 5714
rect 7852 5234 7880 6258
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7944 5914 7972 6122
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7656 5160 7708 5166
rect 7656 5102 7708 5108
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7210 4924 7518 4933
rect 7210 4922 7216 4924
rect 7272 4922 7296 4924
rect 7352 4922 7376 4924
rect 7432 4922 7456 4924
rect 7512 4922 7518 4924
rect 7272 4870 7274 4922
rect 7454 4870 7456 4922
rect 7210 4868 7216 4870
rect 7272 4868 7296 4870
rect 7352 4868 7376 4870
rect 7432 4868 7456 4870
rect 7512 4868 7518 4870
rect 7210 4859 7518 4868
rect 6196 4820 6328 4826
rect 6196 4814 6276 4820
rect 6276 4762 6328 4768
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5816 4684 5868 4690
rect 5816 4626 5868 4632
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5644 4214 5672 4626
rect 5828 4570 5856 4626
rect 6104 4570 6132 4694
rect 5828 4542 6132 4570
rect 6104 4282 6132 4542
rect 6288 4282 6316 4762
rect 7760 4758 7788 4966
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 6276 4276 6328 4282
rect 6276 4218 6328 4224
rect 5632 4208 5684 4214
rect 5632 4150 5684 4156
rect 6380 4146 6408 4558
rect 7944 4554 7972 5170
rect 7932 4548 7984 4554
rect 7932 4490 7984 4496
rect 6550 4380 6858 4389
rect 6550 4378 6556 4380
rect 6612 4378 6636 4380
rect 6692 4378 6716 4380
rect 6772 4378 6796 4380
rect 6852 4378 6858 4380
rect 6612 4326 6614 4378
rect 6794 4326 6796 4378
rect 6550 4324 6556 4326
rect 6612 4324 6636 4326
rect 6692 4324 6716 4326
rect 6772 4324 6796 4326
rect 6852 4324 6858 4326
rect 6550 4315 6858 4324
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 7210 3836 7518 3845
rect 7210 3834 7216 3836
rect 7272 3834 7296 3836
rect 7352 3834 7376 3836
rect 7432 3834 7456 3836
rect 7512 3834 7518 3836
rect 7272 3782 7274 3834
rect 7454 3782 7456 3834
rect 7210 3780 7216 3782
rect 7272 3780 7296 3782
rect 7352 3780 7376 3782
rect 7432 3780 7456 3782
rect 7512 3780 7518 3782
rect 7210 3771 7518 3780
rect 6550 3292 6858 3301
rect 6550 3290 6556 3292
rect 6612 3290 6636 3292
rect 6692 3290 6716 3292
rect 6772 3290 6796 3292
rect 6852 3290 6858 3292
rect 6612 3238 6614 3290
rect 6794 3238 6796 3290
rect 6550 3236 6556 3238
rect 6612 3236 6636 3238
rect 6692 3236 6716 3238
rect 6772 3236 6796 3238
rect 6852 3236 6858 3238
rect 6550 3227 6858 3236
rect 5722 3088 5778 3097
rect 5722 3023 5724 3032
rect 5776 3023 5778 3032
rect 7748 3052 7800 3058
rect 5724 2994 5776 3000
rect 7748 2994 7800 3000
rect 5264 2984 5316 2990
rect 5264 2926 5316 2932
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6656 1442 6684 2858
rect 7210 2748 7518 2757
rect 7210 2746 7216 2748
rect 7272 2746 7296 2748
rect 7352 2746 7376 2748
rect 7432 2746 7456 2748
rect 7512 2746 7518 2748
rect 7272 2694 7274 2746
rect 7454 2694 7456 2746
rect 7210 2692 7216 2694
rect 7272 2692 7296 2694
rect 7352 2692 7376 2694
rect 7432 2692 7456 2694
rect 7512 2692 7518 2694
rect 7210 2683 7518 2692
rect 6472 1414 6684 1442
rect 6472 800 6500 1414
rect 7760 800 7788 2994
rect 8036 2990 8064 8774
rect 8220 7818 8248 8978
rect 8312 8634 8340 10202
rect 8496 10198 8524 10406
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8680 10130 8708 13806
rect 8772 10606 8800 14826
rect 9048 14822 9076 15438
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8864 13802 8892 14554
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8956 12986 8984 13942
rect 9048 13190 9076 14758
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9140 14074 9168 14350
rect 9784 14074 9812 14758
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9876 13734 9904 16934
rect 10140 15972 10192 15978
rect 10140 15914 10192 15920
rect 10152 15706 10180 15914
rect 10244 15910 10272 16934
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 9956 15020 10008 15026
rect 9956 14962 10008 14968
rect 9968 13802 9996 14962
rect 10140 14952 10192 14958
rect 10140 14894 10192 14900
rect 10152 14618 10180 14894
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10048 14544 10100 14550
rect 10048 14486 10100 14492
rect 10060 14074 10088 14486
rect 10244 14414 10272 15846
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10048 13864 10100 13870
rect 10048 13806 10100 13812
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9864 13728 9916 13734
rect 9864 13670 9916 13676
rect 9876 13530 9904 13670
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 9864 13524 9916 13530
rect 9864 13466 9916 13472
rect 9036 13184 9088 13190
rect 9036 13126 9088 13132
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8956 11898 8984 12922
rect 9048 12714 9076 13126
rect 9140 12782 9168 13466
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9140 10606 9168 12718
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9784 11898 9812 12242
rect 9772 11892 9824 11898
rect 9772 11834 9824 11840
rect 9968 11354 9996 13738
rect 10060 11694 10088 13806
rect 10244 12306 10272 14350
rect 10336 13870 10364 15506
rect 10428 15502 10456 17070
rect 10520 16046 10548 17478
rect 10888 17202 10916 18022
rect 11072 17542 11100 19887
rect 11164 19310 11192 21830
rect 11256 20482 11284 22510
rect 11348 22438 11376 23122
rect 11624 22982 11652 23151
rect 11612 22976 11664 22982
rect 11612 22918 11664 22924
rect 11428 22568 11480 22574
rect 11428 22510 11480 22516
rect 11612 22568 11664 22574
rect 11612 22510 11664 22516
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11348 21418 11376 22374
rect 11336 21412 11388 21418
rect 11336 21354 11388 21360
rect 11336 21004 11388 21010
rect 11336 20946 11388 20952
rect 11348 20602 11376 20946
rect 11440 20788 11468 22510
rect 11520 22092 11572 22098
rect 11520 22034 11572 22040
rect 11532 21894 11560 22034
rect 11520 21888 11572 21894
rect 11520 21830 11572 21836
rect 11624 21486 11652 22510
rect 11808 22438 11836 23462
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11900 22710 11928 23122
rect 11888 22704 11940 22710
rect 11888 22646 11940 22652
rect 11992 22642 12020 23598
rect 12176 23050 12204 24006
rect 12360 23526 12388 24142
rect 12452 23730 12480 25162
rect 12728 24614 12756 26726
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12622 23624 12678 23633
rect 12622 23559 12678 23568
rect 12900 23588 12952 23594
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12164 23044 12216 23050
rect 12164 22986 12216 22992
rect 11980 22636 12032 22642
rect 11980 22578 12032 22584
rect 11796 22432 11848 22438
rect 11796 22374 11848 22380
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11716 21729 11744 21830
rect 11702 21720 11758 21729
rect 11702 21655 11758 21664
rect 11612 21480 11664 21486
rect 11532 21440 11612 21468
rect 11532 21078 11560 21440
rect 11612 21422 11664 21428
rect 11704 21480 11756 21486
rect 11704 21422 11756 21428
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11624 21078 11652 21286
rect 11520 21072 11572 21078
rect 11520 21014 11572 21020
rect 11612 21072 11664 21078
rect 11612 21014 11664 21020
rect 11520 20936 11572 20942
rect 11518 20904 11520 20913
rect 11572 20904 11574 20913
rect 11518 20839 11574 20848
rect 11520 20800 11572 20806
rect 11440 20760 11520 20788
rect 11520 20742 11572 20748
rect 11336 20596 11388 20602
rect 11336 20538 11388 20544
rect 11256 20454 11376 20482
rect 11348 19825 11376 20454
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 11440 20058 11468 20334
rect 11532 20058 11560 20742
rect 11716 20466 11744 21422
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11808 20346 11836 22374
rect 11992 21010 12020 22578
rect 12176 22234 12204 22986
rect 12164 22228 12216 22234
rect 12360 22216 12388 23462
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22438 12480 23122
rect 12636 22982 12664 23559
rect 12900 23530 12952 23536
rect 12716 23180 12768 23186
rect 12716 23122 12768 23128
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12728 22658 12756 23122
rect 12636 22630 12756 22658
rect 12636 22574 12664 22630
rect 12624 22568 12676 22574
rect 12624 22510 12676 22516
rect 12716 22568 12768 22574
rect 12716 22510 12768 22516
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12360 22188 12480 22216
rect 12164 22170 12216 22176
rect 12176 22012 12204 22170
rect 12348 22092 12400 22098
rect 12348 22034 12400 22040
rect 12256 22024 12308 22030
rect 12176 21984 12256 22012
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 12084 21554 12112 21830
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 12176 20890 12204 21984
rect 12256 21966 12308 21972
rect 12360 21690 12388 22034
rect 12348 21684 12400 21690
rect 12348 21626 12400 21632
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12268 21350 12296 21558
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12452 21010 12480 22188
rect 12728 22094 12756 22510
rect 12636 22066 12756 22094
rect 12912 22094 12940 23530
rect 13084 22976 13136 22982
rect 13084 22918 13136 22924
rect 13096 22642 13124 22918
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 12912 22066 13124 22094
rect 12636 22030 12664 22066
rect 12624 22024 12676 22030
rect 12624 21966 12676 21972
rect 12636 21554 12664 21966
rect 12624 21548 12676 21554
rect 12624 21490 12676 21496
rect 12714 21040 12770 21049
rect 12256 21004 12308 21010
rect 12256 20946 12308 20952
rect 12440 21004 12492 21010
rect 12770 20998 12848 21026
rect 12714 20975 12770 20984
rect 12440 20946 12492 20952
rect 11992 20862 12204 20890
rect 11886 20496 11942 20505
rect 11886 20431 11942 20440
rect 11624 20318 11836 20346
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11334 19816 11390 19825
rect 11334 19751 11390 19760
rect 11242 19544 11298 19553
rect 11348 19514 11376 19751
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11242 19479 11298 19488
rect 11336 19508 11388 19514
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 11256 19258 11284 19479
rect 11336 19450 11388 19456
rect 11256 19242 11376 19258
rect 11256 19236 11388 19242
rect 11256 19230 11336 19236
rect 11336 19178 11388 19184
rect 11440 18630 11468 19654
rect 11624 19310 11652 20318
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11520 19236 11572 19242
rect 11520 19178 11572 19184
rect 11532 18902 11560 19178
rect 11520 18896 11572 18902
rect 11520 18838 11572 18844
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11060 17536 11112 17542
rect 11060 17478 11112 17484
rect 10876 17196 10928 17202
rect 10876 17138 10928 17144
rect 11072 16726 11100 17478
rect 11716 16946 11744 19858
rect 11900 18970 11928 20431
rect 11992 19378 12020 20862
rect 12268 20380 12296 20946
rect 12348 20460 12400 20466
rect 12348 20402 12400 20408
rect 12176 20352 12296 20380
rect 12072 20256 12124 20262
rect 12072 20198 12124 20204
rect 12084 19990 12112 20198
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 12176 19938 12204 20352
rect 12176 19910 12296 19938
rect 12360 19922 12388 20402
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12176 19258 12204 19790
rect 12084 19230 12204 19258
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11808 18426 11836 18566
rect 11796 18420 11848 18426
rect 11796 18362 11848 18368
rect 11624 16918 11744 16946
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11072 16182 11100 16662
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15162 10456 15438
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10428 13802 10456 15098
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10416 13796 10468 13802
rect 10416 13738 10468 13744
rect 10416 13524 10468 13530
rect 10336 13484 10416 13512
rect 10232 12300 10284 12306
rect 10232 12242 10284 12248
rect 10336 12186 10364 13484
rect 10416 13466 10468 13472
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10244 12158 10364 12186
rect 10140 12096 10192 12102
rect 10140 12038 10192 12044
rect 10152 11830 10180 12038
rect 10140 11824 10192 11830
rect 10140 11766 10192 11772
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9680 11008 9732 11014
rect 9680 10950 9732 10956
rect 9692 10674 9720 10950
rect 9876 10742 9904 11222
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 8772 10266 8800 10542
rect 8852 10532 8904 10538
rect 8852 10474 8904 10480
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8588 9654 8616 9862
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 7812 8260 7818
rect 8208 7754 8260 7760
rect 8220 5846 8248 7754
rect 8312 7342 8340 8570
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8312 6458 8340 7278
rect 8404 6866 8432 9522
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8496 8090 8524 8978
rect 8484 8084 8536 8090
rect 8484 8026 8536 8032
rect 8588 7750 8616 9590
rect 8680 7954 8708 10066
rect 8864 10062 8892 10474
rect 9140 10198 9168 10542
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 9140 8650 9168 10134
rect 9600 10130 9628 10542
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9324 8838 9352 10066
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 9496 8832 9548 8838
rect 9496 8774 9548 8780
rect 9048 8622 9168 8650
rect 8668 7948 8720 7954
rect 8668 7890 8720 7896
rect 8852 7948 8904 7954
rect 8852 7890 8904 7896
rect 8680 7857 8708 7890
rect 8666 7848 8722 7857
rect 8666 7783 8722 7792
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8208 5840 8260 5846
rect 8208 5782 8260 5788
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 4486 8340 5170
rect 8404 5098 8432 5850
rect 8588 5794 8616 7686
rect 8680 7206 8708 7783
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8496 5766 8616 5794
rect 8496 5234 8524 5766
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8588 5370 8616 5646
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 5092 8444 5098
rect 8392 5034 8444 5040
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8404 4706 8432 5034
rect 8404 4678 8524 4706
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8404 4146 8432 4490
rect 8496 4282 8524 4678
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8588 4078 8616 5034
rect 8680 5030 8708 5646
rect 8864 5166 8892 7890
rect 9048 7546 9076 8622
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 6322 9076 7142
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 8668 5024 8720 5030
rect 8668 4966 8720 4972
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8680 3602 8708 4966
rect 9048 4146 9076 6258
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 9048 3738 9076 4082
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 9036 2984 9088 2990
rect 9036 2926 9088 2932
rect 9048 800 9076 2926
rect 9140 2922 9168 8434
rect 9220 8288 9272 8294
rect 9220 8230 9272 8236
rect 9232 8090 9260 8230
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9218 7984 9274 7993
rect 9218 7919 9220 7928
rect 9272 7919 9274 7928
rect 9220 7890 9272 7896
rect 9324 7818 9352 8774
rect 9508 8362 9536 8774
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9324 7410 9352 7754
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 9324 5914 9352 7346
rect 9600 6254 9628 9862
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9692 8090 9720 8366
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9784 7970 9812 9046
rect 9968 8974 9996 9318
rect 10244 9178 10272 12158
rect 10324 11144 10376 11150
rect 10324 11086 10376 11092
rect 10336 10810 10364 11086
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10428 9178 10456 13330
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9692 7942 9812 7970
rect 9968 8044 10272 8072
rect 9692 7886 9720 7942
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9692 7206 9720 7822
rect 9968 7750 9996 8044
rect 10048 7948 10100 7954
rect 10048 7890 10100 7896
rect 9956 7744 10008 7750
rect 9956 7686 10008 7692
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9588 6248 9640 6254
rect 9588 6190 9640 6196
rect 9772 6112 9824 6118
rect 9772 6054 9824 6060
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9784 5370 9812 6054
rect 10060 5914 10088 7890
rect 10244 7886 10272 8044
rect 10520 7954 10548 14758
rect 10612 13462 10640 15846
rect 11164 15638 11192 16730
rect 11336 16040 11388 16046
rect 11336 15982 11388 15988
rect 11348 15706 11376 15982
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11152 15632 11204 15638
rect 11152 15574 11204 15580
rect 11520 15428 11572 15434
rect 11520 15370 11572 15376
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11072 15162 11100 15302
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 11164 15026 11192 15302
rect 11336 15088 11388 15094
rect 11336 15030 11388 15036
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10704 14074 10732 14350
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10600 13456 10652 13462
rect 10600 13398 10652 13404
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10876 12640 10928 12646
rect 10876 12582 10928 12588
rect 10612 12238 10640 12582
rect 10784 12368 10836 12374
rect 10888 12322 10916 12582
rect 10836 12316 10916 12322
rect 10784 12310 10916 12316
rect 10796 12294 10916 12310
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10980 11558 11008 14894
rect 11348 12628 11376 15030
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14550 11468 14758
rect 11428 14544 11480 14550
rect 11428 14486 11480 14492
rect 11428 12640 11480 12646
rect 11348 12600 11428 12628
rect 11428 12582 11480 12588
rect 11152 11688 11204 11694
rect 11152 11630 11204 11636
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10796 11218 10824 11494
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10612 10130 10640 11086
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10508 7948 10560 7954
rect 10508 7890 10560 7896
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 10152 6662 10180 7482
rect 10428 7478 10456 7686
rect 10612 7546 10640 10066
rect 10692 9444 10744 9450
rect 10692 9386 10744 9392
rect 10704 9178 10732 9386
rect 10796 9382 10824 11154
rect 10980 10606 11008 11290
rect 11164 11014 11192 11630
rect 11440 11540 11468 12582
rect 11532 11694 11560 15370
rect 11624 13394 11652 16918
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 11992 15706 12020 16662
rect 11980 15700 12032 15706
rect 11980 15642 12032 15648
rect 12084 14890 12112 19230
rect 12164 19168 12216 19174
rect 12164 19110 12216 19116
rect 12176 18970 12204 19110
rect 12268 18970 12296 19910
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12360 19310 12388 19858
rect 12532 19712 12584 19718
rect 12532 19654 12584 19660
rect 12544 19378 12572 19654
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12348 19304 12400 19310
rect 12820 19281 12848 20998
rect 12900 20868 12952 20874
rect 12900 20810 12952 20816
rect 12348 19246 12400 19252
rect 12806 19272 12862 19281
rect 12806 19207 12862 19216
rect 12440 19168 12492 19174
rect 12912 19156 12940 20810
rect 13096 20806 13124 22066
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 12992 20324 13044 20330
rect 12992 20266 13044 20272
rect 13004 20058 13032 20266
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12440 19110 12492 19116
rect 12728 19128 12940 19156
rect 12164 18964 12216 18970
rect 12164 18906 12216 18912
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12452 18766 12480 19110
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 12176 17338 12204 18566
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12268 17338 12296 17614
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12176 16726 12204 17274
rect 12164 16720 12216 16726
rect 12164 16662 12216 16668
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12176 14890 12204 15438
rect 12072 14884 12124 14890
rect 12072 14826 12124 14832
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 11704 13932 11756 13938
rect 11704 13874 11756 13880
rect 11716 13530 11744 13874
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11716 12850 11744 13466
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11612 12640 11664 12646
rect 11612 12582 11664 12588
rect 11624 12306 11652 12582
rect 11612 12300 11664 12306
rect 11612 12242 11664 12248
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11624 11540 11652 11630
rect 11440 11512 11652 11540
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10888 10266 10916 10542
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10888 9926 10916 10202
rect 11164 10062 11192 10950
rect 11348 10810 11376 11086
rect 11612 11076 11664 11082
rect 11612 11018 11664 11024
rect 11520 11008 11572 11014
rect 11520 10950 11572 10956
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 11532 10198 11560 10950
rect 11520 10192 11572 10198
rect 11520 10134 11572 10140
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8566 11560 9046
rect 11520 8560 11572 8566
rect 11520 8502 11572 8508
rect 11624 7954 11652 11018
rect 11716 10538 11744 12786
rect 11980 12776 12032 12782
rect 11808 12724 11980 12730
rect 11808 12718 12032 12724
rect 11808 12702 12020 12718
rect 11808 10674 11836 12702
rect 12084 12594 12112 13262
rect 12176 12714 12204 14826
rect 12360 13870 12388 17614
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12452 12986 12480 13126
rect 12440 12980 12492 12986
rect 12440 12922 12492 12928
rect 12348 12844 12400 12850
rect 12544 12832 12572 14010
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12400 12804 12572 12832
rect 12348 12786 12400 12792
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 11992 12566 12112 12594
rect 11992 12442 12020 12566
rect 12176 12442 12204 12650
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12544 11898 12572 12804
rect 12636 12442 12664 13874
rect 12728 13818 12756 19128
rect 12900 18828 12952 18834
rect 12900 18770 12952 18776
rect 12912 18630 12940 18770
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 12912 17814 12940 18022
rect 12900 17808 12952 17814
rect 12900 17750 12952 17756
rect 12912 17202 12940 17750
rect 13004 17746 13032 18022
rect 13096 17746 13124 18226
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12806 17096 12862 17105
rect 12806 17031 12808 17040
rect 12860 17031 12862 17040
rect 12808 17002 12860 17008
rect 12820 15502 12848 17002
rect 13096 16658 13124 17682
rect 13188 17184 13216 26846
rect 13636 26794 13688 26800
rect 13648 26738 13676 26794
rect 13556 26710 13676 26738
rect 13556 25974 13584 26710
rect 13740 26586 13768 28970
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13832 27878 13860 28426
rect 13924 28422 13952 29650
rect 14004 29572 14056 29578
rect 14004 29514 14056 29520
rect 14016 29102 14044 29514
rect 14108 29306 14136 29786
rect 14096 29300 14148 29306
rect 14096 29242 14148 29248
rect 14108 29170 14136 29242
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14004 29096 14056 29102
rect 14004 29038 14056 29044
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 13820 27872 13872 27878
rect 13820 27814 13872 27820
rect 13924 27606 13952 28358
rect 14016 28014 14044 29038
rect 14108 28218 14136 29106
rect 14096 28212 14148 28218
rect 14096 28154 14148 28160
rect 14004 28008 14056 28014
rect 14004 27950 14056 27956
rect 14004 27872 14056 27878
rect 14004 27814 14056 27820
rect 13912 27600 13964 27606
rect 13912 27542 13964 27548
rect 13820 27328 13872 27334
rect 13820 27270 13872 27276
rect 13832 26994 13860 27270
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13924 26586 13952 27542
rect 14016 27033 14044 27814
rect 14096 27600 14148 27606
rect 14096 27542 14148 27548
rect 14108 27130 14136 27542
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 14002 27024 14058 27033
rect 14002 26959 14058 26968
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13728 26580 13780 26586
rect 13728 26522 13780 26528
rect 13912 26580 13964 26586
rect 13912 26522 13964 26528
rect 13544 25968 13596 25974
rect 13544 25910 13596 25916
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 13268 25764 13320 25770
rect 13268 25706 13320 25712
rect 13280 25498 13308 25706
rect 13464 25498 13492 25842
rect 13648 25838 13676 26522
rect 13740 25838 13768 26522
rect 13924 26314 13952 26522
rect 13912 26308 13964 26314
rect 13912 26250 13964 26256
rect 14016 26194 14044 26959
rect 14108 26586 14136 27066
rect 14200 26874 14228 30246
rect 14292 29850 14320 31826
rect 14384 31754 14412 32302
rect 14844 31958 14872 32302
rect 14832 31952 14884 31958
rect 14832 31894 14884 31900
rect 14372 31748 14424 31754
rect 14372 31690 14424 31696
rect 14924 31680 14976 31686
rect 15028 31668 15056 32320
rect 15099 32124 15407 32133
rect 15099 32122 15105 32124
rect 15161 32122 15185 32124
rect 15241 32122 15265 32124
rect 15321 32122 15345 32124
rect 15401 32122 15407 32124
rect 15161 32070 15163 32122
rect 15343 32070 15345 32122
rect 15099 32068 15105 32070
rect 15161 32068 15185 32070
rect 15241 32068 15265 32070
rect 15321 32068 15345 32070
rect 15401 32068 15407 32070
rect 15099 32059 15407 32068
rect 15476 32020 15528 32026
rect 15476 31962 15528 31968
rect 15384 31952 15436 31958
rect 15384 31894 15436 31900
rect 14976 31640 15056 31668
rect 14924 31622 14976 31628
rect 14439 31580 14747 31589
rect 14439 31578 14445 31580
rect 14501 31578 14525 31580
rect 14581 31578 14605 31580
rect 14661 31578 14685 31580
rect 14741 31578 14747 31580
rect 14501 31526 14503 31578
rect 14683 31526 14685 31578
rect 14439 31524 14445 31526
rect 14501 31524 14525 31526
rect 14581 31524 14605 31526
rect 14661 31524 14685 31526
rect 14741 31524 14747 31526
rect 14439 31515 14747 31524
rect 14832 30660 14884 30666
rect 14832 30602 14884 30608
rect 14439 30492 14747 30501
rect 14439 30490 14445 30492
rect 14501 30490 14525 30492
rect 14581 30490 14605 30492
rect 14661 30490 14685 30492
rect 14741 30490 14747 30492
rect 14501 30438 14503 30490
rect 14683 30438 14685 30490
rect 14439 30436 14445 30438
rect 14501 30436 14525 30438
rect 14581 30436 14605 30438
rect 14661 30436 14685 30438
rect 14741 30436 14747 30438
rect 14439 30427 14747 30436
rect 14844 30274 14872 30602
rect 14752 30246 14872 30274
rect 14280 29844 14332 29850
rect 14280 29786 14332 29792
rect 14752 29510 14780 30246
rect 14832 29776 14884 29782
rect 14832 29718 14884 29724
rect 14740 29504 14792 29510
rect 14740 29446 14792 29452
rect 14439 29404 14747 29413
rect 14439 29402 14445 29404
rect 14501 29402 14525 29404
rect 14581 29402 14605 29404
rect 14661 29402 14685 29404
rect 14741 29402 14747 29404
rect 14501 29350 14503 29402
rect 14683 29350 14685 29402
rect 14439 29348 14445 29350
rect 14501 29348 14525 29350
rect 14581 29348 14605 29350
rect 14661 29348 14685 29350
rect 14741 29348 14747 29350
rect 14439 29339 14747 29348
rect 14844 29170 14872 29718
rect 14648 29164 14700 29170
rect 14832 29164 14884 29170
rect 14700 29124 14780 29152
rect 14648 29106 14700 29112
rect 14372 29028 14424 29034
rect 14372 28970 14424 28976
rect 14280 28756 14332 28762
rect 14280 28698 14332 28704
rect 14292 28014 14320 28698
rect 14384 28490 14412 28970
rect 14752 28626 14780 29124
rect 14832 29106 14884 29112
rect 14844 28762 14872 29106
rect 14936 29034 14964 31622
rect 15396 31482 15424 31894
rect 15488 31482 15516 31962
rect 15580 31958 15608 32438
rect 15936 32292 15988 32298
rect 15936 32234 15988 32240
rect 15660 32224 15712 32230
rect 15660 32166 15712 32172
rect 15568 31952 15620 31958
rect 15568 31894 15620 31900
rect 15672 31770 15700 32166
rect 15948 32026 15976 32234
rect 15936 32020 15988 32026
rect 15936 31962 15988 31968
rect 15752 31816 15804 31822
rect 15672 31764 15752 31770
rect 15804 31764 15884 31770
rect 15672 31742 15884 31764
rect 15384 31476 15436 31482
rect 15384 31418 15436 31424
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 15099 31036 15407 31045
rect 15099 31034 15105 31036
rect 15161 31034 15185 31036
rect 15241 31034 15265 31036
rect 15321 31034 15345 31036
rect 15401 31034 15407 31036
rect 15161 30982 15163 31034
rect 15343 30982 15345 31034
rect 15099 30980 15105 30982
rect 15161 30980 15185 30982
rect 15241 30980 15265 30982
rect 15321 30980 15345 30982
rect 15401 30980 15407 30982
rect 15099 30971 15407 30980
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15120 30394 15148 30670
rect 15108 30388 15160 30394
rect 15108 30330 15160 30336
rect 15660 30252 15712 30258
rect 15660 30194 15712 30200
rect 15099 29948 15407 29957
rect 15099 29946 15105 29948
rect 15161 29946 15185 29948
rect 15241 29946 15265 29948
rect 15321 29946 15345 29948
rect 15401 29946 15407 29948
rect 15161 29894 15163 29946
rect 15343 29894 15345 29946
rect 15099 29892 15105 29894
rect 15161 29892 15185 29894
rect 15241 29892 15265 29894
rect 15321 29892 15345 29894
rect 15401 29892 15407 29894
rect 15099 29883 15407 29892
rect 15016 29708 15068 29714
rect 15016 29650 15068 29656
rect 15476 29708 15528 29714
rect 15476 29650 15528 29656
rect 15028 29306 15056 29650
rect 15016 29300 15068 29306
rect 15016 29242 15068 29248
rect 14924 29028 14976 29034
rect 14924 28970 14976 28976
rect 14832 28756 14884 28762
rect 14832 28698 14884 28704
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14372 28484 14424 28490
rect 14372 28426 14424 28432
rect 14439 28316 14747 28325
rect 14439 28314 14445 28316
rect 14501 28314 14525 28316
rect 14581 28314 14605 28316
rect 14661 28314 14685 28316
rect 14741 28314 14747 28316
rect 14501 28262 14503 28314
rect 14683 28262 14685 28314
rect 14439 28260 14445 28262
rect 14501 28260 14525 28262
rect 14581 28260 14605 28262
rect 14661 28260 14685 28262
rect 14741 28260 14747 28262
rect 14439 28251 14747 28260
rect 14372 28076 14424 28082
rect 14372 28018 14424 28024
rect 14280 28008 14332 28014
rect 14280 27950 14332 27956
rect 14292 27520 14320 27950
rect 14384 27674 14412 28018
rect 14648 27872 14700 27878
rect 14648 27814 14700 27820
rect 14372 27668 14424 27674
rect 14372 27610 14424 27616
rect 14372 27532 14424 27538
rect 14292 27492 14372 27520
rect 14372 27474 14424 27480
rect 14660 27470 14688 27814
rect 14648 27464 14700 27470
rect 14648 27406 14700 27412
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14292 27062 14320 27270
rect 14439 27228 14747 27237
rect 14439 27226 14445 27228
rect 14501 27226 14525 27228
rect 14581 27226 14605 27228
rect 14661 27226 14685 27228
rect 14741 27226 14747 27228
rect 14501 27174 14503 27226
rect 14683 27174 14685 27226
rect 14439 27172 14445 27174
rect 14501 27172 14525 27174
rect 14581 27172 14605 27174
rect 14661 27172 14685 27174
rect 14741 27172 14747 27174
rect 14439 27163 14747 27172
rect 14844 27130 14872 28698
rect 14936 28626 14964 28970
rect 15028 28626 15056 29242
rect 15099 28860 15407 28869
rect 15099 28858 15105 28860
rect 15161 28858 15185 28860
rect 15241 28858 15265 28860
rect 15321 28858 15345 28860
rect 15401 28858 15407 28860
rect 15161 28806 15163 28858
rect 15343 28806 15345 28858
rect 15099 28804 15105 28806
rect 15161 28804 15185 28806
rect 15241 28804 15265 28806
rect 15321 28804 15345 28806
rect 15401 28804 15407 28806
rect 15099 28795 15407 28804
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 15016 28620 15068 28626
rect 15016 28562 15068 28568
rect 14936 27402 14964 28562
rect 15488 28558 15516 29650
rect 15672 29306 15700 30194
rect 15660 29300 15712 29306
rect 15660 29242 15712 29248
rect 15856 29170 15884 31742
rect 16040 31754 16068 33816
rect 16948 33798 17000 33804
rect 16120 32904 16172 32910
rect 16120 32846 16172 32852
rect 16132 32570 16160 32846
rect 16764 32768 16816 32774
rect 16764 32710 16816 32716
rect 16776 32570 16804 32710
rect 16120 32564 16172 32570
rect 16120 32506 16172 32512
rect 16764 32564 16816 32570
rect 16764 32506 16816 32512
rect 16580 32428 16632 32434
rect 16580 32370 16632 32376
rect 16592 31822 16620 32370
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16040 31726 16160 31754
rect 16028 30184 16080 30190
rect 16028 30126 16080 30132
rect 16040 29850 16068 30126
rect 16028 29844 16080 29850
rect 16028 29786 16080 29792
rect 15844 29164 15896 29170
rect 15844 29106 15896 29112
rect 15844 28620 15896 28626
rect 15844 28562 15896 28568
rect 15476 28552 15528 28558
rect 15476 28494 15528 28500
rect 15752 28212 15804 28218
rect 15752 28154 15804 28160
rect 15476 27940 15528 27946
rect 15476 27882 15528 27888
rect 15099 27772 15407 27781
rect 15099 27770 15105 27772
rect 15161 27770 15185 27772
rect 15241 27770 15265 27772
rect 15321 27770 15345 27772
rect 15401 27770 15407 27772
rect 15161 27718 15163 27770
rect 15343 27718 15345 27770
rect 15099 27716 15105 27718
rect 15161 27716 15185 27718
rect 15241 27716 15265 27718
rect 15321 27716 15345 27718
rect 15401 27716 15407 27718
rect 15099 27707 15407 27716
rect 15488 27674 15516 27882
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 15580 27674 15608 27814
rect 15476 27668 15528 27674
rect 15476 27610 15528 27616
rect 15568 27668 15620 27674
rect 15568 27610 15620 27616
rect 14924 27396 14976 27402
rect 14924 27338 14976 27344
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 14832 27124 14884 27130
rect 14660 27084 14832 27112
rect 14280 27056 14332 27062
rect 14280 26998 14332 27004
rect 14200 26846 14320 26874
rect 14660 26858 14688 27084
rect 14832 27066 14884 27072
rect 15488 26926 15516 27270
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 14188 26784 14240 26790
rect 14188 26726 14240 26732
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 14200 26450 14228 26726
rect 14188 26444 14240 26450
rect 14188 26386 14240 26392
rect 13924 26166 14044 26194
rect 13636 25832 13688 25838
rect 13636 25774 13688 25780
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 13268 25492 13320 25498
rect 13268 25434 13320 25440
rect 13452 25492 13504 25498
rect 13452 25434 13504 25440
rect 13464 24342 13492 25434
rect 13648 25226 13676 25774
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 13636 25220 13688 25226
rect 13636 25162 13688 25168
rect 13648 24818 13676 25162
rect 13740 24954 13768 25298
rect 13728 24948 13780 24954
rect 13728 24890 13780 24896
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13452 24336 13504 24342
rect 13452 24278 13504 24284
rect 13452 24200 13504 24206
rect 13452 24142 13504 24148
rect 13464 23866 13492 24142
rect 13740 23866 13768 24890
rect 13452 23860 13504 23866
rect 13452 23802 13504 23808
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13740 23474 13768 23802
rect 13556 23446 13768 23474
rect 13820 23520 13872 23526
rect 13820 23462 13872 23468
rect 13556 22098 13584 23446
rect 13832 23118 13860 23462
rect 13728 23112 13780 23118
rect 13728 23054 13780 23060
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13740 22778 13768 23054
rect 13728 22772 13780 22778
rect 13728 22714 13780 22720
rect 13924 22420 13952 26166
rect 14188 25696 14240 25702
rect 14188 25638 14240 25644
rect 14200 25430 14228 25638
rect 14188 25424 14240 25430
rect 14188 25366 14240 25372
rect 14292 24426 14320 26846
rect 14648 26852 14700 26858
rect 14648 26794 14700 26800
rect 14832 26852 14884 26858
rect 14832 26794 14884 26800
rect 15660 26852 15712 26858
rect 15660 26794 15712 26800
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14752 26450 14780 26726
rect 14740 26444 14792 26450
rect 14740 26386 14792 26392
rect 14844 26246 14872 26794
rect 15099 26684 15407 26693
rect 15099 26682 15105 26684
rect 15161 26682 15185 26684
rect 15241 26682 15265 26684
rect 15321 26682 15345 26684
rect 15401 26682 15407 26684
rect 15161 26630 15163 26682
rect 15343 26630 15345 26682
rect 15099 26628 15105 26630
rect 15161 26628 15185 26630
rect 15241 26628 15265 26630
rect 15321 26628 15345 26630
rect 15401 26628 15407 26630
rect 15099 26619 15407 26628
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 14832 26240 14884 26246
rect 14832 26182 14884 26188
rect 14439 26140 14747 26149
rect 14439 26138 14445 26140
rect 14501 26138 14525 26140
rect 14581 26138 14605 26140
rect 14661 26138 14685 26140
rect 14741 26138 14747 26140
rect 14501 26086 14503 26138
rect 14683 26086 14685 26138
rect 14439 26084 14445 26086
rect 14501 26084 14525 26086
rect 14581 26084 14605 26086
rect 14661 26084 14685 26086
rect 14741 26084 14747 26086
rect 14439 26075 14747 26084
rect 14844 25906 14872 26182
rect 14832 25900 14884 25906
rect 14832 25842 14884 25848
rect 15476 25764 15528 25770
rect 15476 25706 15528 25712
rect 14464 25696 14516 25702
rect 14464 25638 14516 25644
rect 14476 25294 14504 25638
rect 15099 25596 15407 25605
rect 15099 25594 15105 25596
rect 15161 25594 15185 25596
rect 15241 25594 15265 25596
rect 15321 25594 15345 25596
rect 15401 25594 15407 25596
rect 15161 25542 15163 25594
rect 15343 25542 15345 25594
rect 15099 25540 15105 25542
rect 15161 25540 15185 25542
rect 15241 25540 15265 25542
rect 15321 25540 15345 25542
rect 15401 25540 15407 25542
rect 15099 25531 15407 25540
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14439 25052 14747 25061
rect 14439 25050 14445 25052
rect 14501 25050 14525 25052
rect 14581 25050 14605 25052
rect 14661 25050 14685 25052
rect 14741 25050 14747 25052
rect 14501 24998 14503 25050
rect 14683 24998 14685 25050
rect 14439 24996 14445 24998
rect 14501 24996 14525 24998
rect 14581 24996 14605 24998
rect 14661 24996 14685 24998
rect 14741 24996 14747 24998
rect 14439 24987 14747 24996
rect 14292 24398 14412 24426
rect 14004 24336 14056 24342
rect 14004 24278 14056 24284
rect 14384 24290 14412 24398
rect 14016 23866 14044 24278
rect 14384 24274 14504 24290
rect 14384 24268 14516 24274
rect 14384 24262 14464 24268
rect 14464 24210 14516 24216
rect 14439 23964 14747 23973
rect 14439 23962 14445 23964
rect 14501 23962 14525 23964
rect 14581 23962 14605 23964
rect 14661 23962 14685 23964
rect 14741 23962 14747 23964
rect 14501 23910 14503 23962
rect 14683 23910 14685 23962
rect 14439 23908 14445 23910
rect 14501 23908 14525 23910
rect 14581 23908 14605 23910
rect 14661 23908 14685 23910
rect 14741 23908 14747 23910
rect 14439 23899 14747 23908
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 14188 23520 14240 23526
rect 14188 23462 14240 23468
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14108 22574 14136 23462
rect 14200 23254 14228 23462
rect 14292 23322 14320 23462
rect 14280 23316 14332 23322
rect 14280 23258 14332 23264
rect 14188 23248 14240 23254
rect 14188 23190 14240 23196
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14096 22568 14148 22574
rect 14096 22510 14148 22516
rect 13924 22392 14136 22420
rect 13544 22092 13596 22098
rect 13544 22034 13596 22040
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 13268 19780 13320 19786
rect 13268 19722 13320 19728
rect 13280 19514 13308 19722
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13372 17218 13400 20742
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13464 19378 13492 20198
rect 13556 19922 13584 22034
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 13636 20936 13688 20942
rect 13636 20878 13688 20884
rect 13648 20058 13676 20878
rect 13832 20602 13860 21966
rect 14016 21554 14044 21966
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13912 21480 13964 21486
rect 13912 21422 13964 21428
rect 13820 20596 13872 20602
rect 13820 20538 13872 20544
rect 13818 20088 13874 20097
rect 13636 20052 13688 20058
rect 13818 20023 13874 20032
rect 13636 19994 13688 20000
rect 13832 19990 13860 20023
rect 13820 19984 13872 19990
rect 13820 19926 13872 19932
rect 13544 19916 13596 19922
rect 13544 19858 13596 19864
rect 13832 19514 13860 19926
rect 13924 19854 13952 21422
rect 14004 19984 14056 19990
rect 14004 19926 14056 19932
rect 13912 19848 13964 19854
rect 13912 19790 13964 19796
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13452 19372 13504 19378
rect 13924 19334 13952 19790
rect 14016 19378 14044 19926
rect 13452 19314 13504 19320
rect 13740 19306 13952 19334
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 13740 18034 13768 19306
rect 13912 18828 13964 18834
rect 13912 18770 13964 18776
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13832 18426 13860 18566
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13820 18148 13872 18154
rect 13820 18090 13872 18096
rect 13832 18034 13860 18090
rect 13740 18006 13860 18034
rect 13452 17808 13504 17814
rect 13452 17750 13504 17756
rect 13464 17338 13492 17750
rect 13634 17640 13690 17649
rect 13634 17575 13690 17584
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13372 17190 13492 17218
rect 13188 17156 13308 17184
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 13096 16114 13124 16594
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13188 16250 13216 16458
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12992 15904 13044 15910
rect 12992 15846 13044 15852
rect 12808 15496 12860 15502
rect 12808 15438 12860 15444
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 14006 12848 14214
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12728 13790 12848 13818
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12164 11620 12216 11626
rect 12164 11562 12216 11568
rect 12176 11121 12204 11562
rect 12544 11218 12572 11834
rect 12636 11286 12664 12378
rect 12728 12102 12756 12922
rect 12716 12096 12768 12102
rect 12716 12038 12768 12044
rect 12728 11898 12756 12038
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12162 11112 12218 11121
rect 12162 11047 12218 11056
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11704 10532 11756 10538
rect 11704 10474 11756 10480
rect 11716 9722 11744 10474
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11716 8090 11744 9658
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11808 7954 11836 8502
rect 12084 8430 12112 9522
rect 12176 8566 12204 11047
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 10266 12572 10406
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12532 10056 12584 10062
rect 12532 9998 12584 10004
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11992 7954 12020 8026
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11796 7948 11848 7954
rect 11796 7890 11848 7896
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11980 7948 12032 7954
rect 11980 7890 12032 7896
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10416 7472 10468 7478
rect 10416 7414 10468 7420
rect 10796 7342 10824 7890
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 10784 7336 10836 7342
rect 10784 7278 10836 7284
rect 10232 7200 10284 7206
rect 10232 7142 10284 7148
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10244 6662 10272 7142
rect 10520 6866 10548 7142
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 10060 5098 10088 5510
rect 10152 5234 10180 6598
rect 10416 6316 10468 6322
rect 10416 6258 10468 6264
rect 10428 5710 10456 6258
rect 10796 5778 10824 7278
rect 11428 7200 11480 7206
rect 11428 7142 11480 7148
rect 11440 6866 11468 7142
rect 11428 6860 11480 6866
rect 11428 6802 11480 6808
rect 11520 6316 11572 6322
rect 11520 6258 11572 6264
rect 10876 6180 10928 6186
rect 10876 6122 10928 6128
rect 10888 5914 10916 6122
rect 10876 5908 10928 5914
rect 10876 5850 10928 5856
rect 10784 5772 10836 5778
rect 10784 5714 10836 5720
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 10048 5092 10100 5098
rect 10048 5034 10100 5040
rect 9692 4826 9720 5034
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 10152 4690 10180 5170
rect 10796 4690 10824 5714
rect 11532 5370 11560 6258
rect 11624 5778 11652 7686
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11716 5914 11744 6598
rect 11808 6118 11836 7890
rect 11900 7818 11928 7890
rect 11888 7812 11940 7818
rect 11888 7754 11940 7760
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11808 5846 11836 6054
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11520 5364 11572 5370
rect 11520 5306 11572 5312
rect 11808 4826 11836 5782
rect 11900 5710 11928 6598
rect 11992 5778 12020 7142
rect 12084 5778 12112 8366
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12176 7546 12204 7686
rect 12164 7540 12216 7546
rect 12164 7482 12216 7488
rect 12268 7410 12296 8910
rect 12544 8362 12572 9998
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12544 8090 12572 8298
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12268 6322 12296 7346
rect 12452 7002 12480 8026
rect 12820 7528 12848 13790
rect 12912 13530 12940 13942
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12912 13190 12940 13466
rect 13004 13462 13032 15846
rect 13096 15570 13124 16050
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13188 15638 13216 15914
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 13084 15564 13136 15570
rect 13084 15506 13136 15512
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 14890 13216 15302
rect 13280 15026 13308 17156
rect 13464 16590 13492 17190
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13452 15428 13504 15434
rect 13452 15370 13504 15376
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13176 14884 13228 14890
rect 13176 14826 13228 14832
rect 13280 14482 13308 14962
rect 13268 14476 13320 14482
rect 13268 14418 13320 14424
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13084 13796 13136 13802
rect 13084 13738 13136 13744
rect 13096 13462 13124 13738
rect 12992 13456 13044 13462
rect 12992 13398 13044 13404
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 13004 13274 13032 13398
rect 13188 13394 13216 13874
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 13004 13246 13124 13274
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12986 13032 13126
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12900 12708 12952 12714
rect 12900 12650 12952 12656
rect 12912 12442 12940 12650
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12900 12096 12952 12102
rect 12900 12038 12952 12044
rect 12912 11694 12940 12038
rect 13096 11898 13124 13246
rect 13176 12640 13228 12646
rect 13176 12582 13228 12588
rect 13188 12442 13216 12582
rect 13176 12436 13228 12442
rect 13176 12378 13228 12384
rect 13280 12306 13308 13806
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13372 13326 13400 13670
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13372 11898 13400 13262
rect 13464 12442 13492 15370
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13556 12356 13584 16526
rect 13648 15706 13676 17575
rect 13740 17270 13768 18006
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13820 17060 13872 17066
rect 13820 17002 13872 17008
rect 13832 16114 13860 17002
rect 13924 16998 13952 18770
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 14016 18426 14044 18634
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 13912 16992 13964 16998
rect 13912 16934 13964 16940
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13924 16046 13952 16934
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 14016 16250 14044 16662
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14108 16130 14136 22392
rect 14200 21554 14228 23054
rect 14439 22876 14747 22885
rect 14439 22874 14445 22876
rect 14501 22874 14525 22876
rect 14581 22874 14605 22876
rect 14661 22874 14685 22876
rect 14741 22874 14747 22876
rect 14501 22822 14503 22874
rect 14683 22822 14685 22874
rect 14439 22820 14445 22822
rect 14501 22820 14525 22822
rect 14581 22820 14605 22822
rect 14661 22820 14685 22822
rect 14741 22820 14747 22822
rect 14439 22811 14747 22820
rect 14844 22778 14872 23598
rect 14936 23186 14964 25434
rect 15099 24508 15407 24517
rect 15099 24506 15105 24508
rect 15161 24506 15185 24508
rect 15241 24506 15265 24508
rect 15321 24506 15345 24508
rect 15401 24506 15407 24508
rect 15161 24454 15163 24506
rect 15343 24454 15345 24506
rect 15099 24452 15105 24454
rect 15161 24452 15185 24454
rect 15241 24452 15265 24454
rect 15321 24452 15345 24454
rect 15401 24452 15407 24454
rect 15099 24443 15407 24452
rect 15099 23420 15407 23429
rect 15099 23418 15105 23420
rect 15161 23418 15185 23420
rect 15241 23418 15265 23420
rect 15321 23418 15345 23420
rect 15401 23418 15407 23420
rect 15161 23366 15163 23418
rect 15343 23366 15345 23418
rect 15099 23364 15105 23366
rect 15161 23364 15185 23366
rect 15241 23364 15265 23366
rect 15321 23364 15345 23366
rect 15401 23364 15407 23366
rect 15099 23355 15407 23364
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 14924 23180 14976 23186
rect 14924 23122 14976 23128
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14844 22166 14872 22374
rect 14832 22160 14884 22166
rect 14832 22102 14884 22108
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14439 21788 14747 21797
rect 14439 21786 14445 21788
rect 14501 21786 14525 21788
rect 14581 21786 14605 21788
rect 14661 21786 14685 21788
rect 14741 21786 14747 21788
rect 14501 21734 14503 21786
rect 14683 21734 14685 21786
rect 14439 21732 14445 21734
rect 14501 21732 14525 21734
rect 14581 21732 14605 21734
rect 14661 21732 14685 21734
rect 14741 21732 14747 21734
rect 14439 21723 14747 21732
rect 14372 21684 14424 21690
rect 14372 21626 14424 21632
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14200 19990 14228 21082
rect 14384 21078 14412 21626
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14660 21078 14688 21490
rect 14372 21072 14424 21078
rect 14372 21014 14424 21020
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 14280 20800 14332 20806
rect 14280 20742 14332 20748
rect 14292 20262 14320 20742
rect 14439 20700 14747 20709
rect 14439 20698 14445 20700
rect 14501 20698 14525 20700
rect 14581 20698 14605 20700
rect 14661 20698 14685 20700
rect 14741 20698 14747 20700
rect 14501 20646 14503 20698
rect 14683 20646 14685 20698
rect 14439 20644 14445 20646
rect 14501 20644 14525 20646
rect 14581 20644 14605 20646
rect 14661 20644 14685 20646
rect 14741 20644 14747 20646
rect 14439 20635 14747 20644
rect 14844 20466 14872 21966
rect 14936 21554 14964 23122
rect 15304 23118 15332 23258
rect 15200 23112 15252 23118
rect 15200 23054 15252 23060
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15212 22778 15240 23054
rect 15200 22772 15252 22778
rect 15200 22714 15252 22720
rect 15016 22568 15068 22574
rect 15016 22510 15068 22516
rect 15028 21690 15056 22510
rect 15099 22332 15407 22341
rect 15099 22330 15105 22332
rect 15161 22330 15185 22332
rect 15241 22330 15265 22332
rect 15321 22330 15345 22332
rect 15401 22330 15407 22332
rect 15161 22278 15163 22330
rect 15343 22278 15345 22330
rect 15099 22276 15105 22278
rect 15161 22276 15185 22278
rect 15241 22276 15265 22278
rect 15321 22276 15345 22278
rect 15401 22276 15407 22278
rect 15099 22267 15407 22276
rect 15016 21684 15068 21690
rect 15016 21626 15068 21632
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14188 19984 14240 19990
rect 14186 19952 14188 19961
rect 14240 19952 14242 19961
rect 14186 19887 14242 19896
rect 14439 19612 14747 19621
rect 14439 19610 14445 19612
rect 14501 19610 14525 19612
rect 14581 19610 14605 19612
rect 14661 19610 14685 19612
rect 14741 19610 14747 19612
rect 14501 19558 14503 19610
rect 14683 19558 14685 19610
rect 14439 19556 14445 19558
rect 14501 19556 14525 19558
rect 14581 19556 14605 19558
rect 14661 19556 14685 19558
rect 14741 19556 14747 19558
rect 14439 19547 14747 19556
rect 14370 19272 14426 19281
rect 14292 19230 14370 19258
rect 14292 18193 14320 19230
rect 14370 19207 14426 19216
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14568 18766 14596 19110
rect 14844 18970 14872 20402
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14439 18524 14747 18533
rect 14439 18522 14445 18524
rect 14501 18522 14525 18524
rect 14581 18522 14605 18524
rect 14661 18522 14685 18524
rect 14741 18522 14747 18524
rect 14501 18470 14503 18522
rect 14683 18470 14685 18522
rect 14439 18468 14445 18470
rect 14501 18468 14525 18470
rect 14581 18468 14605 18470
rect 14661 18468 14685 18470
rect 14741 18468 14747 18470
rect 14439 18459 14747 18468
rect 14936 18426 14964 19246
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 14922 18320 14978 18329
rect 14922 18255 14978 18264
rect 14278 18184 14334 18193
rect 14278 18119 14334 18128
rect 14188 17196 14240 17202
rect 14292 17184 14320 18119
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 14439 17436 14747 17445
rect 14439 17434 14445 17436
rect 14501 17434 14525 17436
rect 14581 17434 14605 17436
rect 14661 17434 14685 17436
rect 14741 17434 14747 17436
rect 14501 17382 14503 17434
rect 14683 17382 14685 17434
rect 14439 17380 14445 17382
rect 14501 17380 14525 17382
rect 14581 17380 14605 17382
rect 14661 17380 14685 17382
rect 14741 17380 14747 17382
rect 14439 17371 14747 17380
rect 14372 17196 14424 17202
rect 14292 17156 14372 17184
rect 14188 17138 14240 17144
rect 14372 17138 14424 17144
rect 14200 16998 14228 17138
rect 14844 17134 14872 17614
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14188 16992 14240 16998
rect 14188 16934 14240 16940
rect 14936 16538 14964 18255
rect 15028 17338 15056 21286
rect 15099 21244 15407 21253
rect 15099 21242 15105 21244
rect 15161 21242 15185 21244
rect 15241 21242 15265 21244
rect 15321 21242 15345 21244
rect 15401 21242 15407 21244
rect 15161 21190 15163 21242
rect 15343 21190 15345 21242
rect 15099 21188 15105 21190
rect 15161 21188 15185 21190
rect 15241 21188 15265 21190
rect 15321 21188 15345 21190
rect 15401 21188 15407 21190
rect 15099 21179 15407 21188
rect 15488 21146 15516 25706
rect 15580 25226 15608 26386
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15672 24818 15700 26794
rect 15764 26586 15792 28154
rect 15856 27470 15884 28562
rect 16028 27940 16080 27946
rect 16028 27882 16080 27888
rect 16040 27674 16068 27882
rect 16028 27668 16080 27674
rect 16028 27610 16080 27616
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15856 27130 15884 27406
rect 15844 27124 15896 27130
rect 15844 27066 15896 27072
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15948 27033 15976 27066
rect 15934 27024 15990 27033
rect 15934 26959 15990 26968
rect 15752 26580 15804 26586
rect 15752 26522 15804 26528
rect 15844 26240 15896 26246
rect 15844 26182 15896 26188
rect 15856 25770 15884 26182
rect 15844 25764 15896 25770
rect 15844 25706 15896 25712
rect 15844 25220 15896 25226
rect 15844 25162 15896 25168
rect 15856 24954 15884 25162
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15580 23769 15608 24550
rect 15672 24206 15700 24754
rect 15752 24744 15804 24750
rect 15752 24686 15804 24692
rect 15660 24200 15712 24206
rect 15660 24142 15712 24148
rect 15764 23866 15792 24686
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15566 23760 15622 23769
rect 15566 23695 15622 23704
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 15672 21350 15700 23462
rect 15764 23118 15792 23462
rect 15752 23112 15804 23118
rect 15752 23054 15804 23060
rect 15844 22092 15896 22098
rect 15844 22034 15896 22040
rect 15856 21690 15884 22034
rect 15844 21684 15896 21690
rect 15844 21626 15896 21632
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15476 21140 15528 21146
rect 15476 21082 15528 21088
rect 15936 20800 15988 20806
rect 15936 20742 15988 20748
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15212 20330 15516 20346
rect 15200 20324 15516 20330
rect 15252 20318 15516 20324
rect 15200 20266 15252 20272
rect 15099 20156 15407 20165
rect 15099 20154 15105 20156
rect 15161 20154 15185 20156
rect 15241 20154 15265 20156
rect 15321 20154 15345 20156
rect 15401 20154 15407 20156
rect 15161 20102 15163 20154
rect 15343 20102 15345 20154
rect 15099 20100 15105 20102
rect 15161 20100 15185 20102
rect 15241 20100 15265 20102
rect 15321 20100 15345 20102
rect 15401 20100 15407 20102
rect 15099 20091 15407 20100
rect 15488 19514 15516 20318
rect 15580 20058 15608 20402
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15099 19068 15407 19077
rect 15099 19066 15105 19068
rect 15161 19066 15185 19068
rect 15241 19066 15265 19068
rect 15321 19066 15345 19068
rect 15401 19066 15407 19068
rect 15161 19014 15163 19066
rect 15343 19014 15345 19066
rect 15099 19012 15105 19014
rect 15161 19012 15185 19014
rect 15241 19012 15265 19014
rect 15321 19012 15345 19014
rect 15401 19012 15407 19014
rect 15099 19003 15407 19012
rect 15580 18902 15608 19110
rect 15568 18896 15620 18902
rect 15568 18838 15620 18844
rect 15099 17980 15407 17989
rect 15099 17978 15105 17980
rect 15161 17978 15185 17980
rect 15241 17978 15265 17980
rect 15321 17978 15345 17980
rect 15401 17978 15407 17980
rect 15161 17926 15163 17978
rect 15343 17926 15345 17978
rect 15099 17924 15105 17926
rect 15161 17924 15185 17926
rect 15241 17924 15265 17926
rect 15321 17924 15345 17926
rect 15401 17924 15407 17926
rect 15099 17915 15407 17924
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15016 17332 15068 17338
rect 15016 17274 15068 17280
rect 15488 17270 15516 17478
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15099 16892 15407 16901
rect 15099 16890 15105 16892
rect 15161 16890 15185 16892
rect 15241 16890 15265 16892
rect 15321 16890 15345 16892
rect 15401 16890 15407 16892
rect 15161 16838 15163 16890
rect 15343 16838 15345 16890
rect 15099 16836 15105 16838
rect 15161 16836 15185 16838
rect 15241 16836 15265 16838
rect 15321 16836 15345 16838
rect 15401 16836 15407 16838
rect 15099 16827 15407 16836
rect 15580 16726 15608 17070
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15672 16590 15700 17002
rect 14844 16510 14964 16538
rect 15660 16584 15712 16590
rect 15660 16526 15712 16532
rect 14439 16348 14747 16357
rect 14439 16346 14445 16348
rect 14501 16346 14525 16348
rect 14581 16346 14605 16348
rect 14661 16346 14685 16348
rect 14741 16346 14747 16348
rect 14501 16294 14503 16346
rect 14683 16294 14685 16346
rect 14439 16292 14445 16294
rect 14501 16292 14525 16294
rect 14581 16292 14605 16294
rect 14661 16292 14685 16294
rect 14741 16292 14747 16294
rect 14439 16283 14747 16292
rect 14016 16102 14136 16130
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 14884 13688 14890
rect 13636 14826 13688 14832
rect 13648 14618 13676 14826
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13740 14006 13768 15574
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13924 15026 13952 15438
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13832 14074 13860 14758
rect 13924 14414 13952 14758
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13728 14000 13780 14006
rect 13728 13942 13780 13948
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13832 12986 13860 13398
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13832 12442 13860 12922
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13556 12328 13676 12356
rect 13648 12322 13676 12328
rect 13648 12294 13768 12322
rect 13740 12238 13768 12294
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11150 12940 11494
rect 13096 11218 13124 11834
rect 13372 11354 13400 11834
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 13004 10538 13032 10950
rect 13188 10810 13216 10950
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13464 10606 13492 11698
rect 13740 11354 13768 12174
rect 13924 11801 13952 14350
rect 13910 11792 13966 11801
rect 13910 11727 13966 11736
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13740 11150 13768 11290
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 12992 10532 13044 10538
rect 12992 10474 13044 10480
rect 13084 10532 13136 10538
rect 13084 10474 13136 10480
rect 13096 9382 13124 10474
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13268 10192 13320 10198
rect 13268 10134 13320 10140
rect 13280 9722 13308 10134
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13096 8634 13124 9318
rect 13280 9178 13308 9318
rect 13268 9172 13320 9178
rect 13268 9114 13320 9120
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13556 8430 13584 10202
rect 13924 9518 13952 11727
rect 14016 11014 14044 16102
rect 14740 15632 14792 15638
rect 14844 15620 14872 16510
rect 14924 16448 14976 16454
rect 14924 16390 14976 16396
rect 14792 15592 14872 15620
rect 14740 15574 14792 15580
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14188 14952 14240 14958
rect 14188 14894 14240 14900
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14108 13938 14136 14214
rect 14200 13954 14228 14894
rect 14292 14074 14320 15302
rect 14439 15260 14747 15269
rect 14439 15258 14445 15260
rect 14501 15258 14525 15260
rect 14581 15258 14605 15260
rect 14661 15258 14685 15260
rect 14741 15258 14747 15260
rect 14501 15206 14503 15258
rect 14683 15206 14685 15258
rect 14439 15204 14445 15206
rect 14501 15204 14525 15206
rect 14581 15204 14605 15206
rect 14661 15204 14685 15206
rect 14741 15204 14747 15206
rect 14439 15195 14747 15204
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14464 14816 14516 14822
rect 14464 14758 14516 14764
rect 14476 14618 14504 14758
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14752 14414 14780 14894
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14439 14172 14747 14181
rect 14439 14170 14445 14172
rect 14501 14170 14525 14172
rect 14581 14170 14605 14172
rect 14661 14170 14685 14172
rect 14741 14170 14747 14172
rect 14501 14118 14503 14170
rect 14683 14118 14685 14170
rect 14439 14116 14445 14118
rect 14501 14116 14525 14118
rect 14581 14116 14605 14118
rect 14661 14116 14685 14118
rect 14741 14116 14747 14118
rect 14439 14107 14747 14116
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14844 13954 14872 15098
rect 14936 14482 14964 16390
rect 15672 16182 15700 16526
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15099 15804 15407 15813
rect 15099 15802 15105 15804
rect 15161 15802 15185 15804
rect 15241 15802 15265 15804
rect 15321 15802 15345 15804
rect 15401 15802 15407 15804
rect 15161 15750 15163 15802
rect 15343 15750 15345 15802
rect 15099 15748 15105 15750
rect 15161 15748 15185 15750
rect 15241 15748 15265 15750
rect 15321 15748 15345 15750
rect 15401 15748 15407 15750
rect 15099 15739 15407 15748
rect 15488 15638 15516 15846
rect 15764 15706 15792 19314
rect 15948 16794 15976 20742
rect 16028 20324 16080 20330
rect 16028 20266 16080 20272
rect 16040 20058 16068 20266
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16132 18834 16160 31726
rect 16592 31346 16620 31758
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16488 31272 16540 31278
rect 16488 31214 16540 31220
rect 16304 31136 16356 31142
rect 16304 31078 16356 31084
rect 16316 30190 16344 31078
rect 16500 30938 16528 31214
rect 16580 31204 16632 31210
rect 16580 31146 16632 31152
rect 16488 30932 16540 30938
rect 16488 30874 16540 30880
rect 16592 30802 16620 31146
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16304 30184 16356 30190
rect 16304 30126 16356 30132
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16224 29170 16252 29990
rect 16486 29200 16542 29209
rect 16212 29164 16264 29170
rect 16486 29135 16488 29144
rect 16212 29106 16264 29112
rect 16540 29135 16542 29144
rect 16488 29106 16540 29112
rect 16592 28762 16620 30738
rect 16856 30184 16908 30190
rect 16856 30126 16908 30132
rect 16868 29850 16896 30126
rect 16856 29844 16908 29850
rect 16856 29786 16908 29792
rect 16580 28756 16632 28762
rect 16580 28698 16632 28704
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16408 28218 16436 28562
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 16592 27674 16620 28698
rect 16960 28234 16988 33798
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 18340 32434 18368 32710
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 17776 31816 17828 31822
rect 17776 31758 17828 31764
rect 17224 31680 17276 31686
rect 17224 31622 17276 31628
rect 17236 31346 17264 31622
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17788 30938 17816 31758
rect 17868 31680 17920 31686
rect 17868 31622 17920 31628
rect 17776 30932 17828 30938
rect 17776 30874 17828 30880
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17132 29028 17184 29034
rect 17132 28970 17184 28976
rect 17144 28762 17172 28970
rect 17132 28756 17184 28762
rect 17132 28698 17184 28704
rect 16868 28206 16988 28234
rect 16764 27940 16816 27946
rect 16764 27882 16816 27888
rect 16776 27674 16804 27882
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 16764 27668 16816 27674
rect 16764 27610 16816 27616
rect 16304 26852 16356 26858
rect 16304 26794 16356 26800
rect 16316 26586 16344 26794
rect 16304 26580 16356 26586
rect 16304 26522 16356 26528
rect 16580 26444 16632 26450
rect 16580 26386 16632 26392
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16408 25430 16436 25774
rect 16396 25424 16448 25430
rect 16396 25366 16448 25372
rect 16592 25226 16620 26386
rect 16672 25764 16724 25770
rect 16672 25706 16724 25712
rect 16684 25294 16712 25706
rect 16672 25288 16724 25294
rect 16672 25230 16724 25236
rect 16580 25220 16632 25226
rect 16580 25162 16632 25168
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16408 23798 16436 24754
rect 16592 24698 16620 25162
rect 16670 24848 16726 24857
rect 16868 24818 16896 28206
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 16670 24783 16672 24792
rect 16724 24783 16726 24792
rect 16856 24812 16908 24818
rect 16672 24754 16724 24760
rect 16856 24754 16908 24760
rect 16948 24744 17000 24750
rect 16592 24670 16712 24698
rect 16948 24686 17000 24692
rect 16396 23792 16448 23798
rect 16396 23734 16448 23740
rect 16488 23248 16540 23254
rect 16486 23216 16488 23225
rect 16540 23216 16542 23225
rect 16486 23151 16542 23160
rect 16580 23180 16632 23186
rect 16580 23122 16632 23128
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 16316 22778 16344 22918
rect 16592 22778 16620 23122
rect 16304 22772 16356 22778
rect 16304 22714 16356 22720
rect 16580 22772 16632 22778
rect 16580 22714 16632 22720
rect 16684 22574 16712 24670
rect 16960 24206 16988 24686
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 16856 23656 16908 23662
rect 16856 23598 16908 23604
rect 16868 22982 16896 23598
rect 16856 22976 16908 22982
rect 16856 22918 16908 22924
rect 16672 22568 16724 22574
rect 16672 22510 16724 22516
rect 16684 22094 16712 22510
rect 16684 22066 16804 22094
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16684 21554 16712 21830
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 16776 21418 16804 22066
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16672 21344 16724 21350
rect 16672 21286 16724 21292
rect 16684 20874 16712 21286
rect 16776 20874 16804 21354
rect 16868 21010 16896 22918
rect 16856 21004 16908 21010
rect 16856 20946 16908 20952
rect 16672 20868 16724 20874
rect 16672 20810 16724 20816
rect 16764 20868 16816 20874
rect 16764 20810 16816 20816
rect 16960 20448 16988 24142
rect 16592 20420 16988 20448
rect 16396 19984 16448 19990
rect 16396 19926 16448 19932
rect 16408 19514 16436 19926
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16396 19508 16448 19514
rect 16396 19450 16448 19456
rect 16408 19378 16436 19450
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16500 19310 16528 19790
rect 16488 19304 16540 19310
rect 16488 19246 16540 19252
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16026 17912 16082 17921
rect 16026 17847 16082 17856
rect 16040 17814 16068 17847
rect 16028 17808 16080 17814
rect 16028 17750 16080 17756
rect 16120 17808 16172 17814
rect 16120 17750 16172 17756
rect 16028 17060 16080 17066
rect 16028 17002 16080 17008
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15476 15632 15528 15638
rect 15476 15574 15528 15580
rect 15856 15502 15884 16730
rect 16040 16250 16068 17002
rect 16132 16794 16160 17750
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15856 14958 15884 15438
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15476 14816 15528 14822
rect 15476 14758 15528 14764
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15099 14716 15407 14725
rect 15099 14714 15105 14716
rect 15161 14714 15185 14716
rect 15241 14714 15265 14716
rect 15321 14714 15345 14716
rect 15401 14714 15407 14716
rect 15161 14662 15163 14714
rect 15343 14662 15345 14714
rect 15099 14660 15105 14662
rect 15161 14660 15185 14662
rect 15241 14660 15265 14662
rect 15321 14660 15345 14662
rect 15401 14660 15407 14662
rect 15099 14651 15407 14660
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 14924 14476 14976 14482
rect 14924 14418 14976 14424
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14096 13932 14148 13938
rect 14200 13926 14320 13954
rect 14096 13874 14148 13880
rect 14292 13870 14320 13926
rect 14660 13926 14872 13954
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 14464 13864 14516 13870
rect 14516 13812 14596 13818
rect 14464 13806 14596 13812
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14200 12714 14228 13262
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14200 11762 14228 12650
rect 14292 12442 14320 13806
rect 14476 13790 14596 13806
rect 14464 13728 14516 13734
rect 14464 13670 14516 13676
rect 14476 13530 14504 13670
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14568 13462 14596 13790
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14660 13258 14688 13926
rect 14738 13832 14794 13841
rect 14738 13767 14794 13776
rect 14752 13394 14780 13767
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14752 13274 14780 13330
rect 14648 13252 14700 13258
rect 14752 13246 14872 13274
rect 14648 13194 14700 13200
rect 14439 13084 14747 13093
rect 14439 13082 14445 13084
rect 14501 13082 14525 13084
rect 14581 13082 14605 13084
rect 14661 13082 14685 13084
rect 14741 13082 14747 13084
rect 14501 13030 14503 13082
rect 14683 13030 14685 13082
rect 14439 13028 14445 13030
rect 14501 13028 14525 13030
rect 14581 13028 14605 13030
rect 14661 13028 14685 13030
rect 14741 13028 14747 13030
rect 14439 13019 14747 13028
rect 14280 12436 14332 12442
rect 14844 12434 14872 13246
rect 14936 12646 14964 14214
rect 15212 13818 15240 14554
rect 15488 14113 15516 14758
rect 15474 14104 15530 14113
rect 15580 14074 15608 14758
rect 15856 14618 15884 14894
rect 16132 14822 16160 15506
rect 16224 14890 16252 15846
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 16132 14550 16160 14758
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 15936 14476 15988 14482
rect 15936 14418 15988 14424
rect 15660 14272 15712 14278
rect 15660 14214 15712 14220
rect 15474 14039 15530 14048
rect 15568 14068 15620 14074
rect 15488 13870 15516 14039
rect 15568 14010 15620 14016
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15028 13802 15240 13818
rect 15476 13864 15528 13870
rect 15580 13841 15608 13874
rect 15476 13806 15528 13812
rect 15566 13832 15622 13841
rect 15016 13796 15240 13802
rect 15068 13790 15240 13796
rect 15566 13767 15622 13776
rect 15016 13738 15068 13744
rect 15566 13696 15622 13705
rect 15099 13628 15407 13637
rect 15566 13631 15622 13640
rect 15099 13626 15105 13628
rect 15161 13626 15185 13628
rect 15241 13626 15265 13628
rect 15321 13626 15345 13628
rect 15401 13626 15407 13628
rect 15161 13574 15163 13626
rect 15343 13574 15345 13626
rect 15099 13572 15105 13574
rect 15161 13572 15185 13574
rect 15241 13572 15265 13574
rect 15321 13572 15345 13574
rect 15401 13572 15407 13574
rect 15099 13563 15407 13572
rect 15580 13530 15608 13631
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15580 13394 15608 13466
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15198 13288 15254 13297
rect 15016 13252 15068 13258
rect 15198 13223 15254 13232
rect 15016 13194 15068 13200
rect 15028 12918 15056 13194
rect 15016 12912 15068 12918
rect 15016 12854 15068 12860
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14280 12378 14332 12384
rect 14660 12406 14872 12434
rect 14660 12306 14688 12406
rect 14648 12300 14700 12306
rect 14648 12242 14700 12248
rect 14936 12186 14964 12582
rect 15028 12306 15056 12854
rect 15212 12850 15240 13223
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15488 12889 15516 13126
rect 15474 12880 15530 12889
rect 15200 12844 15252 12850
rect 15474 12815 15476 12824
rect 15200 12786 15252 12792
rect 15528 12815 15530 12824
rect 15476 12786 15528 12792
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15099 12540 15407 12549
rect 15099 12538 15105 12540
rect 15161 12538 15185 12540
rect 15241 12538 15265 12540
rect 15321 12538 15345 12540
rect 15401 12538 15407 12540
rect 15161 12486 15163 12538
rect 15343 12486 15345 12538
rect 15099 12484 15105 12486
rect 15161 12484 15185 12486
rect 15241 12484 15265 12486
rect 15321 12484 15345 12486
rect 15401 12484 15407 12486
rect 15099 12475 15407 12484
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15476 12232 15528 12238
rect 15474 12200 15476 12209
rect 15528 12200 15530 12209
rect 14832 12164 14884 12170
rect 14936 12158 15056 12186
rect 14832 12106 14884 12112
rect 14439 11996 14747 12005
rect 14439 11994 14445 11996
rect 14501 11994 14525 11996
rect 14581 11994 14605 11996
rect 14661 11994 14685 11996
rect 14741 11994 14747 11996
rect 14501 11942 14503 11994
rect 14683 11942 14685 11994
rect 14439 11940 14445 11942
rect 14501 11940 14525 11942
rect 14581 11940 14605 11942
rect 14661 11940 14685 11942
rect 14741 11940 14747 11942
rect 14439 11931 14747 11940
rect 14844 11898 14872 12106
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14188 11756 14240 11762
rect 14188 11698 14240 11704
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14004 11008 14056 11014
rect 14004 10950 14056 10956
rect 14200 10606 14228 11154
rect 14752 11121 14780 11154
rect 14738 11112 14794 11121
rect 14738 11047 14794 11056
rect 14439 10908 14747 10917
rect 14439 10906 14445 10908
rect 14501 10906 14525 10908
rect 14581 10906 14605 10908
rect 14661 10906 14685 10908
rect 14741 10906 14747 10908
rect 14501 10854 14503 10906
rect 14683 10854 14685 10906
rect 14439 10852 14445 10854
rect 14501 10852 14525 10854
rect 14581 10852 14605 10854
rect 14661 10852 14685 10854
rect 14741 10852 14747 10854
rect 14439 10843 14747 10852
rect 14936 10742 14964 12038
rect 15028 11762 15056 12158
rect 15580 12170 15608 12718
rect 15474 12135 15530 12144
rect 15568 12164 15620 12170
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15212 11762 15240 11834
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15099 11452 15407 11461
rect 15099 11450 15105 11452
rect 15161 11450 15185 11452
rect 15241 11450 15265 11452
rect 15321 11450 15345 11452
rect 15401 11450 15407 11452
rect 15161 11398 15163 11450
rect 15343 11398 15345 11450
rect 15099 11396 15105 11398
rect 15161 11396 15185 11398
rect 15241 11396 15265 11398
rect 15321 11396 15345 11398
rect 15401 11396 15407 11398
rect 15099 11387 15407 11396
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14188 10600 14240 10606
rect 14188 10542 14240 10548
rect 14200 9654 14228 10542
rect 14292 10130 14320 10610
rect 15099 10364 15407 10373
rect 15099 10362 15105 10364
rect 15161 10362 15185 10364
rect 15241 10362 15265 10364
rect 15321 10362 15345 10364
rect 15401 10362 15407 10364
rect 15161 10310 15163 10362
rect 15343 10310 15345 10362
rect 15099 10308 15105 10310
rect 15161 10308 15185 10310
rect 15241 10308 15265 10310
rect 15321 10308 15345 10310
rect 15401 10308 15407 10310
rect 15099 10299 15407 10308
rect 14832 10192 14884 10198
rect 14832 10134 14884 10140
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 13912 9512 13964 9518
rect 13912 9454 13964 9460
rect 13924 8956 13952 9454
rect 14200 9194 14228 9590
rect 13832 8928 13952 8956
rect 14108 9166 14228 9194
rect 14292 9194 14320 10066
rect 14439 9820 14747 9829
rect 14439 9818 14445 9820
rect 14501 9818 14525 9820
rect 14581 9818 14605 9820
rect 14661 9818 14685 9820
rect 14741 9818 14747 9820
rect 14501 9766 14503 9818
rect 14683 9766 14685 9818
rect 14439 9764 14445 9766
rect 14501 9764 14525 9766
rect 14581 9764 14605 9766
rect 14661 9764 14685 9766
rect 14741 9764 14747 9766
rect 14439 9755 14747 9764
rect 14844 9722 14872 10134
rect 15488 9738 15516 12135
rect 15568 12106 15620 12112
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15580 11354 15608 11834
rect 15672 11762 15700 14214
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15764 13530 15792 13806
rect 15844 13796 15896 13802
rect 15844 13738 15896 13744
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15856 12322 15884 13738
rect 15948 13190 15976 14418
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16132 14074 16160 14350
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 16040 12918 16068 13942
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15764 12294 15884 12322
rect 15764 12238 15792 12294
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15844 12232 15896 12238
rect 15844 12174 15896 12180
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15580 10198 15608 10406
rect 15568 10192 15620 10198
rect 15568 10134 15620 10140
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 15396 9710 15516 9738
rect 15396 9654 15424 9710
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15099 9276 15407 9285
rect 15099 9274 15105 9276
rect 15161 9274 15185 9276
rect 15241 9274 15265 9276
rect 15321 9274 15345 9276
rect 15401 9274 15407 9276
rect 15161 9222 15163 9274
rect 15343 9222 15345 9274
rect 15099 9220 15105 9222
rect 15161 9220 15185 9222
rect 15241 9220 15265 9222
rect 15321 9220 15345 9222
rect 15401 9220 15407 9222
rect 15099 9211 15407 9220
rect 14292 9166 14412 9194
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 7546 13676 7822
rect 12544 7500 12848 7528
rect 13636 7540 13688 7546
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12440 6792 12492 6798
rect 12440 6734 12492 6740
rect 12452 6458 12480 6734
rect 12440 6452 12492 6458
rect 12440 6394 12492 6400
rect 12256 6316 12308 6322
rect 12256 6258 12308 6264
rect 12544 6254 12572 7500
rect 13636 7482 13688 7488
rect 13544 7200 13596 7206
rect 13544 7142 13596 7148
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12912 6254 12940 6938
rect 13556 6322 13584 7142
rect 13740 6866 13768 8570
rect 13832 8498 13860 8928
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13924 8362 13952 8774
rect 14108 8498 14136 9166
rect 14384 9110 14412 9166
rect 14188 9104 14240 9110
rect 14188 9046 14240 9052
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14554 9072 14610 9081
rect 14200 8634 14228 9046
rect 14554 9007 14610 9016
rect 14924 9036 14976 9042
rect 14568 8974 14596 9007
rect 14924 8978 14976 8984
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14439 8732 14747 8741
rect 14439 8730 14445 8732
rect 14501 8730 14525 8732
rect 14581 8730 14605 8732
rect 14661 8730 14685 8732
rect 14741 8730 14747 8732
rect 14501 8678 14503 8730
rect 14683 8678 14685 8730
rect 14439 8676 14445 8678
rect 14501 8676 14525 8678
rect 14581 8676 14605 8678
rect 14661 8676 14685 8678
rect 14741 8676 14747 8678
rect 14439 8667 14747 8676
rect 14844 8634 14872 8774
rect 14188 8628 14240 8634
rect 14188 8570 14240 8576
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14936 8514 14964 8978
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14752 8486 14964 8514
rect 13912 8356 13964 8362
rect 13912 8298 13964 8304
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13832 6458 13860 7278
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12176 5914 12204 6122
rect 12164 5908 12216 5914
rect 12164 5850 12216 5856
rect 11980 5772 12032 5778
rect 11980 5714 12032 5720
rect 12072 5772 12124 5778
rect 12072 5714 12124 5720
rect 11888 5704 11940 5710
rect 12164 5704 12216 5710
rect 11888 5646 11940 5652
rect 12162 5672 12164 5681
rect 12348 5704 12400 5710
rect 12216 5672 12218 5681
rect 12348 5646 12400 5652
rect 12162 5607 12218 5616
rect 12256 5636 12308 5642
rect 12256 5578 12308 5584
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 11808 4690 11836 4762
rect 10140 4684 10192 4690
rect 10140 4626 10192 4632
rect 10784 4684 10836 4690
rect 10784 4626 10836 4632
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11900 4622 11928 5306
rect 12268 4826 12296 5578
rect 12360 5234 12388 5646
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 9496 4616 9548 4622
rect 9496 4558 9548 4564
rect 11888 4616 11940 4622
rect 11888 4558 11940 4564
rect 9508 4282 9536 4558
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 12544 4146 12572 6190
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12820 5914 12848 6122
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 13372 5846 13400 6054
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13268 5160 13320 5166
rect 13268 5102 13320 5108
rect 13280 5030 13308 5102
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 9680 3392 9732 3398
rect 9680 3334 9732 3340
rect 9692 3194 9720 3334
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 9128 2916 9180 2922
rect 9128 2858 9180 2864
rect 10980 800 11008 2926
rect 12268 800 12296 2994
rect 13280 2990 13308 4966
rect 13372 4622 13400 5782
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13740 5574 13768 5646
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13740 5234 13768 5510
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13648 4282 13676 4558
rect 13636 4276 13688 4282
rect 13636 4218 13688 4224
rect 13740 4146 13768 5170
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13636 3460 13688 3466
rect 13636 3402 13688 3408
rect 13648 3194 13676 3402
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13924 2990 13952 8298
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 4078 14044 7686
rect 14108 7546 14136 8434
rect 14188 8016 14240 8022
rect 14188 7958 14240 7964
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14200 7002 14228 7958
rect 14752 7954 14780 8486
rect 14924 8288 14976 8294
rect 14924 8230 14976 8236
rect 15384 8288 15436 8294
rect 15568 8288 15620 8294
rect 15436 8248 15516 8276
rect 15384 8230 15436 8236
rect 14936 8090 14964 8230
rect 15099 8188 15407 8197
rect 15099 8186 15105 8188
rect 15161 8186 15185 8188
rect 15241 8186 15265 8188
rect 15321 8186 15345 8188
rect 15401 8186 15407 8188
rect 15161 8134 15163 8186
rect 15343 8134 15345 8186
rect 15099 8132 15105 8134
rect 15161 8132 15185 8134
rect 15241 8132 15265 8134
rect 15321 8132 15345 8134
rect 15401 8132 15407 8134
rect 15099 8123 15407 8132
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 15292 8016 15344 8022
rect 15292 7958 15344 7964
rect 14740 7948 14792 7954
rect 14740 7890 14792 7896
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14292 7206 14320 7822
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 14439 7644 14747 7653
rect 14439 7642 14445 7644
rect 14501 7642 14525 7644
rect 14581 7642 14605 7644
rect 14661 7642 14685 7644
rect 14741 7642 14747 7644
rect 14501 7590 14503 7642
rect 14683 7590 14685 7642
rect 14439 7588 14445 7590
rect 14501 7588 14525 7590
rect 14581 7588 14605 7590
rect 14661 7588 14685 7590
rect 14741 7588 14747 7590
rect 14439 7579 14747 7588
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 14439 6556 14747 6565
rect 14439 6554 14445 6556
rect 14501 6554 14525 6556
rect 14581 6554 14605 6556
rect 14661 6554 14685 6556
rect 14741 6554 14747 6556
rect 14501 6502 14503 6554
rect 14683 6502 14685 6554
rect 14439 6500 14445 6502
rect 14501 6500 14525 6502
rect 14581 6500 14605 6502
rect 14661 6500 14685 6502
rect 14741 6500 14747 6502
rect 14439 6491 14747 6500
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14096 5772 14148 5778
rect 14096 5714 14148 5720
rect 14108 5370 14136 5714
rect 14200 5370 14228 6122
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14476 5778 14504 6054
rect 14464 5772 14516 5778
rect 14464 5714 14516 5720
rect 14439 5468 14747 5477
rect 14439 5466 14445 5468
rect 14501 5466 14525 5468
rect 14581 5466 14605 5468
rect 14661 5466 14685 5468
rect 14741 5466 14747 5468
rect 14501 5414 14503 5466
rect 14683 5414 14685 5466
rect 14439 5412 14445 5414
rect 14501 5412 14525 5414
rect 14581 5412 14605 5414
rect 14661 5412 14685 5414
rect 14741 5412 14747 5414
rect 14439 5403 14747 5412
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14188 5364 14240 5370
rect 14188 5306 14240 5312
rect 14844 5166 14872 7414
rect 15212 7274 15240 7686
rect 15304 7342 15332 7958
rect 15488 7546 15516 8248
rect 15568 8230 15620 8236
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15580 7410 15608 8230
rect 15568 7404 15620 7410
rect 15568 7346 15620 7352
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15099 7100 15407 7109
rect 15099 7098 15105 7100
rect 15161 7098 15185 7100
rect 15241 7098 15265 7100
rect 15321 7098 15345 7100
rect 15401 7098 15407 7100
rect 15161 7046 15163 7098
rect 15343 7046 15345 7098
rect 15099 7044 15105 7046
rect 15161 7044 15185 7046
rect 15241 7044 15265 7046
rect 15321 7044 15345 7046
rect 15401 7044 15407 7046
rect 15099 7035 15407 7044
rect 15488 6458 15516 7278
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15672 6254 15700 10950
rect 15764 10606 15792 12038
rect 15856 11830 15884 12174
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15856 11354 15884 11766
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15948 11286 15976 12650
rect 16040 12306 16068 12718
rect 16132 12374 16160 13874
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 16040 11762 16068 12242
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 15936 11280 15988 11286
rect 15934 11248 15936 11257
rect 15988 11248 15990 11257
rect 15934 11183 15990 11192
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10606 15976 10950
rect 16224 10674 16252 14826
rect 16316 14006 16344 18226
rect 16408 17202 16436 18702
rect 16592 17678 16620 20420
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16776 20058 16804 20198
rect 17052 20058 17080 27610
rect 17236 27606 17264 30534
rect 17592 29708 17644 29714
rect 17592 29650 17644 29656
rect 17604 29306 17632 29650
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17696 29186 17724 30738
rect 17880 30734 17908 31622
rect 18432 31482 18460 34002
rect 18708 33454 18736 35678
rect 19996 34134 20024 35678
rect 19984 34128 20036 34134
rect 19984 34070 20036 34076
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 18696 33448 18748 33454
rect 18696 33390 18748 33396
rect 18604 33312 18656 33318
rect 19064 33312 19116 33318
rect 18604 33254 18656 33260
rect 19062 33280 19064 33289
rect 19116 33280 19118 33289
rect 18616 32298 18644 33254
rect 19062 33215 19118 33224
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 18786 32328 18842 32337
rect 18604 32292 18656 32298
rect 18786 32263 18842 32272
rect 18604 32234 18656 32240
rect 18800 32230 18828 32263
rect 18788 32224 18840 32230
rect 18788 32166 18840 32172
rect 18800 31958 18828 32166
rect 18892 32026 18920 32846
rect 19616 32768 19668 32774
rect 19616 32710 19668 32716
rect 19628 32502 19656 32710
rect 19616 32496 19668 32502
rect 19616 32438 19668 32444
rect 19720 32434 19748 33458
rect 21284 33454 21312 35678
rect 22572 34202 22600 35678
rect 22988 34300 23296 34309
rect 22988 34298 22994 34300
rect 23050 34298 23074 34300
rect 23130 34298 23154 34300
rect 23210 34298 23234 34300
rect 23290 34298 23296 34300
rect 23050 34246 23052 34298
rect 23232 34246 23234 34298
rect 22988 34244 22994 34246
rect 23050 34244 23074 34246
rect 23130 34244 23154 34246
rect 23210 34244 23234 34246
rect 23290 34244 23296 34246
rect 22988 34235 23296 34244
rect 22560 34196 22612 34202
rect 22560 34138 22612 34144
rect 23860 34134 23888 35678
rect 23848 34128 23900 34134
rect 23848 34070 23900 34076
rect 22100 34060 22152 34066
rect 22100 34002 22152 34008
rect 24124 34060 24176 34066
rect 24124 34002 24176 34008
rect 21272 33448 21324 33454
rect 21272 33390 21324 33396
rect 21548 33312 21600 33318
rect 21546 33280 21548 33289
rect 21600 33280 21602 33289
rect 21546 33215 21602 33224
rect 19708 32428 19760 32434
rect 19708 32370 19760 32376
rect 19800 32428 19852 32434
rect 19800 32370 19852 32376
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 18788 31952 18840 31958
rect 18788 31894 18840 31900
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 18420 31476 18472 31482
rect 18420 31418 18472 31424
rect 18144 31204 18196 31210
rect 18144 31146 18196 31152
rect 18156 30734 18184 31146
rect 18432 30938 18460 31418
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18800 30938 18828 31282
rect 18420 30932 18472 30938
rect 18420 30874 18472 30880
rect 18788 30932 18840 30938
rect 18788 30874 18840 30880
rect 17868 30728 17920 30734
rect 17868 30670 17920 30676
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 19168 30598 19196 31826
rect 19720 31754 19748 32370
rect 19812 32026 19840 32370
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19720 31726 19840 31754
rect 19708 30728 19760 30734
rect 19708 30670 19760 30676
rect 17868 30592 17920 30598
rect 17868 30534 17920 30540
rect 19156 30592 19208 30598
rect 19156 30534 19208 30540
rect 17604 29158 17724 29186
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17512 28218 17540 28358
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17224 27600 17276 27606
rect 17224 27542 17276 27548
rect 17236 27470 17264 27542
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 17236 26858 17264 27406
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 17604 26586 17632 29158
rect 17684 29096 17736 29102
rect 17684 29038 17736 29044
rect 17696 28014 17724 29038
rect 17684 28008 17736 28014
rect 17684 27950 17736 27956
rect 17696 26994 17724 27950
rect 17776 27872 17828 27878
rect 17776 27814 17828 27820
rect 17788 27674 17816 27814
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 17684 26988 17736 26994
rect 17684 26930 17736 26936
rect 17592 26580 17644 26586
rect 17592 26522 17644 26528
rect 17604 26364 17632 26522
rect 17406 26344 17462 26353
rect 17406 26279 17408 26288
rect 17460 26279 17462 26288
rect 17512 26336 17632 26364
rect 17408 26250 17460 26256
rect 17132 26240 17184 26246
rect 17132 26182 17184 26188
rect 17144 25838 17172 26182
rect 17408 25968 17460 25974
rect 17408 25910 17460 25916
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 17144 22094 17172 25774
rect 17420 25430 17448 25910
rect 17408 25424 17460 25430
rect 17408 25366 17460 25372
rect 17316 24336 17368 24342
rect 17316 24278 17368 24284
rect 17328 23526 17356 24278
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 17236 22234 17264 22510
rect 17224 22228 17276 22234
rect 17224 22170 17276 22176
rect 17144 22066 17264 22094
rect 17130 21584 17186 21593
rect 17130 21519 17132 21528
rect 17184 21519 17186 21528
rect 17132 21490 17184 21496
rect 17130 20496 17186 20505
rect 17130 20431 17186 20440
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16684 18426 16712 18702
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16776 18222 16804 18566
rect 16764 18216 16816 18222
rect 16764 18158 16816 18164
rect 16948 18216 17000 18222
rect 16948 18158 17000 18164
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16856 17672 16908 17678
rect 16856 17614 16908 17620
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16488 16720 16540 16726
rect 16488 16662 16540 16668
rect 16500 16454 16528 16662
rect 16488 16448 16540 16454
rect 16488 16390 16540 16396
rect 16500 15994 16528 16390
rect 16592 16114 16620 16730
rect 16580 16108 16632 16114
rect 16580 16050 16632 16056
rect 16500 15966 16620 15994
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16500 15026 16528 15302
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16408 13462 16436 14554
rect 16500 14482 16528 14962
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16396 13456 16448 13462
rect 16302 13424 16358 13433
rect 16396 13398 16448 13404
rect 16500 13394 16528 13670
rect 16302 13359 16358 13368
rect 16488 13388 16540 13394
rect 16316 12986 16344 13359
rect 16488 13330 16540 13336
rect 16592 13274 16620 15966
rect 16684 14958 16712 17478
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16776 16250 16804 16526
rect 16764 16244 16816 16250
rect 16764 16186 16816 16192
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16776 15366 16804 15914
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16764 15088 16816 15094
rect 16764 15030 16816 15036
rect 16672 14952 16724 14958
rect 16672 14894 16724 14900
rect 16776 13938 16804 15030
rect 16764 13932 16816 13938
rect 16764 13874 16816 13880
rect 16868 13818 16896 17614
rect 16960 16658 16988 18158
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17052 16046 17080 19654
rect 17144 19310 17172 20431
rect 17236 19854 17264 22066
rect 17224 19848 17276 19854
rect 17224 19790 17276 19796
rect 17236 19514 17264 19790
rect 17328 19718 17356 23462
rect 17408 23112 17460 23118
rect 17408 23054 17460 23060
rect 17420 22030 17448 23054
rect 17512 22098 17540 26336
rect 17696 25906 17724 26930
rect 17880 26450 17908 30534
rect 17960 29028 18012 29034
rect 17960 28970 18012 28976
rect 17972 28762 18000 28970
rect 17960 28756 18012 28762
rect 17960 28698 18012 28704
rect 19168 28694 19196 30534
rect 19720 29306 19748 30670
rect 19708 29300 19760 29306
rect 19708 29242 19760 29248
rect 19812 29186 19840 31726
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 19720 29158 19840 29186
rect 19720 29102 19748 29158
rect 19708 29096 19760 29102
rect 19708 29038 19760 29044
rect 19156 28688 19208 28694
rect 19156 28630 19208 28636
rect 19708 28688 19760 28694
rect 19708 28630 19760 28636
rect 19248 28620 19300 28626
rect 19248 28562 19300 28568
rect 19616 28620 19668 28626
rect 19616 28562 19668 28568
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 18064 27674 18092 27814
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 19064 27600 19116 27606
rect 19064 27542 19116 27548
rect 18972 27328 19024 27334
rect 18972 27270 19024 27276
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 17880 25906 17908 26386
rect 18064 26314 18092 26930
rect 18984 26450 19012 27270
rect 19076 27130 19104 27542
rect 19260 27470 19288 28562
rect 19628 28121 19656 28562
rect 19614 28112 19670 28121
rect 19444 28070 19614 28098
rect 19248 27464 19300 27470
rect 19248 27406 19300 27412
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 18972 26444 19024 26450
rect 18972 26386 19024 26392
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18052 26308 18104 26314
rect 18052 26250 18104 26256
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17696 25498 17724 25842
rect 18064 25838 18092 26250
rect 18052 25832 18104 25838
rect 18052 25774 18104 25780
rect 17776 25696 17828 25702
rect 17776 25638 17828 25644
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 17788 25294 17816 25638
rect 17776 25288 17828 25294
rect 17776 25230 17828 25236
rect 17592 24608 17644 24614
rect 17592 24550 17644 24556
rect 17604 24290 17632 24550
rect 17604 24262 17724 24290
rect 17592 24132 17644 24138
rect 17592 24074 17644 24080
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 17408 22024 17460 22030
rect 17408 21966 17460 21972
rect 17604 21962 17632 24074
rect 17592 21956 17644 21962
rect 17592 21898 17644 21904
rect 17696 21672 17724 24262
rect 18052 24064 18104 24070
rect 18052 24006 18104 24012
rect 17868 23588 17920 23594
rect 17868 23530 17920 23536
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17788 22234 17816 22918
rect 17880 22778 17908 23530
rect 18064 23526 18092 24006
rect 18052 23520 18104 23526
rect 18052 23462 18104 23468
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17776 22228 17828 22234
rect 17776 22170 17828 22176
rect 17880 22094 17908 22510
rect 17960 22432 18012 22438
rect 17960 22374 18012 22380
rect 17512 21644 17724 21672
rect 17788 22066 17908 22094
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17224 19508 17276 19514
rect 17276 19468 17356 19496
rect 17224 19450 17276 19456
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 17328 18290 17356 19468
rect 17420 18902 17448 19654
rect 17512 18970 17540 21644
rect 17788 18986 17816 22066
rect 17972 21894 18000 22374
rect 17868 21888 17920 21894
rect 17868 21830 17920 21836
rect 17960 21888 18012 21894
rect 17960 21830 18012 21836
rect 17880 21622 17908 21830
rect 17868 21616 17920 21622
rect 17868 21558 17920 21564
rect 17972 21146 18000 21830
rect 18156 21690 18184 26318
rect 18970 25800 19026 25809
rect 18880 25764 18932 25770
rect 18970 25735 18972 25744
rect 18880 25706 18932 25712
rect 19024 25735 19026 25744
rect 18972 25706 19024 25712
rect 18512 25696 18564 25702
rect 18512 25638 18564 25644
rect 18524 25226 18552 25638
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18696 25288 18748 25294
rect 18696 25230 18748 25236
rect 18512 25220 18564 25226
rect 18512 25162 18564 25168
rect 18616 24954 18644 25230
rect 18236 24948 18288 24954
rect 18236 24890 18288 24896
rect 18604 24948 18656 24954
rect 18604 24890 18656 24896
rect 18248 24206 18276 24890
rect 18512 24812 18564 24818
rect 18512 24754 18564 24760
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18248 22574 18276 24142
rect 18340 24070 18368 24550
rect 18432 24138 18460 24550
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18340 22778 18368 22918
rect 18328 22772 18380 22778
rect 18328 22714 18380 22720
rect 18432 22574 18460 23666
rect 18236 22568 18288 22574
rect 18236 22510 18288 22516
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 18328 22160 18380 22166
rect 18380 22120 18460 22148
rect 18328 22102 18380 22108
rect 18432 21894 18460 22120
rect 18236 21888 18288 21894
rect 18236 21830 18288 21836
rect 18420 21888 18472 21894
rect 18420 21830 18472 21836
rect 18144 21684 18196 21690
rect 18144 21626 18196 21632
rect 17960 21140 18012 21146
rect 17960 21082 18012 21088
rect 17960 20868 18012 20874
rect 17960 20810 18012 20816
rect 17972 20398 18000 20810
rect 18144 20800 18196 20806
rect 18144 20742 18196 20748
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17868 20256 17920 20262
rect 17868 20198 17920 20204
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17604 18958 17816 18986
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17316 18284 17368 18290
rect 17368 18244 17448 18272
rect 17316 18226 17368 18232
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17224 18080 17276 18086
rect 17224 18022 17276 18028
rect 17144 17542 17172 18022
rect 17236 17678 17264 18022
rect 17420 17814 17448 18244
rect 17408 17808 17460 17814
rect 17408 17750 17460 17756
rect 17604 17678 17632 18958
rect 17776 18624 17828 18630
rect 17776 18566 17828 18572
rect 17788 18290 17816 18566
rect 17880 18290 17908 20198
rect 17972 19922 18000 20334
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 18064 19802 18092 20402
rect 17972 19774 18092 19802
rect 17972 19718 18000 19774
rect 17960 19712 18012 19718
rect 17960 19654 18012 19660
rect 17776 18284 17828 18290
rect 17776 18226 17828 18232
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17592 17672 17644 17678
rect 17592 17614 17644 17620
rect 17132 17536 17184 17542
rect 17132 17478 17184 17484
rect 17604 17134 17632 17614
rect 17696 17610 17724 18022
rect 17788 17814 17816 18226
rect 17880 17814 17908 18226
rect 17776 17808 17828 17814
rect 17776 17750 17828 17756
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17592 17128 17644 17134
rect 17592 17070 17644 17076
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16114 17540 16934
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17052 15586 17080 15982
rect 17408 15632 17460 15638
rect 17052 15558 17172 15586
rect 17408 15574 17460 15580
rect 17040 15496 17092 15502
rect 17144 15484 17172 15558
rect 17224 15496 17276 15502
rect 17144 15456 17224 15484
rect 17040 15438 17092 15444
rect 17224 15438 17276 15444
rect 16948 14952 17000 14958
rect 16948 14894 17000 14900
rect 16960 13938 16988 14894
rect 17052 14074 17080 15438
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17144 14618 17172 14962
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17328 14618 17356 14758
rect 17420 14618 17448 15574
rect 17132 14612 17184 14618
rect 17132 14554 17184 14560
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17224 14340 17276 14346
rect 17224 14282 17276 14288
rect 17236 14074 17264 14282
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 17224 14068 17276 14074
rect 17224 14010 17276 14016
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16500 13246 16620 13274
rect 16684 13790 16896 13818
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16316 12102 16344 12718
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16316 11830 16344 12038
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16500 10674 16528 13246
rect 16580 13184 16632 13190
rect 16578 13152 16580 13161
rect 16632 13152 16634 13161
rect 16578 13087 16634 13096
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16592 12374 16620 12718
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16684 11286 16712 13790
rect 16856 13728 16908 13734
rect 17132 13728 17184 13734
rect 16856 13670 16908 13676
rect 16960 13688 17132 13716
rect 16764 13388 16816 13394
rect 16764 13330 16816 13336
rect 16776 12986 16804 13330
rect 16868 13326 16896 13670
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16854 13016 16910 13025
rect 16764 12980 16816 12986
rect 16854 12951 16856 12960
rect 16764 12922 16816 12928
rect 16908 12951 16910 12960
rect 16856 12922 16908 12928
rect 16960 12782 16988 13688
rect 17132 13670 17184 13676
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17144 13161 17172 13262
rect 17130 13152 17186 13161
rect 17130 13087 17186 13096
rect 16764 12776 16816 12782
rect 16764 12718 16816 12724
rect 16948 12776 17000 12782
rect 16948 12718 17000 12724
rect 16776 12628 16804 12718
rect 17040 12640 17092 12646
rect 16776 12600 16896 12628
rect 16868 12374 16896 12600
rect 17040 12582 17092 12588
rect 16856 12368 16908 12374
rect 16856 12310 16908 12316
rect 17052 11762 17080 12582
rect 17144 12374 17172 13087
rect 17132 12368 17184 12374
rect 17132 12310 17184 12316
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17144 11676 17172 12310
rect 17236 12170 17264 14010
rect 17420 14006 17448 14554
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17408 14000 17460 14006
rect 17408 13942 17460 13948
rect 17512 13530 17540 14418
rect 17604 13870 17632 16594
rect 17696 16250 17724 17546
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17880 17134 17908 17478
rect 17868 17128 17920 17134
rect 17868 17070 17920 17076
rect 17684 16244 17736 16250
rect 17684 16186 17736 16192
rect 17684 15632 17736 15638
rect 17684 15574 17736 15580
rect 17696 14958 17724 15574
rect 17972 15162 18000 19654
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 18064 15570 18092 18022
rect 18156 17649 18184 20742
rect 18248 19786 18276 21830
rect 18328 20868 18380 20874
rect 18328 20810 18380 20816
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 18340 19718 18368 20810
rect 18432 19854 18460 21830
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18142 17640 18198 17649
rect 18142 17575 18198 17584
rect 18248 17320 18276 17682
rect 18340 17678 18368 19654
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18432 17542 18460 19790
rect 18524 18834 18552 24754
rect 18708 24750 18736 25230
rect 18892 24750 18920 25706
rect 19076 25242 19104 26794
rect 19260 26466 19288 27406
rect 19168 26438 19288 26466
rect 19168 25838 19196 26438
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19260 26042 19288 26318
rect 19248 26036 19300 26042
rect 19248 25978 19300 25984
rect 19156 25832 19208 25838
rect 19156 25774 19208 25780
rect 19168 25362 19196 25774
rect 19156 25356 19208 25362
rect 19208 25316 19380 25344
rect 19156 25298 19208 25304
rect 19076 25214 19196 25242
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18880 24744 18932 24750
rect 18880 24686 18932 24692
rect 18604 24676 18656 24682
rect 18604 24618 18656 24624
rect 18616 24410 18644 24618
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18972 24064 19024 24070
rect 18972 24006 19024 24012
rect 18604 23792 18656 23798
rect 18604 23734 18656 23740
rect 18616 21026 18644 23734
rect 18696 23180 18748 23186
rect 18696 23122 18748 23128
rect 18708 21962 18736 23122
rect 18984 22386 19012 24006
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 19076 22506 19104 23462
rect 19168 23118 19196 25214
rect 19352 23798 19380 25316
rect 19444 24750 19472 28070
rect 19614 28047 19670 28056
rect 19524 25696 19576 25702
rect 19524 25638 19576 25644
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 19536 25362 19564 25638
rect 19628 25498 19656 25638
rect 19616 25492 19668 25498
rect 19616 25434 19668 25440
rect 19524 25356 19576 25362
rect 19524 25298 19576 25304
rect 19432 24744 19484 24750
rect 19432 24686 19484 24692
rect 19536 24698 19564 25298
rect 19616 25152 19668 25158
rect 19616 25094 19668 25100
rect 19628 24818 19656 25094
rect 19616 24812 19668 24818
rect 19616 24754 19668 24760
rect 19720 24750 19748 28630
rect 20076 28008 20128 28014
rect 20074 27976 20076 27985
rect 20128 27976 20130 27985
rect 20074 27911 20130 27920
rect 20088 27674 20116 27911
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 20272 27334 20300 29582
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 20904 28960 20956 28966
rect 20904 28902 20956 28908
rect 20916 28218 20944 28902
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 20904 28212 20956 28218
rect 20904 28154 20956 28160
rect 20916 28014 20944 28154
rect 20904 28008 20956 28014
rect 20904 27950 20956 27956
rect 20260 27328 20312 27334
rect 20260 27270 20312 27276
rect 20916 26926 20944 27950
rect 20996 27872 21048 27878
rect 20996 27814 21048 27820
rect 21008 27606 21036 27814
rect 20996 27600 21048 27606
rect 20996 27542 21048 27548
rect 21100 27470 21128 28562
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 21100 26926 21128 27406
rect 21192 26926 21220 29446
rect 21272 29028 21324 29034
rect 21272 28970 21324 28976
rect 21548 29028 21600 29034
rect 21548 28970 21600 28976
rect 21284 27334 21312 28970
rect 21560 28762 21588 28970
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21916 28688 21968 28694
rect 21916 28630 21968 28636
rect 21928 27878 21956 28630
rect 21916 27872 21968 27878
rect 21916 27814 21968 27820
rect 21824 27600 21876 27606
rect 21824 27542 21876 27548
rect 21732 27464 21784 27470
rect 21732 27406 21784 27412
rect 21272 27328 21324 27334
rect 21272 27270 21324 27276
rect 21744 27130 21772 27406
rect 21836 27130 21864 27542
rect 21732 27124 21784 27130
rect 21732 27066 21784 27072
rect 21824 27124 21876 27130
rect 21824 27066 21876 27072
rect 21928 26994 21956 27814
rect 22008 27328 22060 27334
rect 22008 27270 22060 27276
rect 22020 27130 22048 27270
rect 22008 27124 22060 27130
rect 22008 27066 22060 27072
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 20904 26920 20956 26926
rect 20904 26862 20956 26868
rect 21088 26920 21140 26926
rect 21088 26862 21140 26868
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21364 26920 21416 26926
rect 21364 26862 21416 26868
rect 20916 26382 20944 26862
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20628 25696 20680 25702
rect 20628 25638 20680 25644
rect 19984 25492 20036 25498
rect 19984 25434 20036 25440
rect 19708 24744 19760 24750
rect 19536 24670 19656 24698
rect 19708 24686 19760 24692
rect 19628 24614 19656 24670
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 19524 24268 19576 24274
rect 19524 24210 19576 24216
rect 19340 23792 19392 23798
rect 19340 23734 19392 23740
rect 19352 23610 19380 23734
rect 19260 23582 19380 23610
rect 19260 23186 19288 23582
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19156 23112 19208 23118
rect 19156 23054 19208 23060
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 18984 22358 19104 22386
rect 18880 22092 18932 22098
rect 18880 22034 18932 22040
rect 18696 21956 18748 21962
rect 18696 21898 18748 21904
rect 18788 21888 18840 21894
rect 18788 21830 18840 21836
rect 18800 21486 18828 21830
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18616 20998 18736 21026
rect 18604 20936 18656 20942
rect 18604 20878 18656 20884
rect 18616 20602 18644 20878
rect 18708 20806 18736 20998
rect 18696 20800 18748 20806
rect 18696 20742 18748 20748
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18708 19922 18736 20742
rect 18696 19916 18748 19922
rect 18696 19858 18748 19864
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18800 18358 18828 21286
rect 18892 20398 18920 22034
rect 19076 22030 19104 22358
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 18984 21486 19012 21966
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18880 20392 18932 20398
rect 18880 20334 18932 20340
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18892 19938 18920 20198
rect 18984 20058 19012 21422
rect 19076 21350 19104 21966
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19076 20369 19104 20538
rect 19168 20466 19196 23054
rect 19352 22982 19380 23462
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19156 20460 19208 20466
rect 19156 20402 19208 20408
rect 19062 20360 19118 20369
rect 19062 20295 19118 20304
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 18892 19910 19012 19938
rect 19168 19922 19196 19994
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18788 18352 18840 18358
rect 18786 18320 18788 18329
rect 18840 18320 18842 18329
rect 18696 18284 18748 18290
rect 18786 18255 18842 18264
rect 18696 18226 18748 18232
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18604 18216 18656 18222
rect 18604 18158 18656 18164
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18340 17338 18368 17478
rect 18156 17292 18276 17320
rect 18328 17332 18380 17338
rect 18156 17202 18184 17292
rect 18328 17274 18380 17280
rect 18432 17218 18460 17478
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18248 17190 18460 17218
rect 18156 17105 18184 17138
rect 18142 17096 18198 17105
rect 18142 17031 18198 17040
rect 18144 16992 18196 16998
rect 18248 16980 18276 17190
rect 18524 17134 18552 18158
rect 18616 18086 18644 18158
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18616 17134 18644 18022
rect 18708 17202 18736 18226
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18800 17338 18828 18158
rect 18892 17882 18920 19314
rect 18984 18222 19012 19910
rect 19156 19916 19208 19922
rect 19156 19858 19208 19864
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19076 18426 19104 19790
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19260 19378 19288 19722
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19352 19334 19380 22918
rect 19536 21622 19564 24210
rect 19628 23662 19656 24550
rect 19616 23656 19668 23662
rect 19616 23598 19668 23604
rect 19720 23322 19748 24686
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19904 23662 19932 24006
rect 19892 23656 19944 23662
rect 19892 23598 19944 23604
rect 19800 23588 19852 23594
rect 19800 23530 19852 23536
rect 19708 23316 19760 23322
rect 19708 23258 19760 23264
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19628 22030 19656 22714
rect 19708 22500 19760 22506
rect 19708 22442 19760 22448
rect 19616 22024 19668 22030
rect 19616 21966 19668 21972
rect 19524 21616 19576 21622
rect 19524 21558 19576 21564
rect 19536 21350 19564 21558
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19628 21146 19656 21966
rect 19720 21894 19748 22442
rect 19708 21888 19760 21894
rect 19708 21830 19760 21836
rect 19616 21140 19668 21146
rect 19616 21082 19668 21088
rect 19720 20777 19748 21830
rect 19706 20768 19762 20777
rect 19706 20703 19762 20712
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19444 19990 19472 20334
rect 19432 19984 19484 19990
rect 19432 19926 19484 19932
rect 19352 19306 19656 19334
rect 19432 18964 19484 18970
rect 19432 18906 19484 18912
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19156 18828 19208 18834
rect 19444 18816 19472 18906
rect 19536 18873 19564 18906
rect 19156 18770 19208 18776
rect 19260 18788 19472 18816
rect 19522 18864 19578 18873
rect 19522 18799 19578 18808
rect 19064 18420 19116 18426
rect 19064 18362 19116 18368
rect 19076 18290 19104 18362
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18972 18216 19024 18222
rect 18972 18158 19024 18164
rect 18880 17876 18932 17882
rect 18880 17818 18932 17824
rect 19064 17740 19116 17746
rect 19064 17682 19116 17688
rect 18788 17332 18840 17338
rect 18788 17274 18840 17280
rect 18696 17196 18748 17202
rect 18696 17138 18748 17144
rect 18328 17128 18380 17134
rect 18328 17070 18380 17076
rect 18512 17128 18564 17134
rect 18512 17070 18564 17076
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18196 16952 18276 16980
rect 18340 16980 18368 17070
rect 18340 16952 18552 16980
rect 18144 16934 18196 16940
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18156 15706 18184 16390
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 17868 15156 17920 15162
rect 17868 15098 17920 15104
rect 17960 15156 18012 15162
rect 17960 15098 18012 15104
rect 17880 15042 17908 15098
rect 18144 15088 18196 15094
rect 17880 15014 18000 15042
rect 18144 15030 18196 15036
rect 17972 14958 18000 15014
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17960 14952 18012 14958
rect 17960 14894 18012 14900
rect 17696 14113 17724 14894
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17776 14476 17828 14482
rect 17776 14418 17828 14424
rect 17868 14476 17920 14482
rect 17868 14418 17920 14424
rect 17682 14104 17738 14113
rect 17682 14039 17738 14048
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17590 13696 17646 13705
rect 17590 13631 17646 13640
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17314 13424 17370 13433
rect 17314 13359 17370 13368
rect 17408 13388 17460 13394
rect 17328 13326 17356 13359
rect 17408 13330 17460 13336
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17420 13274 17448 13330
rect 17420 13246 17540 13274
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17328 12986 17356 13126
rect 17316 12980 17368 12986
rect 17512 12968 17540 13246
rect 17316 12922 17368 12928
rect 17420 12940 17540 12968
rect 17420 12866 17448 12940
rect 17604 12866 17632 13631
rect 17696 13530 17724 14039
rect 17684 13524 17736 13530
rect 17684 13466 17736 13472
rect 17788 13394 17816 14418
rect 17776 13388 17828 13394
rect 17776 13330 17828 13336
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 12918 17724 13262
rect 17328 12838 17448 12866
rect 17512 12838 17632 12866
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17224 12164 17276 12170
rect 17224 12106 17276 12112
rect 17224 11688 17276 11694
rect 17144 11648 17224 11676
rect 17224 11630 17276 11636
rect 16672 11280 16724 11286
rect 16672 11222 16724 11228
rect 16684 10810 16712 11222
rect 17236 11014 17264 11630
rect 17328 11150 17356 12838
rect 17406 12744 17462 12753
rect 17406 12679 17462 12688
rect 17420 12646 17448 12679
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17406 11928 17462 11937
rect 17406 11863 17462 11872
rect 17420 11830 17448 11863
rect 17408 11824 17460 11830
rect 17408 11766 17460 11772
rect 17512 11558 17540 12838
rect 17592 12776 17644 12782
rect 17644 12724 17724 12730
rect 17592 12718 17724 12724
rect 17604 12702 17724 12718
rect 17788 12714 17816 13330
rect 17880 13258 17908 14418
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17972 13025 18000 14554
rect 18052 14272 18104 14278
rect 18052 14214 18104 14220
rect 18064 13802 18092 14214
rect 18052 13796 18104 13802
rect 18052 13738 18104 13744
rect 18064 13462 18092 13738
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17958 13016 18014 13025
rect 18064 12986 18092 13398
rect 18156 12986 18184 15030
rect 17958 12951 18014 12960
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11218 17540 11494
rect 17590 11248 17646 11257
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17500 11212 17552 11218
rect 17590 11183 17592 11192
rect 17500 11154 17552 11160
rect 17644 11183 17646 11192
rect 17592 11154 17644 11160
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17040 11008 17092 11014
rect 16946 10976 17002 10985
rect 17040 10950 17092 10956
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 16946 10911 17002 10920
rect 16960 10810 16988 10911
rect 16672 10804 16724 10810
rect 16672 10746 16724 10752
rect 16948 10804 17000 10810
rect 16948 10746 17000 10752
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15764 10062 15792 10406
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15764 9722 15792 9998
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15764 9382 15792 9658
rect 15856 9586 15884 10406
rect 16316 10266 16344 10542
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 16580 9580 16632 9586
rect 16684 9568 16712 10746
rect 16960 10062 16988 10746
rect 17052 10266 17080 10950
rect 17420 10606 17448 11154
rect 17512 11098 17540 11154
rect 17512 11070 17632 11098
rect 17408 10600 17460 10606
rect 17408 10542 17460 10548
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 16632 9540 16712 9568
rect 16580 9522 16632 9528
rect 16684 9382 16712 9540
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 15764 8090 15792 9318
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 15948 8498 15976 8774
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15752 8084 15804 8090
rect 15752 8026 15804 8032
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15764 7546 15792 7822
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15948 7342 15976 8434
rect 16592 8362 16620 8774
rect 16684 8498 16712 9318
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16776 8090 16804 9386
rect 16868 8906 16896 9998
rect 17052 9722 17080 9998
rect 17040 9716 17092 9722
rect 17040 9658 17092 9664
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16856 8900 16908 8906
rect 16856 8842 16908 8848
rect 16960 8566 16988 8910
rect 17132 8900 17184 8906
rect 17132 8842 17184 8848
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 17144 8498 17172 8842
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17144 8090 17172 8434
rect 17236 8430 17264 10134
rect 17420 9994 17448 10542
rect 17604 10470 17632 11070
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17408 9988 17460 9994
rect 17408 9930 17460 9936
rect 17420 9674 17448 9930
rect 17420 9646 17540 9674
rect 17420 9518 17448 9646
rect 17408 9512 17460 9518
rect 17512 9489 17540 9646
rect 17604 9518 17632 10406
rect 17696 10062 17724 12702
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17868 12368 17920 12374
rect 18050 12336 18106 12345
rect 17868 12310 17920 12316
rect 17880 12102 17908 12310
rect 17972 12294 18050 12322
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 9654 17724 9998
rect 17684 9648 17736 9654
rect 17684 9590 17736 9596
rect 17592 9512 17644 9518
rect 17408 9454 17460 9460
rect 17498 9480 17554 9489
rect 17592 9454 17644 9460
rect 17498 9415 17554 9424
rect 17604 9382 17632 9454
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17604 9042 17632 9318
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 16672 7948 16724 7954
rect 16672 7890 16724 7896
rect 16684 7546 16712 7890
rect 17236 7886 17264 8366
rect 17696 8294 17724 9590
rect 17788 8498 17816 10542
rect 17866 9480 17922 9489
rect 17866 9415 17922 9424
rect 17880 9110 17908 9415
rect 17868 9104 17920 9110
rect 17868 9046 17920 9052
rect 17972 8514 18000 12294
rect 18050 12271 18106 12280
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18064 11801 18092 12174
rect 18050 11792 18106 11801
rect 18050 11727 18106 11736
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10266 18092 10950
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18144 9444 18196 9450
rect 18144 9386 18196 9392
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 18064 9081 18092 9114
rect 18050 9072 18106 9081
rect 18050 9007 18106 9016
rect 18156 8838 18184 9386
rect 18144 8832 18196 8838
rect 18144 8774 18196 8780
rect 17776 8492 17828 8498
rect 17972 8486 18092 8514
rect 17776 8434 17828 8440
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 16672 7540 16724 7546
rect 16672 7482 16724 7488
rect 16776 7342 16804 7686
rect 17328 7546 17356 7822
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17420 7410 17448 8230
rect 17696 8022 17724 8230
rect 17788 8022 17816 8434
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17972 8090 18000 8366
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17776 8016 17828 8022
rect 17776 7958 17828 7964
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 15948 6934 15976 7278
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15099 6012 15407 6021
rect 15099 6010 15105 6012
rect 15161 6010 15185 6012
rect 15241 6010 15265 6012
rect 15321 6010 15345 6012
rect 15401 6010 15407 6012
rect 15161 5958 15163 6010
rect 15343 5958 15345 6010
rect 15099 5956 15105 5958
rect 15161 5956 15185 5958
rect 15241 5956 15265 5958
rect 15321 5956 15345 5958
rect 15401 5956 15407 5958
rect 15099 5947 15407 5956
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 15028 5370 15056 5646
rect 15672 5370 15700 6190
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 16040 5250 16068 5306
rect 15948 5222 16068 5250
rect 16316 5234 16344 6734
rect 16592 6322 16620 6802
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16776 5778 16804 7278
rect 16960 6798 16988 7278
rect 18064 6866 18092 8486
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18156 8090 18184 8434
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 16948 6792 17000 6798
rect 16948 6734 17000 6740
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16670 5672 16726 5681
rect 16670 5607 16726 5616
rect 16396 5568 16448 5574
rect 16396 5510 16448 5516
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16304 5228 16356 5234
rect 14832 5160 14884 5166
rect 14832 5102 14884 5108
rect 14439 4380 14747 4389
rect 14439 4378 14445 4380
rect 14501 4378 14525 4380
rect 14581 4378 14605 4380
rect 14661 4378 14685 4380
rect 14741 4378 14747 4380
rect 14501 4326 14503 4378
rect 14683 4326 14685 4378
rect 14439 4324 14445 4326
rect 14501 4324 14525 4326
rect 14581 4324 14605 4326
rect 14661 4324 14685 4326
rect 14741 4324 14747 4326
rect 14439 4315 14747 4324
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14660 3738 14688 4082
rect 14844 4010 14872 5102
rect 15099 4924 15407 4933
rect 15099 4922 15105 4924
rect 15161 4922 15185 4924
rect 15241 4922 15265 4924
rect 15321 4922 15345 4924
rect 15401 4922 15407 4924
rect 15161 4870 15163 4922
rect 15343 4870 15345 4922
rect 15099 4868 15105 4870
rect 15161 4868 15185 4870
rect 15241 4868 15265 4870
rect 15321 4868 15345 4870
rect 15401 4868 15407 4870
rect 15099 4859 15407 4868
rect 15948 4826 15976 5222
rect 16304 5170 16356 5176
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 15936 4820 15988 4826
rect 15936 4762 15988 4768
rect 16316 4758 16344 4966
rect 15292 4752 15344 4758
rect 15292 4694 15344 4700
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4146 15240 4422
rect 15304 4282 15332 4694
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 15099 3836 15407 3845
rect 15099 3834 15105 3836
rect 15161 3834 15185 3836
rect 15241 3834 15265 3836
rect 15321 3834 15345 3836
rect 15401 3834 15407 3836
rect 15161 3782 15163 3834
rect 15343 3782 15345 3834
rect 15099 3780 15105 3782
rect 15161 3780 15185 3782
rect 15241 3780 15265 3782
rect 15321 3780 15345 3782
rect 15401 3780 15407 3782
rect 15099 3771 15407 3780
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 16408 3602 16436 5510
rect 16592 5234 16620 5510
rect 16580 5228 16632 5234
rect 16580 5170 16632 5176
rect 16684 5166 16712 5607
rect 16868 5234 16896 6258
rect 16960 6254 16988 6734
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16960 5914 16988 6190
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17972 5914 18000 6122
rect 16948 5908 17000 5914
rect 16948 5850 17000 5856
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16764 4616 16816 4622
rect 16764 4558 16816 4564
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 14439 3292 14747 3301
rect 14439 3290 14445 3292
rect 14501 3290 14525 3292
rect 14581 3290 14605 3292
rect 14661 3290 14685 3292
rect 14741 3290 14747 3292
rect 14501 3238 14503 3290
rect 14683 3238 14685 3290
rect 14439 3236 14445 3238
rect 14501 3236 14525 3238
rect 14581 3236 14605 3238
rect 14661 3236 14685 3238
rect 14741 3236 14747 3238
rect 14439 3227 14747 3236
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13648 2774 13676 2926
rect 13556 2746 13676 2774
rect 13556 800 13584 2746
rect 14844 800 14872 2994
rect 15099 2748 15407 2757
rect 15099 2746 15105 2748
rect 15161 2746 15185 2748
rect 15241 2746 15265 2748
rect 15321 2746 15345 2748
rect 15401 2746 15407 2748
rect 15161 2694 15163 2746
rect 15343 2694 15345 2746
rect 15099 2692 15105 2694
rect 15161 2692 15185 2694
rect 15241 2692 15265 2694
rect 15321 2692 15345 2694
rect 15401 2692 15407 2694
rect 15099 2683 15407 2692
rect 16132 800 16160 3470
rect 16776 2990 16804 4558
rect 16868 4282 16896 5170
rect 16960 4826 16988 5850
rect 17868 5772 17920 5778
rect 17868 5714 17920 5720
rect 17880 4826 17908 5714
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 17868 4820 17920 4826
rect 17868 4762 17920 4768
rect 17972 4486 18000 4966
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 18248 4078 18276 16952
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18432 16114 18460 16390
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 18420 15156 18472 15162
rect 18420 15098 18472 15104
rect 18328 14340 18380 14346
rect 18328 14282 18380 14288
rect 18340 11354 18368 14282
rect 18432 14074 18460 15098
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18432 12345 18460 14010
rect 18524 13802 18552 16952
rect 18616 16794 18644 17070
rect 18604 16788 18656 16794
rect 18604 16730 18656 16736
rect 18800 16454 18828 17070
rect 18788 16448 18840 16454
rect 18788 16390 18840 16396
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18892 15366 18920 15506
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18708 14958 18736 15030
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18708 14550 18736 14894
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18696 14544 18748 14550
rect 18616 14504 18696 14532
rect 18512 13796 18564 13802
rect 18512 13738 18564 13744
rect 18616 13394 18644 14504
rect 18696 14486 18748 14492
rect 18788 14544 18840 14550
rect 18788 14486 18840 14492
rect 18696 14272 18748 14278
rect 18696 14214 18748 14220
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18512 12640 18564 12646
rect 18512 12582 18564 12588
rect 18418 12336 18474 12345
rect 18418 12271 18474 12280
rect 18524 11898 18552 12582
rect 18616 12374 18644 12922
rect 18708 12753 18736 14214
rect 18800 14074 18828 14486
rect 18892 14346 18920 14826
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 19076 14090 19104 17682
rect 18984 14074 19104 14090
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18984 14068 19116 14074
rect 18984 14062 19064 14068
rect 18786 13832 18842 13841
rect 18842 13790 18920 13818
rect 18786 13767 18842 13776
rect 18788 13388 18840 13394
rect 18788 13330 18840 13336
rect 18694 12744 18750 12753
rect 18694 12679 18750 12688
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18708 11898 18736 12679
rect 18800 12102 18828 13330
rect 18892 12238 18920 13790
rect 18984 13705 19012 14062
rect 19064 14010 19116 14016
rect 19168 13852 19196 18770
rect 19260 17678 19288 18788
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19536 18057 19564 18566
rect 19522 18048 19578 18057
rect 19522 17983 19578 17992
rect 19522 17776 19578 17785
rect 19522 17711 19524 17720
rect 19576 17711 19578 17720
rect 19524 17682 19576 17688
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19248 16040 19300 16046
rect 19248 15982 19300 15988
rect 19260 15706 19288 15982
rect 19248 15700 19300 15706
rect 19248 15642 19300 15648
rect 19260 15337 19288 15642
rect 19352 15502 19380 16594
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 19444 15502 19472 15846
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19246 15328 19302 15337
rect 19246 15263 19302 15272
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19260 14006 19288 14758
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19352 13870 19380 15438
rect 19444 15162 19472 15438
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19340 13864 19392 13870
rect 19168 13824 19288 13852
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18970 13696 19026 13705
rect 18970 13631 19026 13640
rect 18972 12776 19024 12782
rect 18972 12718 19024 12724
rect 18984 12442 19012 12718
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18340 9926 18368 10066
rect 18328 9920 18380 9926
rect 18328 9862 18380 9868
rect 18708 9674 18736 11018
rect 18892 10810 18920 12174
rect 18984 11694 19012 12378
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18616 9646 18736 9674
rect 18616 9450 18644 9646
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18786 9072 18842 9081
rect 18786 9007 18788 9016
rect 18840 9007 18842 9016
rect 18788 8978 18840 8984
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18420 7744 18472 7750
rect 18420 7686 18472 7692
rect 18432 7342 18460 7686
rect 18420 7336 18472 7342
rect 18420 7278 18472 7284
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 18340 4690 18368 5646
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18236 4072 18288 4078
rect 18236 4014 18288 4020
rect 18524 3398 18552 8910
rect 18984 8838 19012 10542
rect 18972 8832 19024 8838
rect 18972 8774 19024 8780
rect 18984 8650 19012 8774
rect 18892 8634 19012 8650
rect 18880 8628 19012 8634
rect 18932 8622 19012 8628
rect 18880 8570 18932 8576
rect 18972 8560 19024 8566
rect 18972 8502 19024 8508
rect 18786 8256 18842 8265
rect 18786 8191 18842 8200
rect 18602 8120 18658 8129
rect 18602 8055 18658 8064
rect 18616 7818 18644 8055
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18604 7812 18656 7818
rect 18604 7754 18656 7760
rect 18616 5370 18644 7754
rect 18708 7002 18736 7890
rect 18800 7546 18828 8191
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18708 5574 18736 6190
rect 18800 6118 18828 6734
rect 18984 6254 19012 8502
rect 19076 7936 19104 13738
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19260 13682 19288 13824
rect 19340 13806 19392 13812
rect 19628 13784 19656 19306
rect 19720 17921 19748 20334
rect 19812 18970 19840 23530
rect 19996 23186 20024 25434
rect 20640 25294 20668 25638
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20548 24954 20576 25230
rect 20536 24948 20588 24954
rect 20536 24890 20588 24896
rect 20916 24818 20944 26318
rect 21180 25832 21232 25838
rect 21180 25774 21232 25780
rect 21272 25832 21324 25838
rect 21272 25774 21324 25780
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21008 25430 21036 25638
rect 20996 25424 21048 25430
rect 20996 25366 21048 25372
rect 20904 24812 20956 24818
rect 20904 24754 20956 24760
rect 21192 24750 21220 25774
rect 21284 25498 21312 25774
rect 21272 25492 21324 25498
rect 21272 25434 21324 25440
rect 21180 24744 21232 24750
rect 21180 24686 21232 24692
rect 20536 23656 20588 23662
rect 20536 23598 20588 23604
rect 21088 23656 21140 23662
rect 21088 23598 21140 23604
rect 20168 23520 20220 23526
rect 20168 23462 20220 23468
rect 20180 23254 20208 23462
rect 20352 23316 20404 23322
rect 20352 23258 20404 23264
rect 20168 23248 20220 23254
rect 20168 23190 20220 23196
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19996 22778 20024 23122
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 20364 22574 20392 23258
rect 20548 22574 20576 23598
rect 20996 23520 21048 23526
rect 20996 23462 21048 23468
rect 21008 23254 21036 23462
rect 20996 23248 21048 23254
rect 20996 23190 21048 23196
rect 21100 22574 21128 23598
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 21088 22568 21140 22574
rect 21088 22510 21140 22516
rect 21180 22568 21232 22574
rect 21180 22510 21232 22516
rect 20364 22094 20392 22510
rect 20180 22066 20392 22094
rect 19892 20596 19944 20602
rect 19892 20538 19944 20544
rect 19904 20262 19932 20538
rect 19984 20324 20036 20330
rect 19984 20266 20036 20272
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19904 19990 19932 20198
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19996 19854 20024 20266
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 19892 19712 19944 19718
rect 19892 19654 19944 19660
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19800 18828 19852 18834
rect 19800 18770 19852 18776
rect 19812 18358 19840 18770
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19706 17912 19762 17921
rect 19706 17847 19762 17856
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19812 17202 19840 17478
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19904 17082 19932 19654
rect 19812 17054 19932 17082
rect 19812 16046 19840 17054
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 19628 13756 19748 13784
rect 19168 13394 19196 13670
rect 19260 13654 19656 13682
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19168 12442 19196 13330
rect 19628 13258 19656 13654
rect 19616 13252 19668 13258
rect 19616 13194 19668 13200
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19260 12986 19288 13126
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19168 11762 19196 12378
rect 19246 11928 19302 11937
rect 19352 11898 19380 13126
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19536 12442 19564 12718
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19522 12336 19578 12345
rect 19522 12271 19524 12280
rect 19576 12271 19578 12280
rect 19524 12242 19576 12248
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19246 11863 19248 11872
rect 19300 11863 19302 11872
rect 19340 11892 19392 11898
rect 19248 11834 19300 11840
rect 19340 11834 19392 11840
rect 19156 11756 19208 11762
rect 19156 11698 19208 11704
rect 19444 11694 19472 12038
rect 19628 11694 19656 13194
rect 19432 11688 19484 11694
rect 19338 11656 19394 11665
rect 19432 11630 19484 11636
rect 19616 11688 19668 11694
rect 19616 11630 19668 11636
rect 19338 11591 19340 11600
rect 19392 11591 19394 11600
rect 19340 11562 19392 11568
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19168 10606 19196 11494
rect 19444 11218 19472 11630
rect 19432 11212 19484 11218
rect 19432 11154 19484 11160
rect 19628 11098 19656 11630
rect 19260 11070 19656 11098
rect 19260 11014 19288 11070
rect 19248 11008 19300 11014
rect 19248 10950 19300 10956
rect 19156 10600 19208 10606
rect 19156 10542 19208 10548
rect 19260 9518 19288 10950
rect 19720 10674 19748 13756
rect 19708 10668 19760 10674
rect 19708 10610 19760 10616
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 19352 9722 19380 10134
rect 19720 9994 19748 10610
rect 19708 9988 19760 9994
rect 19708 9930 19760 9936
rect 19340 9716 19392 9722
rect 19340 9658 19392 9664
rect 19614 9616 19670 9625
rect 19614 9551 19670 9560
rect 19248 9512 19300 9518
rect 19248 9454 19300 9460
rect 19156 8968 19208 8974
rect 19260 8956 19288 9454
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19208 8928 19288 8956
rect 19156 8910 19208 8916
rect 19260 8498 19288 8928
rect 19352 8906 19380 9318
rect 19628 9042 19656 9551
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19352 8634 19380 8842
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19260 8022 19288 8434
rect 19248 8016 19300 8022
rect 19248 7958 19300 7964
rect 19156 7948 19208 7954
rect 19076 7908 19156 7936
rect 19156 7890 19208 7896
rect 19064 6792 19116 6798
rect 19064 6734 19116 6740
rect 18972 6248 19024 6254
rect 18972 6190 19024 6196
rect 18788 6112 18840 6118
rect 18788 6054 18840 6060
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18604 4616 18656 4622
rect 18604 4558 18656 4564
rect 18616 4282 18644 4558
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18708 4146 18736 5510
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 16764 2984 16816 2990
rect 16764 2926 16816 2932
rect 17420 800 17448 2994
rect 18708 800 18736 2994
rect 18800 2990 18828 6054
rect 18984 5166 19012 6190
rect 19076 5710 19104 6734
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 19168 5234 19196 7890
rect 19352 7750 19380 8570
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19352 7002 19380 7686
rect 19444 7206 19472 8230
rect 19432 7200 19484 7206
rect 19432 7142 19484 7148
rect 19340 6996 19392 7002
rect 19340 6938 19392 6944
rect 19340 6656 19392 6662
rect 19340 6598 19392 6604
rect 19352 6361 19380 6598
rect 19338 6352 19394 6361
rect 19444 6322 19472 7142
rect 19338 6287 19394 6296
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19352 5370 19380 5646
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19536 5234 19564 8910
rect 19628 8634 19656 8978
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19812 8430 19840 15982
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19904 15434 19932 15846
rect 19996 15722 20024 19790
rect 20088 19417 20116 19790
rect 20074 19408 20130 19417
rect 20074 19343 20130 19352
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20088 15858 20116 17614
rect 20180 16017 20208 22066
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20272 20466 20300 20742
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20548 20369 20576 22510
rect 20996 22432 21048 22438
rect 20996 22374 21048 22380
rect 21008 22166 21036 22374
rect 20996 22160 21048 22166
rect 20996 22102 21048 22108
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20640 21010 20668 21286
rect 20720 21072 20772 21078
rect 20720 21014 20772 21020
rect 20628 21004 20680 21010
rect 20628 20946 20680 20952
rect 20534 20360 20590 20369
rect 20534 20295 20590 20304
rect 20548 19990 20576 20295
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18290 20300 19110
rect 20350 18864 20406 18873
rect 20350 18799 20352 18808
rect 20404 18799 20406 18808
rect 20352 18770 20404 18776
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20548 17746 20576 18022
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20272 17338 20300 17614
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 20548 17241 20576 17682
rect 20534 17232 20590 17241
rect 20534 17167 20590 17176
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20364 16046 20392 16390
rect 20352 16040 20404 16046
rect 20166 16008 20222 16017
rect 20352 15982 20404 15988
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 20166 15943 20222 15952
rect 20088 15830 20392 15858
rect 19996 15694 20300 15722
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 19892 15428 19944 15434
rect 19892 15370 19944 15376
rect 19904 15094 19932 15370
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19892 15088 19944 15094
rect 19892 15030 19944 15036
rect 19996 14958 20024 15302
rect 20074 15192 20130 15201
rect 20074 15127 20130 15136
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19904 14618 19932 14758
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 20088 14550 20116 15127
rect 20076 14544 20128 14550
rect 20076 14486 20128 14492
rect 20180 14396 20208 15438
rect 19996 14368 20208 14396
rect 19996 12866 20024 14368
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20076 13728 20128 13734
rect 20074 13696 20076 13705
rect 20128 13696 20130 13705
rect 20074 13631 20130 13640
rect 20088 12986 20116 13631
rect 20180 12986 20208 14010
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 19996 12838 20208 12866
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19904 12442 19932 12582
rect 19892 12436 19944 12442
rect 19892 12378 19944 12384
rect 19996 12102 20024 12650
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19892 11688 19944 11694
rect 19892 11630 19944 11636
rect 19904 11218 19932 11630
rect 20180 11370 20208 12838
rect 19996 11354 20208 11370
rect 19984 11348 20208 11354
rect 20036 11342 20208 11348
rect 19984 11290 20036 11296
rect 19892 11212 19944 11218
rect 19892 11154 19944 11160
rect 19904 10538 19932 11154
rect 19892 10532 19944 10538
rect 19892 10474 19944 10480
rect 19800 8424 19852 8430
rect 19800 8366 19852 8372
rect 19996 8090 20024 11290
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20088 10266 20116 11086
rect 20076 10260 20128 10266
rect 20076 10202 20128 10208
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19708 7812 19760 7818
rect 19708 7754 19760 7760
rect 19720 7546 19748 7754
rect 19708 7540 19760 7546
rect 19708 7482 19760 7488
rect 20272 7342 20300 15694
rect 20364 14618 20392 15830
rect 20456 15162 20484 15982
rect 20548 15706 20576 17167
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20640 15502 20668 20946
rect 20732 20602 20760 21014
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20720 20596 20772 20602
rect 20720 20538 20772 20544
rect 20916 20058 20944 20878
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 21008 19854 21036 21422
rect 21100 20398 21128 22510
rect 21192 22234 21220 22510
rect 21180 22228 21232 22234
rect 21180 22170 21232 22176
rect 21376 22094 21404 26862
rect 21640 26852 21692 26858
rect 21640 26794 21692 26800
rect 21652 26518 21680 26794
rect 21916 26784 21968 26790
rect 21916 26726 21968 26732
rect 21640 26512 21692 26518
rect 21640 26454 21692 26460
rect 21548 26240 21600 26246
rect 21548 26182 21600 26188
rect 21560 25906 21588 26182
rect 21548 25900 21600 25906
rect 21548 25842 21600 25848
rect 21456 25764 21508 25770
rect 21456 25706 21508 25712
rect 21468 25498 21496 25706
rect 21456 25492 21508 25498
rect 21456 25434 21508 25440
rect 21456 24812 21508 24818
rect 21456 24754 21508 24760
rect 21192 22066 21404 22094
rect 21192 20806 21220 22066
rect 21364 21684 21416 21690
rect 21364 21626 21416 21632
rect 21272 21412 21324 21418
rect 21272 21354 21324 21360
rect 21284 21146 21312 21354
rect 21272 21140 21324 21146
rect 21272 21082 21324 21088
rect 21376 21010 21404 21626
rect 21272 21004 21324 21010
rect 21272 20946 21324 20952
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 21284 20806 21312 20946
rect 21180 20800 21232 20806
rect 21180 20742 21232 20748
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21088 20392 21140 20398
rect 21088 20334 21140 20340
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 21100 19310 21128 20334
rect 21192 19514 21220 20742
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21284 20058 21312 20334
rect 21272 20052 21324 20058
rect 21272 19994 21324 20000
rect 21376 19938 21404 20946
rect 21468 20466 21496 24754
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21456 20460 21508 20466
rect 21456 20402 21508 20408
rect 21284 19910 21404 19938
rect 21180 19508 21232 19514
rect 21180 19450 21232 19456
rect 21284 19334 21312 19910
rect 21560 19904 21588 20538
rect 21468 19876 21588 19904
rect 21364 19848 21416 19854
rect 21468 19836 21496 19876
rect 21416 19808 21496 19836
rect 21364 19790 21416 19796
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21192 19306 21312 19334
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18970 20760 19110
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20824 17814 20852 18226
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20824 16726 20852 17750
rect 20812 16720 20864 16726
rect 20812 16662 20864 16668
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 20732 15706 20760 16390
rect 20812 16176 20864 16182
rect 20812 16118 20864 16124
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20444 15156 20496 15162
rect 20444 15098 20496 15104
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20364 14074 20392 14554
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20352 13864 20404 13870
rect 20352 13806 20404 13812
rect 20364 12434 20392 13806
rect 20456 13734 20484 15098
rect 20536 14884 20588 14890
rect 20536 14826 20588 14832
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20548 14482 20576 14826
rect 20628 14816 20680 14822
rect 20628 14758 20680 14764
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20548 14278 20576 14418
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20536 14068 20588 14074
rect 20536 14010 20588 14016
rect 20444 13728 20496 13734
rect 20444 13670 20496 13676
rect 20456 12714 20484 13670
rect 20444 12708 20496 12714
rect 20444 12650 20496 12656
rect 20364 12406 20484 12434
rect 20456 10606 20484 12406
rect 20548 11558 20576 14010
rect 20640 13394 20668 14758
rect 20732 13530 20760 14826
rect 20824 13802 20852 16118
rect 20916 16046 20944 17818
rect 21008 17542 21036 18702
rect 20996 17536 21048 17542
rect 20996 17478 21048 17484
rect 20904 16040 20956 16046
rect 21192 15994 21220 19306
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 21284 17542 21312 17682
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21284 17134 21312 17478
rect 21376 17134 21404 18566
rect 21272 17128 21324 17134
rect 21272 17070 21324 17076
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 21468 16946 21496 19450
rect 21652 19334 21680 26454
rect 21732 24880 21784 24886
rect 21732 24822 21784 24828
rect 21744 24070 21772 24822
rect 21928 24290 21956 26726
rect 22112 25378 22140 34002
rect 22836 33856 22888 33862
rect 22836 33798 22888 33804
rect 22328 33756 22636 33765
rect 22328 33754 22334 33756
rect 22390 33754 22414 33756
rect 22470 33754 22494 33756
rect 22550 33754 22574 33756
rect 22630 33754 22636 33756
rect 22390 33702 22392 33754
rect 22572 33702 22574 33754
rect 22328 33700 22334 33702
rect 22390 33700 22414 33702
rect 22470 33700 22494 33702
rect 22550 33700 22574 33702
rect 22630 33700 22636 33702
rect 22328 33691 22636 33700
rect 22328 32668 22636 32677
rect 22328 32666 22334 32668
rect 22390 32666 22414 32668
rect 22470 32666 22494 32668
rect 22550 32666 22574 32668
rect 22630 32666 22636 32668
rect 22390 32614 22392 32666
rect 22572 32614 22574 32666
rect 22328 32612 22334 32614
rect 22390 32612 22414 32614
rect 22470 32612 22494 32614
rect 22550 32612 22574 32614
rect 22630 32612 22636 32614
rect 22328 32603 22636 32612
rect 22848 31754 22876 33798
rect 22988 33212 23296 33221
rect 22988 33210 22994 33212
rect 23050 33210 23074 33212
rect 23130 33210 23154 33212
rect 23210 33210 23234 33212
rect 23290 33210 23296 33212
rect 23050 33158 23052 33210
rect 23232 33158 23234 33210
rect 22988 33156 22994 33158
rect 23050 33156 23074 33158
rect 23130 33156 23154 33158
rect 23210 33156 23234 33158
rect 23290 33156 23296 33158
rect 22988 33147 23296 33156
rect 23848 32224 23900 32230
rect 23848 32166 23900 32172
rect 24032 32224 24084 32230
rect 24032 32166 24084 32172
rect 22988 32124 23296 32133
rect 22988 32122 22994 32124
rect 23050 32122 23074 32124
rect 23130 32122 23154 32124
rect 23210 32122 23234 32124
rect 23290 32122 23296 32124
rect 23050 32070 23052 32122
rect 23232 32070 23234 32122
rect 22988 32068 22994 32070
rect 23050 32068 23074 32070
rect 23130 32068 23154 32070
rect 23210 32068 23234 32070
rect 23290 32068 23296 32070
rect 22988 32059 23296 32068
rect 22756 31726 22876 31754
rect 22328 31580 22636 31589
rect 22328 31578 22334 31580
rect 22390 31578 22414 31580
rect 22470 31578 22494 31580
rect 22550 31578 22574 31580
rect 22630 31578 22636 31580
rect 22390 31526 22392 31578
rect 22572 31526 22574 31578
rect 22328 31524 22334 31526
rect 22390 31524 22414 31526
rect 22470 31524 22494 31526
rect 22550 31524 22574 31526
rect 22630 31524 22636 31526
rect 22328 31515 22636 31524
rect 22560 31204 22612 31210
rect 22560 31146 22612 31152
rect 22572 30938 22600 31146
rect 22560 30932 22612 30938
rect 22560 30874 22612 30880
rect 22328 30492 22636 30501
rect 22328 30490 22334 30492
rect 22390 30490 22414 30492
rect 22470 30490 22494 30492
rect 22550 30490 22574 30492
rect 22630 30490 22636 30492
rect 22390 30438 22392 30490
rect 22572 30438 22574 30490
rect 22328 30436 22334 30438
rect 22390 30436 22414 30438
rect 22470 30436 22494 30438
rect 22550 30436 22574 30438
rect 22630 30436 22636 30438
rect 22328 30427 22636 30436
rect 22328 29404 22636 29413
rect 22328 29402 22334 29404
rect 22390 29402 22414 29404
rect 22470 29402 22494 29404
rect 22550 29402 22574 29404
rect 22630 29402 22636 29404
rect 22390 29350 22392 29402
rect 22572 29350 22574 29402
rect 22328 29348 22334 29350
rect 22390 29348 22414 29350
rect 22470 29348 22494 29350
rect 22550 29348 22574 29350
rect 22630 29348 22636 29350
rect 22328 29339 22636 29348
rect 22560 29300 22612 29306
rect 22560 29242 22612 29248
rect 22572 28694 22600 29242
rect 22560 28688 22612 28694
rect 22560 28630 22612 28636
rect 22652 28620 22704 28626
rect 22652 28562 22704 28568
rect 22328 28316 22636 28325
rect 22328 28314 22334 28316
rect 22390 28314 22414 28316
rect 22470 28314 22494 28316
rect 22550 28314 22574 28316
rect 22630 28314 22636 28316
rect 22390 28262 22392 28314
rect 22572 28262 22574 28314
rect 22328 28260 22334 28262
rect 22390 28260 22414 28262
rect 22470 28260 22494 28262
rect 22550 28260 22574 28262
rect 22630 28260 22636 28262
rect 22328 28251 22636 28260
rect 22664 27962 22692 28562
rect 22572 27934 22692 27962
rect 22572 27878 22600 27934
rect 22192 27872 22244 27878
rect 22192 27814 22244 27820
rect 22560 27872 22612 27878
rect 22560 27814 22612 27820
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22204 26790 22232 27814
rect 22328 27228 22636 27237
rect 22328 27226 22334 27228
rect 22390 27226 22414 27228
rect 22470 27226 22494 27228
rect 22550 27226 22574 27228
rect 22630 27226 22636 27228
rect 22390 27174 22392 27226
rect 22572 27174 22574 27226
rect 22328 27172 22334 27174
rect 22390 27172 22414 27174
rect 22470 27172 22494 27174
rect 22550 27172 22574 27174
rect 22630 27172 22636 27174
rect 22328 27163 22636 27172
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22192 26444 22244 26450
rect 22192 26386 22244 26392
rect 22204 25430 22232 26386
rect 22328 26140 22636 26149
rect 22328 26138 22334 26140
rect 22390 26138 22414 26140
rect 22470 26138 22494 26140
rect 22550 26138 22574 26140
rect 22630 26138 22636 26140
rect 22390 26086 22392 26138
rect 22572 26086 22574 26138
rect 22328 26084 22334 26086
rect 22390 26084 22414 26086
rect 22470 26084 22494 26086
rect 22550 26084 22574 26086
rect 22630 26084 22636 26086
rect 22328 26075 22636 26084
rect 22560 25764 22612 25770
rect 22560 25706 22612 25712
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22388 25498 22416 25638
rect 22572 25498 22600 25706
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22020 25350 22140 25378
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 22020 24410 22048 25350
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22112 24818 22140 25230
rect 22328 25052 22636 25061
rect 22328 25050 22334 25052
rect 22390 25050 22414 25052
rect 22470 25050 22494 25052
rect 22550 25050 22574 25052
rect 22630 25050 22636 25052
rect 22390 24998 22392 25050
rect 22572 24998 22574 25050
rect 22328 24996 22334 24998
rect 22390 24996 22414 24998
rect 22470 24996 22494 24998
rect 22550 24996 22574 24998
rect 22630 24996 22636 24998
rect 22328 24987 22636 24996
rect 22664 24868 22692 27814
rect 22572 24840 22692 24868
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22572 24614 22600 24840
rect 22560 24608 22612 24614
rect 22560 24550 22612 24556
rect 22008 24404 22060 24410
rect 22008 24346 22060 24352
rect 22100 24404 22152 24410
rect 22100 24346 22152 24352
rect 21928 24262 22048 24290
rect 21732 24064 21784 24070
rect 21732 24006 21784 24012
rect 21744 23662 21772 24006
rect 21732 23656 21784 23662
rect 21732 23598 21784 23604
rect 21744 22030 21772 23598
rect 21824 23180 21876 23186
rect 21824 23122 21876 23128
rect 21836 22506 21864 23122
rect 21824 22500 21876 22506
rect 21824 22442 21876 22448
rect 21916 22432 21968 22438
rect 21916 22374 21968 22380
rect 21928 22234 21956 22374
rect 21916 22228 21968 22234
rect 21916 22170 21968 22176
rect 22020 22114 22048 24262
rect 22112 23610 22140 24346
rect 22572 24342 22600 24550
rect 22560 24336 22612 24342
rect 22560 24278 22612 24284
rect 22652 24200 22704 24206
rect 22652 24142 22704 24148
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22204 23730 22232 24006
rect 22328 23964 22636 23973
rect 22328 23962 22334 23964
rect 22390 23962 22414 23964
rect 22470 23962 22494 23964
rect 22550 23962 22574 23964
rect 22630 23962 22636 23964
rect 22390 23910 22392 23962
rect 22572 23910 22574 23962
rect 22328 23908 22334 23910
rect 22390 23908 22414 23910
rect 22470 23908 22494 23910
rect 22550 23908 22574 23910
rect 22630 23908 22636 23910
rect 22328 23899 22636 23908
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22112 23582 22232 23610
rect 21928 22086 22048 22114
rect 22204 22094 22232 23582
rect 22664 23322 22692 24142
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22328 22876 22636 22885
rect 22328 22874 22334 22876
rect 22390 22874 22414 22876
rect 22470 22874 22494 22876
rect 22550 22874 22574 22876
rect 22630 22874 22636 22876
rect 22390 22822 22392 22874
rect 22572 22822 22574 22874
rect 22328 22820 22334 22822
rect 22390 22820 22414 22822
rect 22470 22820 22494 22822
rect 22550 22820 22574 22822
rect 22630 22820 22636 22822
rect 22328 22811 22636 22820
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22664 22234 22692 22510
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 22756 22094 22784 31726
rect 23296 31680 23348 31686
rect 23296 31622 23348 31628
rect 23308 31346 23336 31622
rect 23296 31340 23348 31346
rect 23296 31282 23348 31288
rect 23308 31124 23336 31282
rect 23664 31272 23716 31278
rect 23664 31214 23716 31220
rect 23308 31096 23428 31124
rect 22988 31036 23296 31045
rect 22988 31034 22994 31036
rect 23050 31034 23074 31036
rect 23130 31034 23154 31036
rect 23210 31034 23234 31036
rect 23290 31034 23296 31036
rect 23050 30982 23052 31034
rect 23232 30982 23234 31034
rect 22988 30980 22994 30982
rect 23050 30980 23074 30982
rect 23130 30980 23154 30982
rect 23210 30980 23234 30982
rect 23290 30980 23296 30982
rect 22988 30971 23296 30980
rect 23400 30258 23428 31096
rect 23480 30592 23532 30598
rect 23480 30534 23532 30540
rect 23492 30326 23520 30534
rect 23676 30326 23704 31214
rect 23480 30320 23532 30326
rect 23480 30262 23532 30268
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 23388 30252 23440 30258
rect 23388 30194 23440 30200
rect 23388 30048 23440 30054
rect 23388 29990 23440 29996
rect 23572 30048 23624 30054
rect 23572 29990 23624 29996
rect 22988 29948 23296 29957
rect 22988 29946 22994 29948
rect 23050 29946 23074 29948
rect 23130 29946 23154 29948
rect 23210 29946 23234 29948
rect 23290 29946 23296 29948
rect 23050 29894 23052 29946
rect 23232 29894 23234 29946
rect 22988 29892 22994 29894
rect 23050 29892 23074 29894
rect 23130 29892 23154 29894
rect 23210 29892 23234 29894
rect 23290 29892 23296 29894
rect 22988 29883 23296 29892
rect 23400 29306 23428 29990
rect 23584 29578 23612 29990
rect 23572 29572 23624 29578
rect 23572 29514 23624 29520
rect 23480 29504 23532 29510
rect 23480 29446 23532 29452
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23492 29102 23520 29446
rect 23480 29096 23532 29102
rect 23480 29038 23532 29044
rect 22836 29028 22888 29034
rect 22836 28970 22888 28976
rect 23388 29028 23440 29034
rect 23388 28970 23440 28976
rect 22848 28762 22876 28970
rect 22988 28860 23296 28869
rect 22988 28858 22994 28860
rect 23050 28858 23074 28860
rect 23130 28858 23154 28860
rect 23210 28858 23234 28860
rect 23290 28858 23296 28860
rect 23050 28806 23052 28858
rect 23232 28806 23234 28858
rect 22988 28804 22994 28806
rect 23050 28804 23074 28806
rect 23130 28804 23154 28806
rect 23210 28804 23234 28806
rect 23290 28804 23296 28806
rect 22988 28795 23296 28804
rect 23400 28762 23428 28970
rect 22836 28756 22888 28762
rect 22836 28698 22888 28704
rect 23388 28756 23440 28762
rect 23388 28698 23440 28704
rect 22836 28620 22888 28626
rect 22836 28562 22888 28568
rect 22848 28150 22876 28562
rect 23400 28218 23428 28698
rect 23492 28694 23520 29038
rect 23480 28688 23532 28694
rect 23480 28630 23532 28636
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 22836 28144 22888 28150
rect 22836 28086 22888 28092
rect 22988 27772 23296 27781
rect 22988 27770 22994 27772
rect 23050 27770 23074 27772
rect 23130 27770 23154 27772
rect 23210 27770 23234 27772
rect 23290 27770 23296 27772
rect 23050 27718 23052 27770
rect 23232 27718 23234 27770
rect 22988 27716 22994 27718
rect 23050 27716 23074 27718
rect 23130 27716 23154 27718
rect 23210 27716 23234 27718
rect 23290 27716 23296 27718
rect 22988 27707 23296 27716
rect 23400 27606 23428 28154
rect 23388 27600 23440 27606
rect 23388 27542 23440 27548
rect 23584 27452 23612 29514
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23768 27606 23796 29038
rect 23756 27600 23808 27606
rect 23756 27542 23808 27548
rect 23400 27424 23612 27452
rect 23296 27328 23348 27334
rect 23296 27270 23348 27276
rect 23308 26858 23336 27270
rect 23296 26852 23348 26858
rect 23296 26794 23348 26800
rect 22988 26684 23296 26693
rect 22988 26682 22994 26684
rect 23050 26682 23074 26684
rect 23130 26682 23154 26684
rect 23210 26682 23234 26684
rect 23290 26682 23296 26684
rect 23050 26630 23052 26682
rect 23232 26630 23234 26682
rect 22988 26628 22994 26630
rect 23050 26628 23074 26630
rect 23130 26628 23154 26630
rect 23210 26628 23234 26630
rect 23290 26628 23296 26630
rect 22988 26619 23296 26628
rect 23400 26568 23428 27424
rect 23308 26540 23428 26568
rect 23308 26042 23336 26540
rect 23860 26518 23888 32166
rect 24044 31958 24072 32166
rect 24032 31952 24084 31958
rect 24032 31894 24084 31900
rect 24136 31142 24164 34002
rect 25148 33998 25176 35678
rect 26056 34060 26108 34066
rect 26056 34002 26108 34008
rect 25136 33992 25188 33998
rect 25136 33934 25188 33940
rect 24492 32428 24544 32434
rect 24492 32370 24544 32376
rect 24124 31136 24176 31142
rect 24124 31078 24176 31084
rect 24032 30728 24084 30734
rect 24032 30670 24084 30676
rect 24044 30394 24072 30670
rect 24032 30388 24084 30394
rect 24032 30330 24084 30336
rect 24032 30252 24084 30258
rect 24032 30194 24084 30200
rect 24044 28422 24072 30194
rect 24504 29628 24532 32370
rect 24860 32224 24912 32230
rect 24860 32166 24912 32172
rect 25228 32224 25280 32230
rect 25228 32166 25280 32172
rect 24872 31890 24900 32166
rect 25240 32026 25268 32166
rect 26068 32026 26096 34002
rect 26436 33522 26464 35678
rect 28368 34134 28396 35678
rect 28356 34128 28408 34134
rect 28356 34070 28408 34076
rect 29656 33998 29684 35678
rect 30944 35578 30972 35678
rect 31036 35578 31064 35686
rect 30944 35550 31064 35578
rect 30877 34300 31185 34309
rect 30877 34298 30883 34300
rect 30939 34298 30963 34300
rect 31019 34298 31043 34300
rect 31099 34298 31123 34300
rect 31179 34298 31185 34300
rect 30939 34246 30941 34298
rect 31121 34246 31123 34298
rect 30877 34244 30883 34246
rect 30939 34244 30963 34246
rect 31019 34244 31043 34246
rect 31099 34244 31123 34246
rect 31179 34244 31185 34246
rect 30877 34235 31185 34244
rect 30012 34060 30064 34066
rect 30012 34002 30064 34008
rect 31208 34060 31260 34066
rect 31208 34002 31260 34008
rect 29644 33992 29696 33998
rect 29644 33934 29696 33940
rect 26424 33516 26476 33522
rect 26424 33458 26476 33464
rect 26516 33448 26568 33454
rect 26516 33390 26568 33396
rect 25228 32020 25280 32026
rect 25228 31962 25280 31968
rect 26056 32020 26108 32026
rect 26056 31962 26108 31968
rect 24860 31884 24912 31890
rect 24860 31826 24912 31832
rect 26528 31770 26556 33390
rect 29276 32972 29328 32978
rect 29276 32914 29328 32920
rect 26792 32564 26844 32570
rect 26792 32506 26844 32512
rect 26436 31742 26556 31770
rect 24768 31136 24820 31142
rect 24768 31078 24820 31084
rect 24780 30802 24808 31078
rect 24768 30796 24820 30802
rect 24768 30738 24820 30744
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 24952 30592 25004 30598
rect 24952 30534 25004 30540
rect 24964 30258 24992 30534
rect 24952 30252 25004 30258
rect 24952 30194 25004 30200
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 25056 30054 25084 30194
rect 25044 30048 25096 30054
rect 25044 29990 25096 29996
rect 25228 30048 25280 30054
rect 25228 29990 25280 29996
rect 24768 29640 24820 29646
rect 24504 29600 24768 29628
rect 24768 29582 24820 29588
rect 24780 29510 24808 29582
rect 24768 29504 24820 29510
rect 24768 29446 24820 29452
rect 24952 29504 25004 29510
rect 24952 29446 25004 29452
rect 24676 28960 24728 28966
rect 24676 28902 24728 28908
rect 24688 28694 24716 28902
rect 24676 28688 24728 28694
rect 24676 28630 24728 28636
rect 24768 28552 24820 28558
rect 24768 28494 24820 28500
rect 24032 28416 24084 28422
rect 24032 28358 24084 28364
rect 24044 28218 24072 28358
rect 24032 28212 24084 28218
rect 24032 28154 24084 28160
rect 24044 26994 24072 28154
rect 24216 28008 24268 28014
rect 24216 27950 24268 27956
rect 24228 27538 24256 27950
rect 24676 27600 24728 27606
rect 24676 27542 24728 27548
rect 24216 27532 24268 27538
rect 24216 27474 24268 27480
rect 24308 27464 24360 27470
rect 24308 27406 24360 27412
rect 24124 27328 24176 27334
rect 24124 27270 24176 27276
rect 24136 27130 24164 27270
rect 24124 27124 24176 27130
rect 24124 27066 24176 27072
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 23848 26512 23900 26518
rect 23900 26472 23980 26500
rect 23848 26454 23900 26460
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 22836 26036 22888 26042
rect 22836 25978 22888 25984
rect 23296 26036 23348 26042
rect 23296 25978 23348 25984
rect 22848 24818 22876 25978
rect 22988 25596 23296 25605
rect 22988 25594 22994 25596
rect 23050 25594 23074 25596
rect 23130 25594 23154 25596
rect 23210 25594 23234 25596
rect 23290 25594 23296 25596
rect 23050 25542 23052 25594
rect 23232 25542 23234 25594
rect 22988 25540 22994 25542
rect 23050 25540 23074 25542
rect 23130 25540 23154 25542
rect 23210 25540 23234 25542
rect 23290 25540 23296 25542
rect 22988 25531 23296 25540
rect 23112 25492 23164 25498
rect 23112 25434 23164 25440
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 22836 24812 22888 24818
rect 22836 24754 22888 24760
rect 22940 24682 22968 25298
rect 23124 24750 23152 25434
rect 23400 25430 23428 26386
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23388 25424 23440 25430
rect 23388 25366 23440 25372
rect 23492 25378 23520 26318
rect 23492 25350 23612 25378
rect 23480 25288 23532 25294
rect 23480 25230 23532 25236
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 23308 24818 23336 25094
rect 23492 24954 23520 25230
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23296 24812 23348 24818
rect 23296 24754 23348 24760
rect 23112 24744 23164 24750
rect 23112 24686 23164 24692
rect 22928 24676 22980 24682
rect 22928 24618 22980 24624
rect 22988 24508 23296 24517
rect 22988 24506 22994 24508
rect 23050 24506 23074 24508
rect 23130 24506 23154 24508
rect 23210 24506 23234 24508
rect 23290 24506 23296 24508
rect 23050 24454 23052 24506
rect 23232 24454 23234 24506
rect 22988 24452 22994 24454
rect 23050 24452 23074 24454
rect 23130 24452 23154 24454
rect 23210 24452 23234 24454
rect 23290 24452 23296 24454
rect 22988 24443 23296 24452
rect 23388 24336 23440 24342
rect 23584 24290 23612 25350
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23768 24954 23796 25230
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 23756 24608 23808 24614
rect 23756 24550 23808 24556
rect 23388 24278 23440 24284
rect 22988 23420 23296 23429
rect 22988 23418 22994 23420
rect 23050 23418 23074 23420
rect 23130 23418 23154 23420
rect 23210 23418 23234 23420
rect 23290 23418 23296 23420
rect 23050 23366 23052 23418
rect 23232 23366 23234 23418
rect 22988 23364 22994 23366
rect 23050 23364 23074 23366
rect 23130 23364 23154 23366
rect 23210 23364 23234 23366
rect 23290 23364 23296 23366
rect 22988 23355 23296 23364
rect 22836 22432 22888 22438
rect 22836 22374 22888 22380
rect 22848 22216 22876 22374
rect 22988 22332 23296 22341
rect 22988 22330 22994 22332
rect 23050 22330 23074 22332
rect 23130 22330 23154 22332
rect 23210 22330 23234 22332
rect 23290 22330 23296 22332
rect 23050 22278 23052 22330
rect 23232 22278 23234 22330
rect 22988 22276 22994 22278
rect 23050 22276 23074 22278
rect 23130 22276 23154 22278
rect 23210 22276 23234 22278
rect 23290 22276 23296 22278
rect 22988 22267 23296 22276
rect 22848 22188 22968 22216
rect 22940 22098 22968 22188
rect 23296 22160 23348 22166
rect 23202 22128 23258 22137
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21928 21894 21956 22086
rect 22204 22066 22600 22094
rect 22756 22066 22876 22094
rect 22572 21894 22600 22066
rect 22744 22024 22796 22030
rect 22664 21984 22744 22012
rect 21916 21888 21968 21894
rect 21916 21830 21968 21836
rect 22008 21888 22060 21894
rect 22008 21830 22060 21836
rect 22192 21888 22244 21894
rect 22192 21830 22244 21836
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 21928 21298 21956 21830
rect 22020 21418 22048 21830
rect 22008 21412 22060 21418
rect 22008 21354 22060 21360
rect 21928 21270 22048 21298
rect 21916 20936 21968 20942
rect 21916 20878 21968 20884
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21836 20398 21864 20538
rect 21928 20398 21956 20878
rect 21824 20392 21876 20398
rect 21916 20392 21968 20398
rect 21824 20334 21876 20340
rect 21914 20360 21916 20369
rect 21968 20360 21970 20369
rect 21652 19306 21772 19334
rect 21640 18624 21692 18630
rect 21640 18566 21692 18572
rect 21548 18148 21600 18154
rect 21548 18090 21600 18096
rect 21560 17338 21588 18090
rect 21652 17746 21680 18566
rect 21640 17740 21692 17746
rect 21640 17682 21692 17688
rect 21548 17332 21600 17338
rect 21548 17274 21600 17280
rect 20904 15982 20956 15988
rect 21100 15966 21220 15994
rect 21376 16918 21496 16946
rect 20902 15872 20958 15881
rect 20958 15830 21036 15858
rect 20902 15807 20958 15816
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20916 14958 20944 15438
rect 20904 14952 20956 14958
rect 20904 14894 20956 14900
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 20824 13530 20852 13738
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20732 11898 20760 12378
rect 20916 12306 20944 13330
rect 21008 12442 21036 15830
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20996 12300 21048 12306
rect 20996 12242 21048 12248
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 20720 11892 20772 11898
rect 20720 11834 20772 11840
rect 20824 11558 20852 12174
rect 20916 11694 20944 12242
rect 20904 11688 20956 11694
rect 20904 11630 20956 11636
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20444 10600 20496 10606
rect 20444 10542 20496 10548
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20364 9178 20392 9454
rect 20456 9382 20484 10542
rect 20548 9586 20576 11494
rect 21008 11354 21036 12242
rect 21100 12238 21128 15966
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21192 14550 21220 15846
rect 21180 14544 21232 14550
rect 21180 14486 21232 14492
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21192 13530 21220 14350
rect 21284 13870 21312 14350
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 21180 13524 21232 13530
rect 21180 13466 21232 13472
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 21008 10606 21036 10950
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20640 10266 20668 10406
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20260 7336 20312 7342
rect 20260 7278 20312 7284
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19628 6458 19656 6598
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19616 6112 19668 6118
rect 19616 6054 19668 6060
rect 19628 5234 19656 6054
rect 19812 5370 19840 6258
rect 19904 6254 19932 7142
rect 20272 6322 20300 7278
rect 20352 7268 20404 7274
rect 20456 7256 20484 9318
rect 20548 8430 20576 9522
rect 20732 9178 20760 9998
rect 20812 9648 20864 9654
rect 20812 9590 20864 9596
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20824 8566 20852 9590
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20916 9042 20944 9318
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 21100 8786 21128 12174
rect 21272 12164 21324 12170
rect 21272 12106 21324 12112
rect 21284 11801 21312 12106
rect 21270 11792 21326 11801
rect 21270 11727 21326 11736
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21284 10538 21312 10950
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 21192 9926 21220 10406
rect 21180 9920 21232 9926
rect 21180 9862 21232 9868
rect 21192 8974 21220 9862
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21008 8758 21128 8786
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 21008 8294 21036 8758
rect 21088 8424 21140 8430
rect 21088 8366 21140 8372
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20404 7228 20484 7256
rect 20352 7210 20404 7216
rect 20364 7002 20392 7210
rect 20720 7200 20772 7206
rect 20720 7142 20772 7148
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 19892 6248 19944 6254
rect 19892 6190 19944 6196
rect 20272 5914 20300 6258
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 19800 5364 19852 5370
rect 19800 5306 19852 5312
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19524 5228 19576 5234
rect 19524 5170 19576 5176
rect 19616 5228 19668 5234
rect 19616 5170 19668 5176
rect 20364 5166 20392 6938
rect 20732 6934 20760 7142
rect 20720 6928 20772 6934
rect 20720 6870 20772 6876
rect 21008 6866 21036 7142
rect 20996 6860 21048 6866
rect 20996 6802 21048 6808
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20824 5234 20852 5510
rect 20812 5228 20864 5234
rect 20812 5170 20864 5176
rect 18972 5160 19024 5166
rect 18972 5102 19024 5108
rect 20352 5160 20404 5166
rect 20352 5102 20404 5108
rect 20076 5092 20128 5098
rect 20076 5034 20128 5040
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19168 4758 19196 4966
rect 20088 4826 20116 5034
rect 20076 4820 20128 4826
rect 20076 4762 20128 4768
rect 19156 4752 19208 4758
rect 19156 4694 19208 4700
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19352 3602 19380 4422
rect 20088 4146 20116 4762
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19340 3596 19392 3602
rect 19340 3538 19392 3544
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 18788 2984 18840 2990
rect 18788 2926 18840 2932
rect 20640 800 20668 3470
rect 21100 2922 21128 8366
rect 21192 7750 21220 8910
rect 21180 7744 21232 7750
rect 21180 7686 21232 7692
rect 21192 6662 21220 7686
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 21284 7342 21312 7414
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21376 7256 21404 16918
rect 21652 16794 21680 17682
rect 21640 16788 21692 16794
rect 21640 16730 21692 16736
rect 21652 15910 21680 16730
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21640 15904 21692 15910
rect 21640 15846 21692 15852
rect 21468 12714 21496 15846
rect 21640 15088 21692 15094
rect 21640 15030 21692 15036
rect 21548 14816 21600 14822
rect 21548 14758 21600 14764
rect 21560 14074 21588 14758
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21652 13870 21680 15030
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21744 13190 21772 19306
rect 21836 15858 21864 20334
rect 21914 20295 21970 20304
rect 22020 19334 22048 21270
rect 22204 20058 22232 21830
rect 22328 21788 22636 21797
rect 22328 21786 22334 21788
rect 22390 21786 22414 21788
rect 22470 21786 22494 21788
rect 22550 21786 22574 21788
rect 22630 21786 22636 21788
rect 22390 21734 22392 21786
rect 22572 21734 22574 21786
rect 22328 21732 22334 21734
rect 22390 21732 22414 21734
rect 22470 21732 22494 21734
rect 22550 21732 22574 21734
rect 22630 21732 22636 21734
rect 22328 21723 22636 21732
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 22376 21072 22428 21078
rect 22376 21014 22428 21020
rect 22388 20806 22416 21014
rect 22572 20890 22600 21558
rect 22664 21350 22692 21984
rect 22744 21966 22796 21972
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22652 21344 22704 21350
rect 22652 21286 22704 21292
rect 22664 21010 22692 21286
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22572 20862 22692 20890
rect 22664 20806 22692 20862
rect 22376 20800 22428 20806
rect 22376 20742 22428 20748
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22328 20700 22636 20709
rect 22328 20698 22334 20700
rect 22390 20698 22414 20700
rect 22470 20698 22494 20700
rect 22550 20698 22574 20700
rect 22630 20698 22636 20700
rect 22390 20646 22392 20698
rect 22572 20646 22574 20698
rect 22328 20644 22334 20646
rect 22390 20644 22414 20646
rect 22470 20644 22494 20646
rect 22550 20644 22574 20646
rect 22630 20644 22636 20646
rect 22328 20635 22636 20644
rect 22560 20460 22612 20466
rect 22560 20402 22612 20408
rect 22192 20052 22244 20058
rect 22192 19994 22244 20000
rect 22100 19984 22152 19990
rect 22100 19926 22152 19932
rect 22112 19514 22140 19926
rect 22572 19786 22600 20402
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22328 19612 22636 19621
rect 22328 19610 22334 19612
rect 22390 19610 22414 19612
rect 22470 19610 22494 19612
rect 22550 19610 22574 19612
rect 22630 19610 22636 19612
rect 22390 19558 22392 19610
rect 22572 19558 22574 19610
rect 22328 19556 22334 19558
rect 22390 19556 22414 19558
rect 22470 19556 22494 19558
rect 22550 19556 22574 19558
rect 22630 19556 22636 19558
rect 22328 19547 22636 19556
rect 22100 19508 22152 19514
rect 22100 19450 22152 19456
rect 22020 19306 22140 19334
rect 21916 17808 21968 17814
rect 21916 17750 21968 17756
rect 21928 16114 21956 17750
rect 22008 16652 22060 16658
rect 22008 16594 22060 16600
rect 21916 16108 21968 16114
rect 21916 16050 21968 16056
rect 21836 15830 21956 15858
rect 21824 15360 21876 15366
rect 21824 15302 21876 15308
rect 21836 15026 21864 15302
rect 21824 15020 21876 15026
rect 21824 14962 21876 14968
rect 21822 14784 21878 14793
rect 21822 14719 21878 14728
rect 21732 13184 21784 13190
rect 21732 13126 21784 13132
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21456 12708 21508 12714
rect 21456 12650 21508 12656
rect 21468 8022 21496 12650
rect 21548 12096 21600 12102
rect 21548 12038 21600 12044
rect 21456 8016 21508 8022
rect 21456 7958 21508 7964
rect 21560 7750 21588 12038
rect 21652 11694 21680 12854
rect 21640 11688 21692 11694
rect 21640 11630 21692 11636
rect 21836 9994 21864 14719
rect 21928 11898 21956 15830
rect 22020 15706 22048 16594
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22112 15450 22140 19306
rect 22328 18524 22636 18533
rect 22328 18522 22334 18524
rect 22390 18522 22414 18524
rect 22470 18522 22494 18524
rect 22550 18522 22574 18524
rect 22630 18522 22636 18524
rect 22390 18470 22392 18522
rect 22572 18470 22574 18522
rect 22328 18468 22334 18470
rect 22390 18468 22414 18470
rect 22470 18468 22494 18470
rect 22550 18468 22574 18470
rect 22630 18468 22636 18470
rect 22328 18459 22636 18468
rect 22192 18080 22244 18086
rect 22192 18022 22244 18028
rect 22204 17134 22232 18022
rect 22664 17785 22692 20742
rect 22756 17882 22784 21830
rect 22744 17876 22796 17882
rect 22744 17818 22796 17824
rect 22848 17796 22876 22066
rect 22928 22092 22980 22098
rect 23296 22102 23348 22108
rect 23202 22063 23258 22072
rect 22928 22034 22980 22040
rect 22940 21622 22968 22034
rect 23216 22030 23244 22063
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23308 21894 23336 22102
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23400 21690 23428 24278
rect 23492 24262 23612 24290
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 22928 21616 22980 21622
rect 22928 21558 22980 21564
rect 22988 21244 23296 21253
rect 22988 21242 22994 21244
rect 23050 21242 23074 21244
rect 23130 21242 23154 21244
rect 23210 21242 23234 21244
rect 23290 21242 23296 21244
rect 23050 21190 23052 21242
rect 23232 21190 23234 21242
rect 22988 21188 22994 21190
rect 23050 21188 23074 21190
rect 23130 21188 23154 21190
rect 23210 21188 23234 21190
rect 23290 21188 23296 21190
rect 22988 21179 23296 21188
rect 22988 20156 23296 20165
rect 22988 20154 22994 20156
rect 23050 20154 23074 20156
rect 23130 20154 23154 20156
rect 23210 20154 23234 20156
rect 23290 20154 23296 20156
rect 23050 20102 23052 20154
rect 23232 20102 23234 20154
rect 22988 20100 22994 20102
rect 23050 20100 23074 20102
rect 23130 20100 23154 20102
rect 23210 20100 23234 20102
rect 23290 20100 23296 20102
rect 22988 20091 23296 20100
rect 22988 19068 23296 19077
rect 22988 19066 22994 19068
rect 23050 19066 23074 19068
rect 23130 19066 23154 19068
rect 23210 19066 23234 19068
rect 23290 19066 23296 19068
rect 23050 19014 23052 19066
rect 23232 19014 23234 19066
rect 22988 19012 22994 19014
rect 23050 19012 23074 19014
rect 23130 19012 23154 19014
rect 23210 19012 23234 19014
rect 23290 19012 23296 19014
rect 22988 19003 23296 19012
rect 23400 18630 23428 21626
rect 23492 21554 23520 24262
rect 23768 24206 23796 24550
rect 23756 24200 23808 24206
rect 23662 24168 23718 24177
rect 23756 24142 23808 24148
rect 23662 24103 23718 24112
rect 23572 24064 23624 24070
rect 23572 24006 23624 24012
rect 23584 23798 23612 24006
rect 23676 23798 23704 24103
rect 23572 23792 23624 23798
rect 23572 23734 23624 23740
rect 23664 23792 23716 23798
rect 23664 23734 23716 23740
rect 23676 23186 23704 23734
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23480 21548 23532 21554
rect 23480 21490 23532 21496
rect 23584 20602 23612 23054
rect 23768 22574 23796 24142
rect 23756 22568 23808 22574
rect 23756 22510 23808 22516
rect 23848 22432 23900 22438
rect 23848 22374 23900 22380
rect 23860 22166 23888 22374
rect 23848 22160 23900 22166
rect 23848 22102 23900 22108
rect 23952 21570 23980 26472
rect 24044 25906 24072 26930
rect 24320 26246 24348 27406
rect 24688 26926 24716 27542
rect 24780 26926 24808 28494
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 24872 27130 24900 27406
rect 24860 27124 24912 27130
rect 24860 27066 24912 27072
rect 24492 26920 24544 26926
rect 24492 26862 24544 26868
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24768 26920 24820 26926
rect 24768 26862 24820 26868
rect 24308 26240 24360 26246
rect 24308 26182 24360 26188
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 24032 23724 24084 23730
rect 24032 23666 24084 23672
rect 24044 22642 24072 23666
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 24044 21876 24072 22578
rect 24124 21888 24176 21894
rect 24044 21848 24124 21876
rect 24044 21622 24072 21848
rect 24124 21830 24176 21836
rect 23676 21542 23980 21570
rect 24032 21616 24084 21622
rect 24032 21558 24084 21564
rect 23676 20942 23704 21542
rect 23756 21480 23808 21486
rect 23756 21422 23808 21428
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23572 20596 23624 20602
rect 23572 20538 23624 20544
rect 23664 19916 23716 19922
rect 23664 19858 23716 19864
rect 23480 19848 23532 19854
rect 23480 19790 23532 19796
rect 23492 19378 23520 19790
rect 23572 19780 23624 19786
rect 23572 19722 23624 19728
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23480 18760 23532 18766
rect 23480 18702 23532 18708
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 23492 18426 23520 18702
rect 23480 18420 23532 18426
rect 23480 18362 23532 18368
rect 23584 18290 23612 19722
rect 23676 19242 23704 19858
rect 23768 19378 23796 21422
rect 24044 21128 24072 21558
rect 23952 21100 24072 21128
rect 23952 20466 23980 21100
rect 24504 21078 24532 26862
rect 24584 26852 24636 26858
rect 24584 26794 24636 26800
rect 24596 26586 24624 26794
rect 24584 26580 24636 26586
rect 24584 26522 24636 26528
rect 24780 25498 24808 26862
rect 24860 26784 24912 26790
rect 24860 26726 24912 26732
rect 24872 26450 24900 26726
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24964 26382 24992 29446
rect 25056 29306 25084 29990
rect 25240 29850 25268 29990
rect 25516 29850 25544 30670
rect 26240 30592 26292 30598
rect 26240 30534 26292 30540
rect 25780 30320 25832 30326
rect 25780 30262 25832 30268
rect 25228 29844 25280 29850
rect 25228 29786 25280 29792
rect 25504 29844 25556 29850
rect 25504 29786 25556 29792
rect 25136 29708 25188 29714
rect 25136 29650 25188 29656
rect 25044 29300 25096 29306
rect 25044 29242 25096 29248
rect 25148 28994 25176 29650
rect 25792 29578 25820 30262
rect 26252 29782 26280 30534
rect 26240 29776 26292 29782
rect 26240 29718 26292 29724
rect 26148 29640 26200 29646
rect 26148 29582 26200 29588
rect 26240 29640 26292 29646
rect 26240 29582 26292 29588
rect 25780 29572 25832 29578
rect 25780 29514 25832 29520
rect 26160 29306 26188 29582
rect 26148 29300 26200 29306
rect 26148 29242 26200 29248
rect 25148 28966 25452 28994
rect 25228 28552 25280 28558
rect 25228 28494 25280 28500
rect 25240 28218 25268 28494
rect 25228 28212 25280 28218
rect 25228 28154 25280 28160
rect 25042 28112 25098 28121
rect 25042 28047 25044 28056
rect 25096 28047 25098 28056
rect 25044 28018 25096 28024
rect 25136 27872 25188 27878
rect 25136 27814 25188 27820
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 24860 26240 24912 26246
rect 24860 26182 24912 26188
rect 24872 25906 24900 26182
rect 24860 25900 24912 25906
rect 24860 25842 24912 25848
rect 24768 25492 24820 25498
rect 24768 25434 24820 25440
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24872 24750 24900 25298
rect 24860 24744 24912 24750
rect 24860 24686 24912 24692
rect 25044 23588 25096 23594
rect 25044 23530 25096 23536
rect 25056 23322 25084 23530
rect 25044 23316 25096 23322
rect 25044 23258 25096 23264
rect 24768 22976 24820 22982
rect 24768 22918 24820 22924
rect 24780 22778 24808 22918
rect 24768 22772 24820 22778
rect 24768 22714 24820 22720
rect 25148 22234 25176 27814
rect 25424 26246 25452 28966
rect 26148 28960 26200 28966
rect 26148 28902 26200 28908
rect 25872 28552 25924 28558
rect 25872 28494 25924 28500
rect 25884 28218 25912 28494
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 26160 28014 26188 28902
rect 26148 28008 26200 28014
rect 26148 27950 26200 27956
rect 26160 27606 26188 27950
rect 26148 27600 26200 27606
rect 26148 27542 26200 27548
rect 25688 26920 25740 26926
rect 25688 26862 25740 26868
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25412 25764 25464 25770
rect 25412 25706 25464 25712
rect 25320 25288 25372 25294
rect 25320 25230 25372 25236
rect 25332 23050 25360 25230
rect 25424 24954 25452 25706
rect 25700 25498 25728 26862
rect 26252 26858 26280 29582
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 26344 27130 26372 27406
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26240 26852 26292 26858
rect 26240 26794 26292 26800
rect 26332 26852 26384 26858
rect 26332 26794 26384 26800
rect 25872 26512 25924 26518
rect 25872 26454 25924 26460
rect 25884 26042 25912 26454
rect 25964 26376 26016 26382
rect 26252 26330 26280 26794
rect 25964 26318 26016 26324
rect 25872 26036 25924 26042
rect 25872 25978 25924 25984
rect 25688 25492 25740 25498
rect 25688 25434 25740 25440
rect 25412 24948 25464 24954
rect 25412 24890 25464 24896
rect 25596 24676 25648 24682
rect 25596 24618 25648 24624
rect 25412 23860 25464 23866
rect 25412 23802 25464 23808
rect 25424 23118 25452 23802
rect 25608 23730 25636 24618
rect 25596 23724 25648 23730
rect 25596 23666 25648 23672
rect 25412 23112 25464 23118
rect 25412 23054 25464 23060
rect 25872 23112 25924 23118
rect 25872 23054 25924 23060
rect 25320 23044 25372 23050
rect 25320 22986 25372 22992
rect 25688 23044 25740 23050
rect 25688 22986 25740 22992
rect 25412 22568 25464 22574
rect 25412 22510 25464 22516
rect 25424 22234 25452 22510
rect 25700 22438 25728 22986
rect 25884 22778 25912 23054
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25688 22432 25740 22438
rect 25688 22374 25740 22380
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25412 22228 25464 22234
rect 25412 22170 25464 22176
rect 25700 22030 25728 22374
rect 25976 22234 26004 26318
rect 26160 26302 26280 26330
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 25964 22228 26016 22234
rect 25964 22170 26016 22176
rect 26068 22137 26096 26182
rect 26160 25838 26188 26302
rect 26240 26240 26292 26246
rect 26240 26182 26292 26188
rect 26148 25832 26200 25838
rect 26148 25774 26200 25780
rect 26252 25702 26280 26182
rect 26344 26042 26372 26794
rect 26436 26042 26464 31742
rect 26516 31680 26568 31686
rect 26516 31622 26568 31628
rect 26528 31346 26556 31622
rect 26804 31482 26832 32506
rect 28264 32224 28316 32230
rect 28264 32166 28316 32172
rect 28816 32224 28868 32230
rect 28816 32166 28868 32172
rect 29184 32224 29236 32230
rect 29184 32166 29236 32172
rect 27620 31884 27672 31890
rect 27620 31826 27672 31832
rect 27528 31748 27580 31754
rect 27528 31690 27580 31696
rect 26884 31680 26936 31686
rect 26884 31622 26936 31628
rect 26792 31476 26844 31482
rect 26792 31418 26844 31424
rect 26516 31340 26568 31346
rect 26516 31282 26568 31288
rect 26804 30258 26832 31418
rect 26896 31346 26924 31622
rect 26884 31340 26936 31346
rect 26884 31282 26936 31288
rect 27540 30938 27568 31690
rect 27528 30932 27580 30938
rect 27528 30874 27580 30880
rect 26792 30252 26844 30258
rect 26792 30194 26844 30200
rect 26700 30184 26752 30190
rect 26700 30126 26752 30132
rect 26712 28014 26740 30126
rect 26804 29034 26832 30194
rect 26884 30048 26936 30054
rect 26884 29990 26936 29996
rect 26896 29782 26924 29990
rect 26884 29776 26936 29782
rect 26884 29718 26936 29724
rect 27540 29510 27568 30874
rect 27632 30598 27660 31826
rect 27804 31680 27856 31686
rect 27804 31622 27856 31628
rect 27816 31210 27844 31622
rect 27804 31204 27856 31210
rect 27804 31146 27856 31152
rect 27804 30796 27856 30802
rect 27804 30738 27856 30744
rect 27620 30592 27672 30598
rect 27620 30534 27672 30540
rect 27620 30048 27672 30054
rect 27620 29990 27672 29996
rect 27712 30048 27764 30054
rect 27712 29990 27764 29996
rect 27528 29504 27580 29510
rect 27528 29446 27580 29452
rect 27540 29170 27568 29446
rect 27528 29164 27580 29170
rect 27528 29106 27580 29112
rect 27252 29096 27304 29102
rect 27252 29038 27304 29044
rect 26792 29028 26844 29034
rect 26792 28970 26844 28976
rect 26700 28008 26752 28014
rect 26700 27950 26752 27956
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 26332 26036 26384 26042
rect 26332 25978 26384 25984
rect 26424 26036 26476 26042
rect 26424 25978 26476 25984
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 26528 25838 26556 25910
rect 26516 25832 26568 25838
rect 26712 25809 26740 27270
rect 26804 26450 26832 28970
rect 27264 28762 27292 29038
rect 27436 28960 27488 28966
rect 27436 28902 27488 28908
rect 27252 28756 27304 28762
rect 27252 28698 27304 28704
rect 26884 28688 26936 28694
rect 26884 28630 26936 28636
rect 26896 28218 26924 28630
rect 27448 28626 27476 28902
rect 27540 28626 27568 29106
rect 27632 28642 27660 29990
rect 27724 29578 27752 29990
rect 27816 29850 27844 30738
rect 28276 30734 28304 32166
rect 28540 31884 28592 31890
rect 28540 31826 28592 31832
rect 28552 31754 28580 31826
rect 28552 31726 28764 31754
rect 28736 31210 28764 31726
rect 28724 31204 28776 31210
rect 28724 31146 28776 31152
rect 28540 31136 28592 31142
rect 28540 31078 28592 31084
rect 28552 30938 28580 31078
rect 28540 30932 28592 30938
rect 28540 30874 28592 30880
rect 28264 30728 28316 30734
rect 28264 30670 28316 30676
rect 28540 30184 28592 30190
rect 28540 30126 28592 30132
rect 27988 30048 28040 30054
rect 27988 29990 28040 29996
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27712 29572 27764 29578
rect 27712 29514 27764 29520
rect 27724 29073 27752 29514
rect 27710 29064 27766 29073
rect 27710 28999 27766 29008
rect 27816 28762 27844 29786
rect 27896 29708 27948 29714
rect 27896 29650 27948 29656
rect 27804 28756 27856 28762
rect 27804 28698 27856 28704
rect 27632 28626 27844 28642
rect 27908 28626 27936 29650
rect 28000 29170 28028 29990
rect 28552 29850 28580 30126
rect 28540 29844 28592 29850
rect 28540 29786 28592 29792
rect 27988 29164 28040 29170
rect 27988 29106 28040 29112
rect 28448 29164 28500 29170
rect 28448 29106 28500 29112
rect 28264 28960 28316 28966
rect 28264 28902 28316 28908
rect 28276 28762 28304 28902
rect 28264 28756 28316 28762
rect 28264 28698 28316 28704
rect 27436 28620 27488 28626
rect 27436 28562 27488 28568
rect 27528 28620 27580 28626
rect 27632 28620 27856 28626
rect 27632 28614 27804 28620
rect 27528 28562 27580 28568
rect 27804 28562 27856 28568
rect 27896 28620 27948 28626
rect 27896 28562 27948 28568
rect 26884 28212 26936 28218
rect 26884 28154 26936 28160
rect 27540 27946 27568 28562
rect 27816 28422 27844 28562
rect 27804 28416 27856 28422
rect 27804 28358 27856 28364
rect 27528 27940 27580 27946
rect 27528 27882 27580 27888
rect 27620 27940 27672 27946
rect 27620 27882 27672 27888
rect 27160 27464 27212 27470
rect 27160 27406 27212 27412
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 27080 26994 27108 27270
rect 27068 26988 27120 26994
rect 27068 26930 27120 26936
rect 26884 26852 26936 26858
rect 26884 26794 26936 26800
rect 26896 26586 26924 26794
rect 26976 26784 27028 26790
rect 26976 26726 27028 26732
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 26792 26444 26844 26450
rect 26792 26386 26844 26392
rect 26792 26308 26844 26314
rect 26792 26250 26844 26256
rect 26516 25774 26568 25780
rect 26698 25800 26754 25809
rect 26240 25696 26292 25702
rect 26240 25638 26292 25644
rect 26252 24342 26280 25638
rect 26240 24336 26292 24342
rect 26240 24278 26292 24284
rect 26332 23656 26384 23662
rect 26332 23598 26384 23604
rect 26344 23322 26372 23598
rect 26332 23316 26384 23322
rect 26332 23258 26384 23264
rect 26528 23202 26556 25774
rect 26698 25735 26754 25744
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26620 24070 26648 25638
rect 26700 25288 26752 25294
rect 26700 25230 26752 25236
rect 26608 24064 26660 24070
rect 26606 24032 26608 24041
rect 26660 24032 26662 24041
rect 26606 23967 26662 23976
rect 26712 23662 26740 25230
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26608 23316 26660 23322
rect 26712 23304 26740 23598
rect 26660 23276 26740 23304
rect 26608 23258 26660 23264
rect 26528 23174 26648 23202
rect 26516 23112 26568 23118
rect 26516 23054 26568 23060
rect 26332 22568 26384 22574
rect 26332 22510 26384 22516
rect 26344 22234 26372 22510
rect 26528 22506 26556 23054
rect 26424 22500 26476 22506
rect 26424 22442 26476 22448
rect 26516 22500 26568 22506
rect 26516 22442 26568 22448
rect 26436 22234 26464 22442
rect 26332 22228 26384 22234
rect 26332 22170 26384 22176
rect 26424 22228 26476 22234
rect 26424 22170 26476 22176
rect 26054 22128 26110 22137
rect 26054 22063 26110 22072
rect 25688 22024 25740 22030
rect 25688 21966 25740 21972
rect 24492 21072 24544 21078
rect 24492 21014 24544 21020
rect 24768 21072 24820 21078
rect 24768 21014 24820 21020
rect 24032 21004 24084 21010
rect 24032 20946 24084 20952
rect 24044 20806 24072 20946
rect 24032 20800 24084 20806
rect 24032 20742 24084 20748
rect 24492 20800 24544 20806
rect 24492 20742 24544 20748
rect 24504 20466 24532 20742
rect 23940 20460 23992 20466
rect 23940 20402 23992 20408
rect 24124 20460 24176 20466
rect 24124 20402 24176 20408
rect 24492 20460 24544 20466
rect 24492 20402 24544 20408
rect 24136 20262 24164 20402
rect 23848 20256 23900 20262
rect 23848 20198 23900 20204
rect 24124 20256 24176 20262
rect 24124 20198 24176 20204
rect 24676 20256 24728 20262
rect 24676 20198 24728 20204
rect 23860 19922 23888 20198
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23664 19236 23716 19242
rect 23664 19178 23716 19184
rect 24136 18834 24164 20198
rect 24688 19990 24716 20198
rect 24676 19984 24728 19990
rect 24676 19926 24728 19932
rect 24124 18828 24176 18834
rect 24124 18770 24176 18776
rect 23940 18692 23992 18698
rect 23940 18634 23992 18640
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23480 18148 23532 18154
rect 23480 18090 23532 18096
rect 22988 17980 23296 17989
rect 22988 17978 22994 17980
rect 23050 17978 23074 17980
rect 23130 17978 23154 17980
rect 23210 17978 23234 17980
rect 23290 17978 23296 17980
rect 23050 17926 23052 17978
rect 23232 17926 23234 17978
rect 22988 17924 22994 17926
rect 23050 17924 23074 17926
rect 23130 17924 23154 17926
rect 23210 17924 23234 17926
rect 23290 17924 23296 17926
rect 22988 17915 23296 17924
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 22650 17776 22706 17785
rect 22848 17768 22968 17796
rect 22650 17711 22706 17720
rect 22940 17626 22968 17768
rect 22664 17598 22968 17626
rect 23020 17672 23072 17678
rect 23020 17614 23072 17620
rect 22328 17436 22636 17445
rect 22328 17434 22334 17436
rect 22390 17434 22414 17436
rect 22470 17434 22494 17436
rect 22550 17434 22574 17436
rect 22630 17434 22636 17436
rect 22390 17382 22392 17434
rect 22572 17382 22574 17434
rect 22328 17380 22334 17382
rect 22390 17380 22414 17382
rect 22470 17380 22494 17382
rect 22550 17380 22574 17382
rect 22630 17380 22636 17382
rect 22328 17371 22636 17380
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22376 17264 22428 17270
rect 22376 17206 22428 17212
rect 22296 17134 22324 17206
rect 22192 17128 22244 17134
rect 22192 17070 22244 17076
rect 22284 17128 22336 17134
rect 22284 17070 22336 17076
rect 22388 16794 22416 17206
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22388 16538 22416 16730
rect 22204 16510 22416 16538
rect 22204 15570 22232 16510
rect 22572 16454 22600 17138
rect 22560 16448 22612 16454
rect 22560 16390 22612 16396
rect 22328 16348 22636 16357
rect 22328 16346 22334 16348
rect 22390 16346 22414 16348
rect 22470 16346 22494 16348
rect 22550 16346 22574 16348
rect 22630 16346 22636 16348
rect 22390 16294 22392 16346
rect 22572 16294 22574 16346
rect 22328 16292 22334 16294
rect 22390 16292 22414 16294
rect 22470 16292 22494 16294
rect 22550 16292 22574 16294
rect 22630 16292 22636 16294
rect 22328 16283 22636 16292
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 22112 15422 22232 15450
rect 22100 14884 22152 14890
rect 22100 14826 22152 14832
rect 22008 14816 22060 14822
rect 22008 14758 22060 14764
rect 22020 13870 22048 14758
rect 22112 14006 22140 14826
rect 22204 14793 22232 15422
rect 22328 15260 22636 15269
rect 22328 15258 22334 15260
rect 22390 15258 22414 15260
rect 22470 15258 22494 15260
rect 22550 15258 22574 15260
rect 22630 15258 22636 15260
rect 22390 15206 22392 15258
rect 22572 15206 22574 15258
rect 22328 15204 22334 15206
rect 22390 15204 22414 15206
rect 22470 15204 22494 15206
rect 22550 15204 22574 15206
rect 22630 15204 22636 15206
rect 22328 15195 22636 15204
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22190 14784 22246 14793
rect 22190 14719 22246 14728
rect 22480 14618 22508 14894
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22204 14362 22232 14554
rect 22480 14482 22508 14554
rect 22664 14482 22692 17598
rect 22836 17332 22888 17338
rect 22836 17274 22888 17280
rect 22848 16794 22876 17274
rect 23032 17202 23060 17614
rect 23020 17196 23072 17202
rect 23020 17138 23072 17144
rect 23308 17048 23336 17818
rect 23492 17542 23520 18090
rect 23480 17536 23532 17542
rect 23480 17478 23532 17484
rect 23308 17020 23428 17048
rect 22988 16892 23296 16901
rect 22988 16890 22994 16892
rect 23050 16890 23074 16892
rect 23130 16890 23154 16892
rect 23210 16890 23234 16892
rect 23290 16890 23296 16892
rect 23050 16838 23052 16890
rect 23232 16838 23234 16890
rect 22988 16836 22994 16838
rect 23050 16836 23074 16838
rect 23130 16836 23154 16838
rect 23210 16836 23234 16838
rect 23290 16836 23296 16838
rect 22988 16827 23296 16836
rect 22836 16788 22888 16794
rect 22836 16730 22888 16736
rect 23400 16590 23428 17020
rect 23492 16658 23520 17478
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23584 16522 23612 18226
rect 23756 16992 23808 16998
rect 23756 16934 23808 16940
rect 23848 16992 23900 16998
rect 23848 16934 23900 16940
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22652 14476 22704 14482
rect 22652 14418 22704 14424
rect 22204 14346 22324 14362
rect 22204 14340 22336 14346
rect 22204 14334 22284 14340
rect 22284 14282 22336 14288
rect 22192 14272 22244 14278
rect 22192 14214 22244 14220
rect 22100 14000 22152 14006
rect 22100 13942 22152 13948
rect 22008 13864 22060 13870
rect 22008 13806 22060 13812
rect 22008 13728 22060 13734
rect 22006 13696 22008 13705
rect 22060 13696 22062 13705
rect 22006 13631 22062 13640
rect 22008 13320 22060 13326
rect 22008 13262 22060 13268
rect 22020 12986 22048 13262
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22112 12986 22140 13126
rect 22204 12986 22232 14214
rect 22328 14172 22636 14181
rect 22328 14170 22334 14172
rect 22390 14170 22414 14172
rect 22470 14170 22494 14172
rect 22550 14170 22574 14172
rect 22630 14170 22636 14172
rect 22390 14118 22392 14170
rect 22572 14118 22574 14170
rect 22328 14116 22334 14118
rect 22390 14116 22414 14118
rect 22470 14116 22494 14118
rect 22550 14116 22574 14118
rect 22630 14116 22636 14118
rect 22328 14107 22636 14116
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22296 13190 22324 13874
rect 22388 13190 22416 13942
rect 22848 13410 22876 16390
rect 23584 16250 23612 16458
rect 23572 16244 23624 16250
rect 23572 16186 23624 16192
rect 23768 16114 23796 16934
rect 23860 16794 23888 16934
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23848 16652 23900 16658
rect 23848 16594 23900 16600
rect 23756 16108 23808 16114
rect 23756 16050 23808 16056
rect 23756 15972 23808 15978
rect 23756 15914 23808 15920
rect 22988 15804 23296 15813
rect 22988 15802 22994 15804
rect 23050 15802 23074 15804
rect 23130 15802 23154 15804
rect 23210 15802 23234 15804
rect 23290 15802 23296 15804
rect 23050 15750 23052 15802
rect 23232 15750 23234 15802
rect 22988 15748 22994 15750
rect 23050 15748 23074 15750
rect 23130 15748 23154 15750
rect 23210 15748 23234 15750
rect 23290 15748 23296 15750
rect 22988 15739 23296 15748
rect 23768 15706 23796 15914
rect 23756 15700 23808 15706
rect 23756 15642 23808 15648
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23756 15564 23808 15570
rect 23860 15552 23888 16594
rect 23808 15524 23888 15552
rect 23756 15506 23808 15512
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23400 14822 23428 15302
rect 23492 15162 23520 15506
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 22988 14716 23296 14725
rect 22988 14714 22994 14716
rect 23050 14714 23074 14716
rect 23130 14714 23154 14716
rect 23210 14714 23234 14716
rect 23290 14714 23296 14716
rect 23050 14662 23052 14714
rect 23232 14662 23234 14714
rect 22988 14660 22994 14662
rect 23050 14660 23074 14662
rect 23130 14660 23154 14662
rect 23210 14660 23234 14662
rect 23290 14660 23296 14662
rect 22988 14651 23296 14660
rect 23400 14414 23428 14758
rect 23768 14482 23796 15506
rect 23952 14521 23980 18634
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24412 18290 24440 18566
rect 24400 18284 24452 18290
rect 24400 18226 24452 18232
rect 24216 17808 24268 17814
rect 24216 17750 24268 17756
rect 24228 16794 24256 17750
rect 24308 17128 24360 17134
rect 24308 17070 24360 17076
rect 24400 17128 24452 17134
rect 24400 17070 24452 17076
rect 24320 16794 24348 17070
rect 24216 16788 24268 16794
rect 24216 16730 24268 16736
rect 24308 16788 24360 16794
rect 24308 16730 24360 16736
rect 24412 16658 24440 17070
rect 24400 16652 24452 16658
rect 24400 16594 24452 16600
rect 24584 16244 24636 16250
rect 24584 16186 24636 16192
rect 24400 15972 24452 15978
rect 24400 15914 24452 15920
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 24044 15706 24072 15846
rect 24032 15700 24084 15706
rect 24032 15642 24084 15648
rect 24044 14618 24072 15642
rect 24412 15094 24440 15914
rect 24400 15088 24452 15094
rect 24400 15030 24452 15036
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 23938 14512 23994 14521
rect 23756 14476 23808 14482
rect 23938 14447 23994 14456
rect 23756 14418 23808 14424
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 22940 13938 22968 14214
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 23216 13870 23244 14350
rect 23388 14272 23440 14278
rect 23388 14214 23440 14220
rect 23400 13977 23428 14214
rect 23386 13968 23442 13977
rect 23386 13903 23388 13912
rect 23440 13903 23442 13912
rect 23480 13932 23532 13938
rect 23388 13874 23440 13880
rect 23480 13874 23532 13880
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 22988 13628 23296 13637
rect 22988 13626 22994 13628
rect 23050 13626 23074 13628
rect 23130 13626 23154 13628
rect 23210 13626 23234 13628
rect 23290 13626 23296 13628
rect 23050 13574 23052 13626
rect 23232 13574 23234 13626
rect 22988 13572 22994 13574
rect 23050 13572 23074 13574
rect 23130 13572 23154 13574
rect 23210 13572 23234 13574
rect 23290 13572 23296 13574
rect 22988 13563 23296 13572
rect 23492 13530 23520 13874
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 22652 13388 22704 13394
rect 22848 13382 22968 13410
rect 22652 13330 22704 13336
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22376 13184 22428 13190
rect 22376 13126 22428 13132
rect 22328 13084 22636 13093
rect 22328 13082 22334 13084
rect 22390 13082 22414 13084
rect 22470 13082 22494 13084
rect 22550 13082 22574 13084
rect 22630 13082 22636 13084
rect 22390 13030 22392 13082
rect 22572 13030 22574 13082
rect 22328 13028 22334 13030
rect 22390 13028 22414 13030
rect 22470 13028 22494 13030
rect 22550 13028 22574 13030
rect 22630 13028 22636 13030
rect 22328 13019 22636 13028
rect 22008 12980 22060 12986
rect 22008 12922 22060 12928
rect 22100 12980 22152 12986
rect 22100 12922 22152 12928
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21916 11892 21968 11898
rect 21916 11834 21968 11840
rect 21824 9988 21876 9994
rect 21824 9930 21876 9936
rect 21732 9444 21784 9450
rect 21732 9386 21784 9392
rect 21744 8634 21772 9386
rect 21824 9376 21876 9382
rect 21824 9318 21876 9324
rect 21836 8974 21864 9318
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21928 8537 21956 11834
rect 22020 11665 22048 12174
rect 22328 11996 22636 12005
rect 22328 11994 22334 11996
rect 22390 11994 22414 11996
rect 22470 11994 22494 11996
rect 22550 11994 22574 11996
rect 22630 11994 22636 11996
rect 22390 11942 22392 11994
rect 22572 11942 22574 11994
rect 22328 11940 22334 11942
rect 22390 11940 22414 11942
rect 22470 11940 22494 11942
rect 22550 11940 22574 11942
rect 22630 11940 22636 11942
rect 22328 11931 22636 11940
rect 22664 11898 22692 13330
rect 22836 12980 22888 12986
rect 22836 12922 22888 12928
rect 22744 12776 22796 12782
rect 22744 12718 22796 12724
rect 22756 12102 22784 12718
rect 22744 12096 22796 12102
rect 22744 12038 22796 12044
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22848 11762 22876 12922
rect 22940 12782 22968 13382
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 23308 12986 23336 13126
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23756 12844 23808 12850
rect 23756 12786 23808 12792
rect 22928 12776 22980 12782
rect 22928 12718 22980 12724
rect 23768 12714 23796 12786
rect 23756 12708 23808 12714
rect 23756 12650 23808 12656
rect 22988 12540 23296 12549
rect 22988 12538 22994 12540
rect 23050 12538 23074 12540
rect 23130 12538 23154 12540
rect 23210 12538 23234 12540
rect 23290 12538 23296 12540
rect 23050 12486 23052 12538
rect 23232 12486 23234 12538
rect 22988 12484 22994 12486
rect 23050 12484 23074 12486
rect 23130 12484 23154 12486
rect 23210 12484 23234 12486
rect 23290 12484 23296 12486
rect 22988 12475 23296 12484
rect 23860 12434 23888 13262
rect 23952 13002 23980 14447
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24504 14074 24532 14282
rect 24492 14068 24544 14074
rect 24492 14010 24544 14016
rect 24228 13938 24440 13954
rect 24216 13932 24440 13938
rect 24268 13926 24440 13932
rect 24216 13874 24268 13880
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24044 13326 24072 13670
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24136 13190 24164 13806
rect 24216 13728 24268 13734
rect 24216 13670 24268 13676
rect 24228 13530 24256 13670
rect 24216 13524 24268 13530
rect 24216 13466 24268 13472
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 23952 12974 24164 13002
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 23952 12442 23980 12650
rect 23768 12406 23888 12434
rect 23940 12436 23992 12442
rect 23768 12374 23796 12406
rect 24136 12434 24164 12974
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24320 12434 24348 12582
rect 23940 12378 23992 12384
rect 24044 12406 24164 12434
rect 24228 12406 24348 12434
rect 23756 12368 23808 12374
rect 23570 12336 23626 12345
rect 23756 12310 23808 12316
rect 23570 12271 23572 12280
rect 23624 12271 23626 12280
rect 23572 12242 23624 12248
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 22836 11756 22888 11762
rect 22836 11698 22888 11704
rect 22100 11688 22152 11694
rect 22006 11656 22062 11665
rect 22100 11630 22152 11636
rect 22190 11656 22246 11665
rect 22006 11591 22062 11600
rect 22112 10130 22140 11630
rect 22190 11591 22246 11600
rect 22100 10124 22152 10130
rect 22100 10066 22152 10072
rect 22100 9988 22152 9994
rect 22100 9930 22152 9936
rect 22112 8945 22140 9930
rect 22204 9450 22232 11591
rect 22652 11144 22704 11150
rect 22652 11086 22704 11092
rect 22328 10908 22636 10917
rect 22328 10906 22334 10908
rect 22390 10906 22414 10908
rect 22470 10906 22494 10908
rect 22550 10906 22574 10908
rect 22630 10906 22636 10908
rect 22390 10854 22392 10906
rect 22572 10854 22574 10906
rect 22328 10852 22334 10854
rect 22390 10852 22414 10854
rect 22470 10852 22494 10854
rect 22550 10852 22574 10854
rect 22630 10852 22636 10854
rect 22328 10843 22636 10852
rect 22664 9926 22692 11086
rect 22848 10674 22876 11698
rect 22988 11452 23296 11461
rect 22988 11450 22994 11452
rect 23050 11450 23074 11452
rect 23130 11450 23154 11452
rect 23210 11450 23234 11452
rect 23290 11450 23296 11452
rect 23050 11398 23052 11450
rect 23232 11398 23234 11450
rect 22988 11396 22994 11398
rect 23050 11396 23074 11398
rect 23130 11396 23154 11398
rect 23210 11396 23234 11398
rect 23290 11396 23296 11398
rect 22988 11387 23296 11396
rect 23400 11354 23428 12038
rect 22928 11348 22980 11354
rect 22928 11290 22980 11296
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22744 10600 22796 10606
rect 22940 10554 22968 11290
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 23296 11212 23348 11218
rect 23296 11154 23348 11160
rect 23664 11212 23716 11218
rect 23664 11154 23716 11160
rect 23032 10742 23060 11154
rect 23308 11098 23336 11154
rect 23480 11144 23532 11150
rect 23308 11070 23428 11098
rect 23480 11086 23532 11092
rect 23020 10736 23072 10742
rect 23020 10678 23072 10684
rect 22744 10542 22796 10548
rect 22756 10266 22784 10542
rect 22848 10526 22968 10554
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22744 10124 22796 10130
rect 22744 10066 22796 10072
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 22328 9820 22636 9829
rect 22328 9818 22334 9820
rect 22390 9818 22414 9820
rect 22470 9818 22494 9820
rect 22550 9818 22574 9820
rect 22630 9818 22636 9820
rect 22390 9766 22392 9818
rect 22572 9766 22574 9818
rect 22328 9764 22334 9766
rect 22390 9764 22414 9766
rect 22470 9764 22494 9766
rect 22550 9764 22574 9766
rect 22630 9764 22636 9766
rect 22328 9755 22636 9764
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22652 9376 22704 9382
rect 22652 9318 22704 9324
rect 22098 8936 22154 8945
rect 22098 8871 22154 8880
rect 22008 8832 22060 8838
rect 22060 8792 22140 8820
rect 22008 8774 22060 8780
rect 22112 8634 22140 8792
rect 22328 8732 22636 8741
rect 22328 8730 22334 8732
rect 22390 8730 22414 8732
rect 22470 8730 22494 8732
rect 22550 8730 22574 8732
rect 22630 8730 22636 8732
rect 22390 8678 22392 8730
rect 22572 8678 22574 8730
rect 22328 8676 22334 8678
rect 22390 8676 22414 8678
rect 22470 8676 22494 8678
rect 22550 8676 22574 8678
rect 22630 8676 22636 8678
rect 22328 8667 22636 8676
rect 22664 8650 22692 9318
rect 22756 9058 22784 10066
rect 22848 9586 22876 10526
rect 22988 10364 23296 10373
rect 22988 10362 22994 10364
rect 23050 10362 23074 10364
rect 23130 10362 23154 10364
rect 23210 10362 23234 10364
rect 23290 10362 23296 10364
rect 23050 10310 23052 10362
rect 23232 10310 23234 10362
rect 22988 10308 22994 10310
rect 23050 10308 23074 10310
rect 23130 10308 23154 10310
rect 23210 10308 23234 10310
rect 23290 10308 23296 10310
rect 22988 10299 23296 10308
rect 23400 9994 23428 11070
rect 23492 10810 23520 11086
rect 23480 10804 23532 10810
rect 23480 10746 23532 10752
rect 23676 10062 23704 11154
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23952 10538 23980 10950
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 23940 10124 23992 10130
rect 23940 10066 23992 10072
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23756 10056 23808 10062
rect 23756 9998 23808 10004
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22940 9518 22968 9862
rect 23308 9674 23336 9862
rect 23124 9646 23336 9674
rect 23124 9586 23152 9646
rect 23112 9580 23164 9586
rect 23112 9522 23164 9528
rect 22928 9512 22980 9518
rect 22928 9454 22980 9460
rect 22988 9276 23296 9285
rect 22988 9274 22994 9276
rect 23050 9274 23074 9276
rect 23130 9274 23154 9276
rect 23210 9274 23234 9276
rect 23290 9274 23296 9276
rect 23050 9222 23052 9274
rect 23232 9222 23234 9274
rect 22988 9220 22994 9222
rect 23050 9220 23074 9222
rect 23130 9220 23154 9222
rect 23210 9220 23234 9222
rect 23290 9220 23296 9222
rect 22988 9211 23296 9220
rect 22756 9030 22968 9058
rect 22664 8634 22876 8650
rect 22100 8628 22152 8634
rect 22664 8628 22888 8634
rect 22664 8622 22836 8628
rect 22100 8570 22152 8576
rect 22836 8570 22888 8576
rect 21914 8528 21970 8537
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21824 8492 21876 8498
rect 21914 8463 21970 8472
rect 21824 8434 21876 8440
rect 21652 8022 21680 8434
rect 21640 8016 21692 8022
rect 21640 7958 21692 7964
rect 21744 7954 21772 8434
rect 21732 7948 21784 7954
rect 21732 7890 21784 7896
rect 21548 7744 21600 7750
rect 21548 7686 21600 7692
rect 21732 7268 21784 7274
rect 21376 7228 21732 7256
rect 21732 7210 21784 7216
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21560 6458 21588 6598
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21732 6180 21784 6186
rect 21732 6122 21784 6128
rect 21744 5370 21772 6122
rect 21732 5364 21784 5370
rect 21732 5306 21784 5312
rect 21180 4480 21232 4486
rect 21180 4422 21232 4428
rect 21192 4146 21220 4422
rect 21180 4140 21232 4146
rect 21180 4082 21232 4088
rect 21192 2990 21220 4082
rect 21744 4078 21772 5306
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21836 3534 21864 8434
rect 21928 7478 21956 8463
rect 22112 8412 22140 8570
rect 22940 8514 22968 9030
rect 23400 8566 23428 9930
rect 23768 9518 23796 9998
rect 23756 9512 23808 9518
rect 23756 9454 23808 9460
rect 23848 9512 23900 9518
rect 23848 9454 23900 9460
rect 23572 9036 23624 9042
rect 23572 8978 23624 8984
rect 23584 8634 23612 8978
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23388 8560 23440 8566
rect 22848 8486 22968 8514
rect 23110 8528 23166 8537
rect 23388 8502 23440 8508
rect 22284 8424 22336 8430
rect 22112 8384 22284 8412
rect 22284 8366 22336 8372
rect 22848 8090 22876 8486
rect 23110 8463 23112 8472
rect 23164 8463 23166 8472
rect 23112 8434 23164 8440
rect 23386 8392 23442 8401
rect 23386 8327 23442 8336
rect 22988 8188 23296 8197
rect 22988 8186 22994 8188
rect 23050 8186 23074 8188
rect 23130 8186 23154 8188
rect 23210 8186 23234 8188
rect 23290 8186 23296 8188
rect 23050 8134 23052 8186
rect 23232 8134 23234 8186
rect 22988 8132 22994 8134
rect 23050 8132 23074 8134
rect 23130 8132 23154 8134
rect 23210 8132 23234 8134
rect 23290 8132 23296 8134
rect 22988 8123 23296 8132
rect 23400 8090 23428 8327
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22744 7948 22796 7954
rect 22744 7890 22796 7896
rect 22664 7750 22692 7890
rect 22756 7750 22784 7890
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22020 7546 22048 7686
rect 22328 7644 22636 7653
rect 22328 7642 22334 7644
rect 22390 7642 22414 7644
rect 22470 7642 22494 7644
rect 22550 7642 22574 7644
rect 22630 7642 22636 7644
rect 22390 7590 22392 7642
rect 22572 7590 22574 7642
rect 22328 7588 22334 7590
rect 22390 7588 22414 7590
rect 22470 7588 22494 7590
rect 22550 7588 22574 7590
rect 22630 7588 22636 7590
rect 22328 7579 22636 7588
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21916 7472 21968 7478
rect 21916 7414 21968 7420
rect 21928 5914 21956 7414
rect 22468 7336 22520 7342
rect 22468 7278 22520 7284
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 22112 6866 22140 7142
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22204 6118 22232 6802
rect 22480 6662 22508 7278
rect 22468 6656 22520 6662
rect 22468 6598 22520 6604
rect 22328 6556 22636 6565
rect 22328 6554 22334 6556
rect 22390 6554 22414 6556
rect 22470 6554 22494 6556
rect 22550 6554 22574 6556
rect 22630 6554 22636 6556
rect 22390 6502 22392 6554
rect 22572 6502 22574 6554
rect 22328 6500 22334 6502
rect 22390 6500 22414 6502
rect 22470 6500 22494 6502
rect 22550 6500 22574 6502
rect 22630 6500 22636 6502
rect 22328 6491 22636 6500
rect 22192 6112 22244 6118
rect 22192 6054 22244 6060
rect 21916 5908 21968 5914
rect 21916 5850 21968 5856
rect 22204 5778 22232 6054
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22664 5642 22692 7686
rect 23400 7546 23428 8026
rect 23860 7886 23888 9454
rect 23952 8906 23980 10066
rect 23940 8900 23992 8906
rect 23940 8842 23992 8848
rect 23572 7880 23624 7886
rect 23572 7822 23624 7828
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 23388 7540 23440 7546
rect 23388 7482 23440 7488
rect 23480 7200 23532 7206
rect 23480 7142 23532 7148
rect 22988 7100 23296 7109
rect 22988 7098 22994 7100
rect 23050 7098 23074 7100
rect 23130 7098 23154 7100
rect 23210 7098 23234 7100
rect 23290 7098 23296 7100
rect 23050 7046 23052 7098
rect 23232 7046 23234 7098
rect 22988 7044 22994 7046
rect 23050 7044 23074 7046
rect 23130 7044 23154 7046
rect 23210 7044 23234 7046
rect 23290 7044 23296 7046
rect 22988 7035 23296 7044
rect 23020 6792 23072 6798
rect 23020 6734 23072 6740
rect 22836 6656 22888 6662
rect 22836 6598 22888 6604
rect 22652 5636 22704 5642
rect 22652 5578 22704 5584
rect 22328 5468 22636 5477
rect 22328 5466 22334 5468
rect 22390 5466 22414 5468
rect 22470 5466 22494 5468
rect 22550 5466 22574 5468
rect 22630 5466 22636 5468
rect 22390 5414 22392 5466
rect 22572 5414 22574 5466
rect 22328 5412 22334 5414
rect 22390 5412 22414 5414
rect 22470 5412 22494 5414
rect 22550 5412 22574 5414
rect 22630 5412 22636 5414
rect 22328 5403 22636 5412
rect 22848 5234 22876 6598
rect 23032 6458 23060 6734
rect 23492 6458 23520 7142
rect 23584 7002 23612 7822
rect 23756 7744 23808 7750
rect 23756 7686 23808 7692
rect 23572 6996 23624 7002
rect 23572 6938 23624 6944
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23584 6254 23612 6938
rect 23768 6866 23796 7686
rect 23860 7410 23888 7822
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23860 6322 23888 7346
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 24044 6254 24072 12406
rect 24124 12300 24176 12306
rect 24124 12242 24176 12248
rect 24136 7478 24164 12242
rect 24228 11762 24256 12406
rect 24216 11756 24268 11762
rect 24216 11698 24268 11704
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24228 10674 24256 10950
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24216 8628 24268 8634
rect 24216 8570 24268 8576
rect 24124 7472 24176 7478
rect 24124 7414 24176 7420
rect 24122 6896 24178 6905
rect 24122 6831 24124 6840
rect 24176 6831 24178 6840
rect 24124 6802 24176 6808
rect 23572 6248 23624 6254
rect 23572 6190 23624 6196
rect 23664 6248 23716 6254
rect 23664 6190 23716 6196
rect 23756 6248 23808 6254
rect 23756 6190 23808 6196
rect 24032 6248 24084 6254
rect 24032 6190 24084 6196
rect 23388 6112 23440 6118
rect 23388 6054 23440 6060
rect 22988 6012 23296 6021
rect 22988 6010 22994 6012
rect 23050 6010 23074 6012
rect 23130 6010 23154 6012
rect 23210 6010 23234 6012
rect 23290 6010 23296 6012
rect 23050 5958 23052 6010
rect 23232 5958 23234 6010
rect 22988 5956 22994 5958
rect 23050 5956 23074 5958
rect 23130 5956 23154 5958
rect 23210 5956 23234 5958
rect 23290 5956 23296 5958
rect 22988 5947 23296 5956
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 23400 5166 23428 6054
rect 23584 5370 23612 6190
rect 23676 6118 23704 6190
rect 23664 6112 23716 6118
rect 23664 6054 23716 6060
rect 23676 5846 23704 6054
rect 23664 5840 23716 5846
rect 23664 5782 23716 5788
rect 23768 5370 23796 6190
rect 24228 5778 24256 8570
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24320 8090 24348 8230
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 24320 6254 24348 7142
rect 24308 6248 24360 6254
rect 24308 6190 24360 6196
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 24228 5370 24256 5714
rect 24308 5704 24360 5710
rect 24308 5646 24360 5652
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 24216 5364 24268 5370
rect 24216 5306 24268 5312
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 22988 4924 23296 4933
rect 22988 4922 22994 4924
rect 23050 4922 23074 4924
rect 23130 4922 23154 4924
rect 23210 4922 23234 4924
rect 23290 4922 23296 4924
rect 23050 4870 23052 4922
rect 23232 4870 23234 4922
rect 22988 4868 22994 4870
rect 23050 4868 23074 4870
rect 23130 4868 23154 4870
rect 23210 4868 23234 4870
rect 23290 4868 23296 4870
rect 22988 4859 23296 4868
rect 23400 4826 23428 5102
rect 23388 4820 23440 4826
rect 23388 4762 23440 4768
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22328 4380 22636 4389
rect 22328 4378 22334 4380
rect 22390 4378 22414 4380
rect 22470 4378 22494 4380
rect 22550 4378 22574 4380
rect 22630 4378 22636 4380
rect 22390 4326 22392 4378
rect 22572 4326 22574 4378
rect 22328 4324 22334 4326
rect 22390 4324 22414 4326
rect 22470 4324 22494 4326
rect 22550 4324 22574 4326
rect 22630 4324 22636 4326
rect 22328 4315 22636 4324
rect 22848 3942 22876 4558
rect 23664 4480 23716 4486
rect 23664 4422 23716 4428
rect 23676 3942 23704 4422
rect 23768 4078 23796 5306
rect 23848 5024 23900 5030
rect 23848 4966 23900 4972
rect 23860 4690 23888 4966
rect 23848 4684 23900 4690
rect 23848 4626 23900 4632
rect 23756 4072 23808 4078
rect 23756 4014 23808 4020
rect 22836 3936 22888 3942
rect 22836 3878 22888 3884
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 22988 3836 23296 3845
rect 22988 3834 22994 3836
rect 23050 3834 23074 3836
rect 23130 3834 23154 3836
rect 23210 3834 23234 3836
rect 23290 3834 23296 3836
rect 23050 3782 23052 3834
rect 23232 3782 23234 3834
rect 22988 3780 22994 3782
rect 23050 3780 23074 3782
rect 23130 3780 23154 3782
rect 23210 3780 23234 3782
rect 23290 3780 23296 3782
rect 22988 3771 23296 3780
rect 21824 3528 21876 3534
rect 21824 3470 21876 3476
rect 22328 3292 22636 3301
rect 22328 3290 22334 3292
rect 22390 3290 22414 3292
rect 22470 3290 22494 3292
rect 22550 3290 22574 3292
rect 22630 3290 22636 3292
rect 22390 3238 22392 3290
rect 22572 3238 22574 3290
rect 22328 3236 22334 3238
rect 22390 3236 22414 3238
rect 22470 3236 22494 3238
rect 22550 3236 22574 3238
rect 22630 3236 22636 3238
rect 22328 3227 22636 3236
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 22020 1442 22048 2994
rect 23676 2990 23704 3878
rect 24320 3126 24348 5646
rect 24412 3466 24440 13926
rect 24596 13716 24624 16186
rect 24676 14884 24728 14890
rect 24676 14826 24728 14832
rect 24688 14618 24716 14826
rect 24676 14612 24728 14618
rect 24676 14554 24728 14560
rect 24504 13688 24624 13716
rect 24504 13326 24532 13688
rect 24676 13388 24728 13394
rect 24676 13330 24728 13336
rect 24492 13320 24544 13326
rect 24492 13262 24544 13268
rect 24504 11150 24532 13262
rect 24688 12918 24716 13330
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24688 12434 24716 12854
rect 24596 12406 24716 12434
rect 24596 12306 24624 12406
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 24780 9217 24808 21014
rect 25596 21004 25648 21010
rect 25596 20946 25648 20952
rect 25608 20602 25636 20946
rect 25596 20596 25648 20602
rect 25596 20538 25648 20544
rect 25320 19984 25372 19990
rect 25320 19926 25372 19932
rect 24952 19712 25004 19718
rect 24952 19654 25004 19660
rect 24964 19514 24992 19654
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 25332 19310 25360 19926
rect 25700 19922 25728 21966
rect 26056 21548 26108 21554
rect 26056 21490 26108 21496
rect 25780 21480 25832 21486
rect 25780 21422 25832 21428
rect 25792 20806 25820 21422
rect 26068 21078 26096 21490
rect 26148 21480 26200 21486
rect 26200 21428 26280 21434
rect 26148 21422 26280 21428
rect 26160 21406 26280 21422
rect 26056 21072 26108 21078
rect 26056 21014 26108 21020
rect 25780 20800 25832 20806
rect 25780 20742 25832 20748
rect 26252 20602 26280 21406
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26332 20800 26384 20806
rect 26332 20742 26384 20748
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26344 20466 26372 20742
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26056 20392 26108 20398
rect 26056 20334 26108 20340
rect 25780 20324 25832 20330
rect 25780 20266 25832 20272
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25792 19718 25820 20266
rect 26068 19786 26096 20334
rect 26148 20324 26200 20330
rect 26332 20324 26384 20330
rect 26200 20284 26280 20312
rect 26148 20266 26200 20272
rect 26252 19922 26280 20284
rect 26332 20266 26384 20272
rect 26344 20058 26372 20266
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26240 19916 26292 19922
rect 26240 19858 26292 19864
rect 26056 19780 26108 19786
rect 26056 19722 26108 19728
rect 25780 19712 25832 19718
rect 25780 19654 25832 19660
rect 26252 19502 26372 19530
rect 26436 19514 26464 20538
rect 25320 19304 25372 19310
rect 25320 19246 25372 19252
rect 26056 19168 26108 19174
rect 26056 19110 26108 19116
rect 26068 18970 26096 19110
rect 26056 18964 26108 18970
rect 26056 18906 26108 18912
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 25700 18426 25728 18770
rect 25688 18420 25740 18426
rect 25688 18362 25740 18368
rect 24952 18080 25004 18086
rect 24952 18022 25004 18028
rect 24964 17678 24992 18022
rect 24952 17672 25004 17678
rect 24952 17614 25004 17620
rect 25228 17536 25280 17542
rect 25228 17478 25280 17484
rect 25240 17338 25268 17478
rect 25228 17332 25280 17338
rect 25228 17274 25280 17280
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 25044 16720 25096 16726
rect 25044 16662 25096 16668
rect 25056 16250 25084 16662
rect 25044 16244 25096 16250
rect 25044 16186 25096 16192
rect 24952 16040 25004 16046
rect 24952 15982 25004 15988
rect 24964 14482 24992 15982
rect 25148 15910 25176 17070
rect 25136 15904 25188 15910
rect 25136 15846 25188 15852
rect 24952 14476 25004 14482
rect 24952 14418 25004 14424
rect 24964 12238 24992 14418
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25056 12850 25084 13126
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25240 12442 25268 17274
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25608 16658 25636 16934
rect 25884 16794 25912 17070
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 26056 16176 26108 16182
rect 26056 16118 26108 16124
rect 26068 14550 26096 16118
rect 26148 15904 26200 15910
rect 26148 15846 26200 15852
rect 26056 14544 26108 14550
rect 26056 14486 26108 14492
rect 25780 14476 25832 14482
rect 25780 14418 25832 14424
rect 25964 14476 26016 14482
rect 25964 14418 26016 14424
rect 25792 14074 25820 14418
rect 25976 14074 26004 14418
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 25964 14068 26016 14074
rect 25964 14010 26016 14016
rect 25688 14000 25740 14006
rect 25688 13942 25740 13948
rect 25700 13530 25728 13942
rect 25688 13524 25740 13530
rect 25688 13466 25740 13472
rect 26160 13462 26188 15846
rect 26252 13705 26280 19502
rect 26344 19446 26372 19502
rect 26424 19508 26476 19514
rect 26424 19450 26476 19456
rect 26332 19440 26384 19446
rect 26332 19382 26384 19388
rect 26332 16992 26384 16998
rect 26332 16934 26384 16940
rect 26344 16658 26372 16934
rect 26528 16658 26556 21354
rect 26620 20482 26648 23174
rect 26712 22710 26740 23276
rect 26700 22704 26752 22710
rect 26700 22646 26752 22652
rect 26700 22228 26752 22234
rect 26700 22170 26752 22176
rect 26712 22098 26740 22170
rect 26700 22092 26752 22098
rect 26700 22034 26752 22040
rect 26700 20936 26752 20942
rect 26700 20878 26752 20884
rect 26712 20602 26740 20878
rect 26700 20596 26752 20602
rect 26700 20538 26752 20544
rect 26620 20454 26740 20482
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26620 19718 26648 20334
rect 26608 19712 26660 19718
rect 26608 19654 26660 19660
rect 26712 19446 26740 20454
rect 26804 19922 26832 26250
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26896 21146 26924 25638
rect 26988 25498 27016 26726
rect 27080 26466 27108 26930
rect 27172 26586 27200 27406
rect 27632 27402 27660 27882
rect 27816 27554 27844 28358
rect 27724 27538 27844 27554
rect 27712 27532 27844 27538
rect 27764 27526 27844 27532
rect 27712 27474 27764 27480
rect 27620 27396 27672 27402
rect 27620 27338 27672 27344
rect 27160 26580 27212 26586
rect 27160 26522 27212 26528
rect 27080 26450 27200 26466
rect 27080 26444 27212 26450
rect 27080 26438 27160 26444
rect 27160 26386 27212 26392
rect 27172 25838 27200 26386
rect 27344 25968 27396 25974
rect 27344 25910 27396 25916
rect 27160 25832 27212 25838
rect 27160 25774 27212 25780
rect 27356 25498 27384 25910
rect 26976 25492 27028 25498
rect 26976 25434 27028 25440
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27068 25288 27120 25294
rect 27068 25230 27120 25236
rect 27540 25242 27568 25298
rect 27080 24954 27108 25230
rect 27540 25214 27660 25242
rect 27068 24948 27120 24954
rect 27068 24890 27120 24896
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27172 24138 27200 24550
rect 27160 24132 27212 24138
rect 27160 24074 27212 24080
rect 27632 24070 27660 25214
rect 27724 25158 27752 27474
rect 27908 26042 27936 28562
rect 28460 28490 28488 29106
rect 28632 28620 28684 28626
rect 28632 28562 28684 28568
rect 28448 28484 28500 28490
rect 28448 28426 28500 28432
rect 28356 28212 28408 28218
rect 28356 28154 28408 28160
rect 28172 27668 28224 27674
rect 28172 27610 28224 27616
rect 27986 27568 28042 27577
rect 27986 27503 28042 27512
rect 28000 26790 28028 27503
rect 28184 27334 28212 27610
rect 28368 27606 28396 28154
rect 28356 27600 28408 27606
rect 28356 27542 28408 27548
rect 28644 27538 28672 28562
rect 28828 28218 28856 32166
rect 29196 31958 29224 32166
rect 29184 31952 29236 31958
rect 29184 31894 29236 31900
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 28908 30048 28960 30054
rect 28908 29990 28960 29996
rect 28920 29850 28948 29990
rect 28908 29844 28960 29850
rect 28908 29786 28960 29792
rect 29104 29782 29132 30534
rect 29092 29776 29144 29782
rect 29092 29718 29144 29724
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 29012 28762 29040 28970
rect 29000 28756 29052 28762
rect 29000 28698 29052 28704
rect 28816 28212 28868 28218
rect 28816 28154 28868 28160
rect 28908 28144 28960 28150
rect 28908 28086 28960 28092
rect 28724 28008 28776 28014
rect 28920 27985 28948 28086
rect 28724 27950 28776 27956
rect 28906 27976 28962 27985
rect 28736 27674 28764 27950
rect 28906 27911 28962 27920
rect 28724 27668 28776 27674
rect 28724 27610 28776 27616
rect 28632 27532 28684 27538
rect 28632 27474 28684 27480
rect 28908 27532 28960 27538
rect 28908 27474 28960 27480
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 28080 26988 28132 26994
rect 28080 26930 28132 26936
rect 27988 26784 28040 26790
rect 27988 26726 28040 26732
rect 27896 26036 27948 26042
rect 27896 25978 27948 25984
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 27712 25152 27764 25158
rect 27712 25094 27764 25100
rect 27816 24954 27844 25230
rect 27804 24948 27856 24954
rect 27804 24890 27856 24896
rect 27712 24676 27764 24682
rect 27712 24618 27764 24624
rect 27724 24206 27752 24618
rect 27712 24200 27764 24206
rect 27712 24142 27764 24148
rect 27620 24064 27672 24070
rect 27620 24006 27672 24012
rect 27436 23656 27488 23662
rect 27436 23598 27488 23604
rect 27344 23520 27396 23526
rect 27344 23462 27396 23468
rect 27356 23186 27384 23462
rect 27448 23322 27476 23598
rect 27632 23594 27660 24006
rect 27712 23656 27764 23662
rect 27712 23598 27764 23604
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 27632 23474 27660 23530
rect 27540 23446 27660 23474
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 27344 23180 27396 23186
rect 27344 23122 27396 23128
rect 27068 22500 27120 22506
rect 27068 22442 27120 22448
rect 27080 22098 27108 22442
rect 27160 22432 27212 22438
rect 27160 22374 27212 22380
rect 27068 22092 27120 22098
rect 26988 22052 27068 22080
rect 26988 21962 27016 22052
rect 27068 22034 27120 22040
rect 26976 21956 27028 21962
rect 26976 21898 27028 21904
rect 27068 21956 27120 21962
rect 27068 21898 27120 21904
rect 26884 21140 26936 21146
rect 26884 21082 26936 21088
rect 26988 21010 27016 21898
rect 27080 21010 27108 21898
rect 26976 21004 27028 21010
rect 26976 20946 27028 20952
rect 27068 21004 27120 21010
rect 27068 20946 27120 20952
rect 27172 20602 27200 22374
rect 27448 22234 27476 23258
rect 27436 22228 27488 22234
rect 27436 22170 27488 22176
rect 27344 21004 27396 21010
rect 27344 20946 27396 20952
rect 27252 20936 27304 20942
rect 27252 20878 27304 20884
rect 27160 20596 27212 20602
rect 27160 20538 27212 20544
rect 26792 19916 26844 19922
rect 26792 19858 26844 19864
rect 27068 19780 27120 19786
rect 27068 19722 27120 19728
rect 26792 19508 26844 19514
rect 26792 19450 26844 19456
rect 26700 19440 26752 19446
rect 26700 19382 26752 19388
rect 26804 18222 26832 19450
rect 26608 18216 26660 18222
rect 26608 18158 26660 18164
rect 26792 18216 26844 18222
rect 26792 18158 26844 18164
rect 26620 17338 26648 18158
rect 27080 18086 27108 19722
rect 27172 19310 27200 20538
rect 27160 19304 27212 19310
rect 27160 19246 27212 19252
rect 27264 19242 27292 20878
rect 27356 19922 27384 20946
rect 27540 20398 27568 23446
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 27632 22166 27660 23122
rect 27724 23050 27752 23598
rect 27816 23186 27844 24890
rect 27908 24342 27936 25230
rect 28000 24614 28028 26726
rect 28092 26450 28120 26930
rect 28184 26450 28212 27270
rect 28644 26926 28672 27474
rect 28632 26920 28684 26926
rect 28632 26862 28684 26868
rect 28080 26444 28132 26450
rect 28080 26386 28132 26392
rect 28172 26444 28224 26450
rect 28172 26386 28224 26392
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 27896 24336 27948 24342
rect 27896 24278 27948 24284
rect 28092 23866 28120 26386
rect 28172 26240 28224 26246
rect 28172 26182 28224 26188
rect 28184 25770 28212 26182
rect 28172 25764 28224 25770
rect 28172 25706 28224 25712
rect 28920 25498 28948 27474
rect 29000 25968 29052 25974
rect 29000 25910 29052 25916
rect 28908 25492 28960 25498
rect 28908 25434 28960 25440
rect 28632 25356 28684 25362
rect 28632 25298 28684 25304
rect 28448 25152 28500 25158
rect 28448 25094 28500 25100
rect 28264 24608 28316 24614
rect 28264 24550 28316 24556
rect 28276 24410 28304 24550
rect 28264 24404 28316 24410
rect 28264 24346 28316 24352
rect 28080 23860 28132 23866
rect 28080 23802 28132 23808
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 28356 23656 28408 23662
rect 28356 23598 28408 23604
rect 28092 23322 28120 23598
rect 28080 23316 28132 23322
rect 28080 23258 28132 23264
rect 28368 23186 28396 23598
rect 27804 23180 27856 23186
rect 27804 23122 27856 23128
rect 28356 23180 28408 23186
rect 28356 23122 28408 23128
rect 28172 23112 28224 23118
rect 28172 23054 28224 23060
rect 27712 23044 27764 23050
rect 27712 22986 27764 22992
rect 27988 23044 28040 23050
rect 27988 22986 28040 22992
rect 27620 22160 27672 22166
rect 27618 22128 27620 22137
rect 27672 22128 27674 22137
rect 27618 22063 27674 22072
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27632 20602 27660 21830
rect 27724 21128 27752 22986
rect 27896 22704 27948 22710
rect 27896 22646 27948 22652
rect 27908 22098 27936 22646
rect 28000 22420 28028 22986
rect 28184 22778 28212 23054
rect 28172 22772 28224 22778
rect 28172 22714 28224 22720
rect 28368 22710 28396 23122
rect 28356 22704 28408 22710
rect 28356 22646 28408 22652
rect 28460 22574 28488 25094
rect 28644 24818 28672 25298
rect 29012 24818 29040 25910
rect 29104 25378 29132 29718
rect 29184 28552 29236 28558
rect 29184 28494 29236 28500
rect 29196 26994 29224 28494
rect 29288 28218 29316 32914
rect 30024 31346 30052 34002
rect 30217 33756 30525 33765
rect 30217 33754 30223 33756
rect 30279 33754 30303 33756
rect 30359 33754 30383 33756
rect 30439 33754 30463 33756
rect 30519 33754 30525 33756
rect 30279 33702 30281 33754
rect 30461 33702 30463 33754
rect 30217 33700 30223 33702
rect 30279 33700 30303 33702
rect 30359 33700 30383 33702
rect 30439 33700 30463 33702
rect 30519 33700 30525 33702
rect 30217 33691 30525 33700
rect 30877 33212 31185 33221
rect 30877 33210 30883 33212
rect 30939 33210 30963 33212
rect 31019 33210 31043 33212
rect 31099 33210 31123 33212
rect 31179 33210 31185 33212
rect 30939 33158 30941 33210
rect 31121 33158 31123 33210
rect 30877 33156 30883 33158
rect 30939 33156 30963 33158
rect 31019 33156 31043 33158
rect 31099 33156 31123 33158
rect 31179 33156 31185 33158
rect 30877 33147 31185 33156
rect 30217 32668 30525 32677
rect 30217 32666 30223 32668
rect 30279 32666 30303 32668
rect 30359 32666 30383 32668
rect 30439 32666 30463 32668
rect 30519 32666 30525 32668
rect 30279 32614 30281 32666
rect 30461 32614 30463 32666
rect 30217 32612 30223 32614
rect 30279 32612 30303 32614
rect 30359 32612 30383 32614
rect 30439 32612 30463 32614
rect 30519 32612 30525 32614
rect 30217 32603 30525 32612
rect 31220 32434 31248 34002
rect 31312 33522 31340 35686
rect 32218 35678 32274 36478
rect 33506 35678 33562 36478
rect 34794 35678 34850 36478
rect 36082 35678 36138 36478
rect 31300 33516 31352 33522
rect 31300 33458 31352 33464
rect 31392 33448 31444 33454
rect 31392 33390 31444 33396
rect 30380 32428 30432 32434
rect 30380 32370 30432 32376
rect 31208 32428 31260 32434
rect 31208 32370 31260 32376
rect 30392 32026 30420 32370
rect 30877 32124 31185 32133
rect 30877 32122 30883 32124
rect 30939 32122 30963 32124
rect 31019 32122 31043 32124
rect 31099 32122 31123 32124
rect 31179 32122 31185 32124
rect 30939 32070 30941 32122
rect 31121 32070 31123 32122
rect 30877 32068 30883 32070
rect 30939 32068 30963 32070
rect 31019 32068 31043 32070
rect 31099 32068 31123 32070
rect 31179 32068 31185 32070
rect 30877 32059 31185 32068
rect 30380 32020 30432 32026
rect 30380 31962 30432 31968
rect 31300 31952 31352 31958
rect 31300 31894 31352 31900
rect 30564 31816 30616 31822
rect 30564 31758 30616 31764
rect 30217 31580 30525 31589
rect 30217 31578 30223 31580
rect 30279 31578 30303 31580
rect 30359 31578 30383 31580
rect 30439 31578 30463 31580
rect 30519 31578 30525 31580
rect 30279 31526 30281 31578
rect 30461 31526 30463 31578
rect 30217 31524 30223 31526
rect 30279 31524 30303 31526
rect 30359 31524 30383 31526
rect 30439 31524 30463 31526
rect 30519 31524 30525 31526
rect 30217 31515 30525 31524
rect 30012 31340 30064 31346
rect 30012 31282 30064 31288
rect 30196 31136 30248 31142
rect 30196 31078 30248 31084
rect 30208 30938 30236 31078
rect 30196 30932 30248 30938
rect 30196 30874 30248 30880
rect 30217 30492 30525 30501
rect 30217 30490 30223 30492
rect 30279 30490 30303 30492
rect 30359 30490 30383 30492
rect 30439 30490 30463 30492
rect 30519 30490 30525 30492
rect 30279 30438 30281 30490
rect 30461 30438 30463 30490
rect 30217 30436 30223 30438
rect 30279 30436 30303 30438
rect 30359 30436 30383 30438
rect 30439 30436 30463 30438
rect 30519 30436 30525 30438
rect 30217 30427 30525 30436
rect 30576 30274 30604 31758
rect 31312 31482 31340 31894
rect 31300 31476 31352 31482
rect 31300 31418 31352 31424
rect 30748 31272 30800 31278
rect 30748 31214 30800 31220
rect 30760 30394 30788 31214
rect 30877 31036 31185 31045
rect 30877 31034 30883 31036
rect 30939 31034 30963 31036
rect 31019 31034 31043 31036
rect 31099 31034 31123 31036
rect 31179 31034 31185 31036
rect 30939 30982 30941 31034
rect 31121 30982 31123 31034
rect 30877 30980 30883 30982
rect 30939 30980 30963 30982
rect 31019 30980 31043 30982
rect 31099 30980 31123 30982
rect 31179 30980 31185 30982
rect 30877 30971 31185 30980
rect 31404 30802 31432 33390
rect 32232 32842 32260 35678
rect 33046 34096 33102 34105
rect 33046 34031 33102 34040
rect 33060 33658 33088 34031
rect 33048 33652 33100 33658
rect 33048 33594 33100 33600
rect 32680 33380 32732 33386
rect 32680 33322 32732 33328
rect 32312 32972 32364 32978
rect 32312 32914 32364 32920
rect 32220 32836 32272 32842
rect 32220 32778 32272 32784
rect 32220 31884 32272 31890
rect 32220 31826 32272 31832
rect 31852 31816 31904 31822
rect 31852 31758 31904 31764
rect 32128 31816 32180 31822
rect 32128 31758 32180 31764
rect 31864 31226 31892 31758
rect 32140 31385 32168 31758
rect 32126 31376 32182 31385
rect 32126 31311 32182 31320
rect 31576 31204 31628 31210
rect 31864 31198 31984 31226
rect 31576 31146 31628 31152
rect 31588 30938 31616 31146
rect 31852 31136 31904 31142
rect 31852 31078 31904 31084
rect 31864 30938 31892 31078
rect 31576 30932 31628 30938
rect 31576 30874 31628 30880
rect 31852 30932 31904 30938
rect 31852 30874 31904 30880
rect 31392 30796 31444 30802
rect 31392 30738 31444 30744
rect 31588 30598 31616 30874
rect 30840 30592 30892 30598
rect 30840 30534 30892 30540
rect 31208 30592 31260 30598
rect 31208 30534 31260 30540
rect 31392 30592 31444 30598
rect 31392 30534 31444 30540
rect 31576 30592 31628 30598
rect 31576 30534 31628 30540
rect 30748 30388 30800 30394
rect 30748 30330 30800 30336
rect 30392 30246 30604 30274
rect 30852 30258 30880 30534
rect 30840 30252 30892 30258
rect 30392 30190 30420 30246
rect 30840 30194 30892 30200
rect 31220 30190 31248 30534
rect 29368 30184 29420 30190
rect 29368 30126 29420 30132
rect 30380 30184 30432 30190
rect 30380 30126 30432 30132
rect 30472 30184 30524 30190
rect 30472 30126 30524 30132
rect 30656 30184 30708 30190
rect 30656 30126 30708 30132
rect 31208 30184 31260 30190
rect 31208 30126 31260 30132
rect 29380 29306 29408 30126
rect 30392 29782 30420 30126
rect 30484 29850 30512 30126
rect 30472 29844 30524 29850
rect 30472 29786 30524 29792
rect 30380 29776 30432 29782
rect 30380 29718 30432 29724
rect 30104 29708 30156 29714
rect 30104 29650 30156 29656
rect 29368 29300 29420 29306
rect 29368 29242 29420 29248
rect 30116 29034 30144 29650
rect 30668 29510 30696 30126
rect 30877 29948 31185 29957
rect 30877 29946 30883 29948
rect 30939 29946 30963 29948
rect 31019 29946 31043 29948
rect 31099 29946 31123 29948
rect 31179 29946 31185 29948
rect 30939 29894 30941 29946
rect 31121 29894 31123 29946
rect 30877 29892 30883 29894
rect 30939 29892 30963 29894
rect 31019 29892 31043 29894
rect 31099 29892 31123 29894
rect 31179 29892 31185 29894
rect 30877 29883 31185 29892
rect 30656 29504 30708 29510
rect 30656 29446 30708 29452
rect 30217 29404 30525 29413
rect 30217 29402 30223 29404
rect 30279 29402 30303 29404
rect 30359 29402 30383 29404
rect 30439 29402 30463 29404
rect 30519 29402 30525 29404
rect 30279 29350 30281 29402
rect 30461 29350 30463 29402
rect 30217 29348 30223 29350
rect 30279 29348 30303 29350
rect 30359 29348 30383 29350
rect 30439 29348 30463 29350
rect 30519 29348 30525 29350
rect 30217 29339 30525 29348
rect 30104 29028 30156 29034
rect 30104 28970 30156 28976
rect 29368 28960 29420 28966
rect 29368 28902 29420 28908
rect 29276 28212 29328 28218
rect 29276 28154 29328 28160
rect 29380 27878 29408 28902
rect 29460 28552 29512 28558
rect 29460 28494 29512 28500
rect 29472 28218 29500 28494
rect 29460 28212 29512 28218
rect 29460 28154 29512 28160
rect 30012 28008 30064 28014
rect 30012 27950 30064 27956
rect 29368 27872 29420 27878
rect 29368 27814 29420 27820
rect 29276 27532 29328 27538
rect 29276 27474 29328 27480
rect 29288 27334 29316 27474
rect 29552 27464 29604 27470
rect 29552 27406 29604 27412
rect 29276 27328 29328 27334
rect 29328 27288 29408 27316
rect 29276 27270 29328 27276
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 29196 25906 29224 26930
rect 29276 26784 29328 26790
rect 29276 26726 29328 26732
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 29288 25770 29316 26726
rect 29380 25906 29408 27288
rect 29564 26858 29592 27406
rect 29552 26852 29604 26858
rect 29552 26794 29604 26800
rect 30024 26234 30052 27950
rect 30116 27606 30144 28970
rect 30564 28620 30616 28626
rect 30564 28562 30616 28568
rect 30217 28316 30525 28325
rect 30217 28314 30223 28316
rect 30279 28314 30303 28316
rect 30359 28314 30383 28316
rect 30439 28314 30463 28316
rect 30519 28314 30525 28316
rect 30279 28262 30281 28314
rect 30461 28262 30463 28314
rect 30217 28260 30223 28262
rect 30279 28260 30303 28262
rect 30359 28260 30383 28262
rect 30439 28260 30463 28262
rect 30519 28260 30525 28262
rect 30217 28251 30525 28260
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30104 27600 30156 27606
rect 30104 27542 30156 27548
rect 30392 27538 30420 27950
rect 30576 27674 30604 28562
rect 30668 28558 30696 29446
rect 31208 29096 31260 29102
rect 31208 29038 31260 29044
rect 30877 28860 31185 28869
rect 30877 28858 30883 28860
rect 30939 28858 30963 28860
rect 31019 28858 31043 28860
rect 31099 28858 31123 28860
rect 31179 28858 31185 28860
rect 30939 28806 30941 28858
rect 31121 28806 31123 28858
rect 30877 28804 30883 28806
rect 30939 28804 30963 28806
rect 31019 28804 31043 28806
rect 31099 28804 31123 28806
rect 31179 28804 31185 28806
rect 30877 28795 31185 28804
rect 31220 28762 31248 29038
rect 31404 28966 31432 30534
rect 31668 29776 31720 29782
rect 31668 29718 31720 29724
rect 31300 28960 31352 28966
rect 31300 28902 31352 28908
rect 31392 28960 31444 28966
rect 31392 28902 31444 28908
rect 31208 28756 31260 28762
rect 31208 28698 31260 28704
rect 31312 28694 31340 28902
rect 31300 28688 31352 28694
rect 31300 28630 31352 28636
rect 30656 28552 30708 28558
rect 30656 28494 30708 28500
rect 31024 28552 31076 28558
rect 31024 28494 31076 28500
rect 31036 28014 31064 28494
rect 31404 28082 31432 28902
rect 31680 28082 31708 29718
rect 31852 29096 31904 29102
rect 31852 29038 31904 29044
rect 31864 28218 31892 29038
rect 31852 28212 31904 28218
rect 31852 28154 31904 28160
rect 31392 28076 31444 28082
rect 31392 28018 31444 28024
rect 31668 28076 31720 28082
rect 31668 28018 31720 28024
rect 31024 28008 31076 28014
rect 31024 27950 31076 27956
rect 30656 27872 30708 27878
rect 30656 27814 30708 27820
rect 30564 27668 30616 27674
rect 30564 27610 30616 27616
rect 30380 27532 30432 27538
rect 30380 27474 30432 27480
rect 30104 27464 30156 27470
rect 30104 27406 30156 27412
rect 30564 27464 30616 27470
rect 30564 27406 30616 27412
rect 30116 26586 30144 27406
rect 30217 27228 30525 27237
rect 30217 27226 30223 27228
rect 30279 27226 30303 27228
rect 30359 27226 30383 27228
rect 30439 27226 30463 27228
rect 30519 27226 30525 27228
rect 30279 27174 30281 27226
rect 30461 27174 30463 27226
rect 30217 27172 30223 27174
rect 30279 27172 30303 27174
rect 30359 27172 30383 27174
rect 30439 27172 30463 27174
rect 30519 27172 30525 27174
rect 30217 27163 30525 27172
rect 30576 27130 30604 27406
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30668 26926 30696 27814
rect 30877 27772 31185 27781
rect 30877 27770 30883 27772
rect 30939 27770 30963 27772
rect 31019 27770 31043 27772
rect 31099 27770 31123 27772
rect 31179 27770 31185 27772
rect 30939 27718 30941 27770
rect 31121 27718 31123 27770
rect 30877 27716 30883 27718
rect 30939 27716 30963 27718
rect 31019 27716 31043 27718
rect 31099 27716 31123 27718
rect 31179 27716 31185 27718
rect 30877 27707 31185 27716
rect 31680 27674 31708 28018
rect 31668 27668 31720 27674
rect 31668 27610 31720 27616
rect 31392 27600 31444 27606
rect 31392 27542 31444 27548
rect 31404 27334 31432 27542
rect 30748 27328 30800 27334
rect 30748 27270 30800 27276
rect 31392 27328 31444 27334
rect 31392 27270 31444 27276
rect 30656 26920 30708 26926
rect 30656 26862 30708 26868
rect 30104 26580 30156 26586
rect 30104 26522 30156 26528
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30024 26206 30144 26234
rect 29368 25900 29420 25906
rect 29368 25842 29420 25848
rect 29276 25764 29328 25770
rect 29276 25706 29328 25712
rect 29104 25350 29316 25378
rect 30116 25362 30144 26206
rect 30217 26140 30525 26149
rect 30217 26138 30223 26140
rect 30279 26138 30303 26140
rect 30359 26138 30383 26140
rect 30439 26138 30463 26140
rect 30519 26138 30525 26140
rect 30279 26086 30281 26138
rect 30461 26086 30463 26138
rect 30217 26084 30223 26086
rect 30279 26084 30303 26086
rect 30359 26084 30383 26086
rect 30439 26084 30463 26086
rect 30519 26084 30525 26086
rect 30217 26075 30525 26084
rect 30576 25702 30604 26318
rect 30760 25770 30788 27270
rect 31852 26988 31904 26994
rect 31852 26930 31904 26936
rect 31484 26852 31536 26858
rect 31484 26794 31536 26800
rect 30877 26684 31185 26693
rect 30877 26682 30883 26684
rect 30939 26682 30963 26684
rect 31019 26682 31043 26684
rect 31099 26682 31123 26684
rect 31179 26682 31185 26684
rect 30939 26630 30941 26682
rect 31121 26630 31123 26682
rect 30877 26628 30883 26630
rect 30939 26628 30963 26630
rect 31019 26628 31043 26630
rect 31099 26628 31123 26630
rect 31179 26628 31185 26630
rect 30877 26619 31185 26628
rect 31496 26586 31524 26794
rect 31484 26580 31536 26586
rect 31484 26522 31536 26528
rect 30932 26376 30984 26382
rect 30932 26318 30984 26324
rect 30944 26042 30972 26318
rect 31864 26314 31892 26930
rect 31852 26308 31904 26314
rect 31852 26250 31904 26256
rect 31956 26234 31984 31198
rect 32036 31204 32088 31210
rect 32036 31146 32088 31152
rect 32048 29646 32076 31146
rect 32232 30274 32260 31826
rect 32140 30246 32260 30274
rect 32140 30054 32168 30246
rect 32220 30116 32272 30122
rect 32220 30058 32272 30064
rect 32128 30048 32180 30054
rect 32128 29990 32180 29996
rect 32036 29640 32088 29646
rect 32088 29600 32168 29628
rect 32036 29582 32088 29588
rect 32036 28960 32088 28966
rect 32036 28902 32088 28908
rect 32048 28694 32076 28902
rect 32036 28688 32088 28694
rect 32036 28630 32088 28636
rect 32036 27668 32088 27674
rect 32036 27610 32088 27616
rect 32048 27470 32076 27610
rect 32140 27470 32168 29600
rect 32232 29306 32260 30058
rect 32220 29300 32272 29306
rect 32220 29242 32272 29248
rect 32324 28506 32352 32914
rect 32404 32904 32456 32910
rect 32404 32846 32456 32852
rect 32232 28478 32352 28506
rect 32036 27464 32088 27470
rect 32036 27406 32088 27412
rect 32128 27464 32180 27470
rect 32128 27406 32180 27412
rect 32036 27328 32088 27334
rect 32036 27270 32088 27276
rect 32048 26586 32076 27270
rect 32232 26994 32260 28478
rect 32312 28416 32364 28422
rect 32312 28358 32364 28364
rect 32324 27946 32352 28358
rect 32312 27940 32364 27946
rect 32312 27882 32364 27888
rect 32416 27470 32444 32846
rect 32496 31272 32548 31278
rect 32496 31214 32548 31220
rect 32508 29850 32536 31214
rect 32496 29844 32548 29850
rect 32496 29786 32548 29792
rect 32588 29096 32640 29102
rect 32588 29038 32640 29044
rect 32600 28422 32628 29038
rect 32588 28416 32640 28422
rect 32588 28358 32640 28364
rect 32692 27946 32720 33322
rect 33048 32360 33100 32366
rect 33048 32302 33100 32308
rect 32772 31272 32824 31278
rect 32772 31214 32824 31220
rect 32784 30394 32812 31214
rect 33060 30938 33088 32302
rect 33520 31958 33548 35678
rect 33782 35456 33838 35465
rect 33782 35391 33838 35400
rect 33508 31952 33560 31958
rect 33508 31894 33560 31900
rect 33796 31346 33824 35391
rect 34808 33046 34836 35678
rect 36096 33046 36124 35678
rect 34796 33040 34848 33046
rect 34796 32982 34848 32988
rect 36084 33040 36136 33046
rect 36084 32982 36136 32988
rect 34886 32736 34942 32745
rect 34886 32671 34942 32680
rect 34900 32434 34928 32671
rect 34888 32428 34940 32434
rect 34888 32370 34940 32376
rect 33784 31340 33836 31346
rect 33784 31282 33836 31288
rect 33048 30932 33100 30938
rect 33048 30874 33100 30880
rect 32772 30388 32824 30394
rect 32772 30330 32824 30336
rect 32784 29714 32812 30330
rect 33060 29850 33088 30874
rect 35164 30184 35216 30190
rect 35164 30126 35216 30132
rect 34060 30116 34112 30122
rect 34060 30058 34112 30064
rect 33048 29844 33100 29850
rect 33048 29786 33100 29792
rect 32772 29708 32824 29714
rect 32772 29650 32824 29656
rect 33048 29708 33100 29714
rect 33048 29650 33100 29656
rect 32864 28416 32916 28422
rect 32864 28358 32916 28364
rect 32876 28082 32904 28358
rect 32864 28076 32916 28082
rect 32864 28018 32916 28024
rect 32680 27940 32732 27946
rect 32680 27882 32732 27888
rect 32692 27674 32720 27882
rect 32496 27668 32548 27674
rect 32496 27610 32548 27616
rect 32680 27668 32732 27674
rect 32680 27610 32732 27616
rect 32404 27464 32456 27470
rect 32404 27406 32456 27412
rect 32220 26988 32272 26994
rect 32220 26930 32272 26936
rect 32508 26790 32536 27610
rect 33060 27577 33088 29650
rect 33784 29028 33836 29034
rect 33784 28970 33836 28976
rect 33140 28960 33192 28966
rect 33140 28902 33192 28908
rect 33152 28626 33180 28902
rect 33796 28665 33824 28970
rect 33782 28656 33838 28665
rect 33140 28620 33192 28626
rect 33782 28591 33838 28600
rect 33140 28562 33192 28568
rect 33046 27568 33102 27577
rect 33046 27503 33102 27512
rect 33048 27464 33100 27470
rect 33048 27406 33100 27412
rect 32588 27396 32640 27402
rect 32588 27338 32640 27344
rect 32600 27130 32628 27338
rect 33060 27130 33088 27406
rect 32588 27124 32640 27130
rect 32588 27066 32640 27072
rect 33048 27124 33100 27130
rect 33048 27066 33100 27072
rect 33060 27010 33088 27066
rect 33152 27062 33180 28562
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33428 27470 33456 28494
rect 33876 28416 33928 28422
rect 33876 28358 33928 28364
rect 33888 28014 33916 28358
rect 33876 28008 33928 28014
rect 33876 27950 33928 27956
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 33784 27328 33836 27334
rect 33784 27270 33836 27276
rect 32692 26982 33088 27010
rect 33140 27056 33192 27062
rect 33140 26998 33192 27004
rect 32496 26784 32548 26790
rect 32496 26726 32548 26732
rect 32036 26580 32088 26586
rect 32036 26522 32088 26528
rect 31956 26206 32352 26234
rect 30932 26036 30984 26042
rect 30932 25978 30984 25984
rect 30748 25764 30800 25770
rect 30748 25706 30800 25712
rect 30564 25696 30616 25702
rect 30564 25638 30616 25644
rect 30877 25596 31185 25605
rect 30877 25594 30883 25596
rect 30939 25594 30963 25596
rect 31019 25594 31043 25596
rect 31099 25594 31123 25596
rect 31179 25594 31185 25596
rect 30939 25542 30941 25594
rect 31121 25542 31123 25594
rect 30877 25540 30883 25542
rect 30939 25540 30963 25542
rect 31019 25540 31043 25542
rect 31099 25540 31123 25542
rect 31179 25540 31185 25542
rect 30877 25531 31185 25540
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 29000 24812 29052 24818
rect 29000 24754 29052 24760
rect 28816 24744 28868 24750
rect 28816 24686 28868 24692
rect 28540 24676 28592 24682
rect 28540 24618 28592 24624
rect 28552 24274 28580 24618
rect 28724 24336 28776 24342
rect 28724 24278 28776 24284
rect 28540 24268 28592 24274
rect 28540 24210 28592 24216
rect 28736 24177 28764 24278
rect 28722 24168 28778 24177
rect 28722 24103 28778 24112
rect 28724 24064 28776 24070
rect 28724 24006 28776 24012
rect 28540 23520 28592 23526
rect 28540 23462 28592 23468
rect 28448 22568 28500 22574
rect 28448 22510 28500 22516
rect 28172 22432 28224 22438
rect 28000 22392 28172 22420
rect 28172 22374 28224 22380
rect 28448 22432 28500 22438
rect 28552 22420 28580 23462
rect 28736 23186 28764 24006
rect 28828 23866 28856 24686
rect 29184 24200 29236 24206
rect 29184 24142 29236 24148
rect 28816 23860 28868 23866
rect 28816 23802 28868 23808
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 28920 23526 28948 23802
rect 28908 23520 28960 23526
rect 28908 23462 28960 23468
rect 28724 23180 28776 23186
rect 28724 23122 28776 23128
rect 29092 23180 29144 23186
rect 29092 23122 29144 23128
rect 28500 22392 28580 22420
rect 28448 22374 28500 22380
rect 27986 22128 28042 22137
rect 27896 22092 27948 22098
rect 27986 22063 28042 22072
rect 27896 22034 27948 22040
rect 28000 22012 28028 22063
rect 28080 22024 28132 22030
rect 28000 21984 28080 22012
rect 28080 21966 28132 21972
rect 28184 21894 28212 22374
rect 28172 21888 28224 21894
rect 28172 21830 28224 21836
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 27988 21140 28040 21146
rect 27724 21100 27844 21128
rect 27816 21010 27844 21100
rect 27988 21082 28040 21088
rect 27712 21004 27764 21010
rect 27712 20946 27764 20952
rect 27804 21004 27856 21010
rect 27804 20946 27856 20952
rect 27724 20602 27752 20946
rect 28000 20890 28028 21082
rect 28184 21078 28212 21422
rect 28460 21146 28488 22374
rect 29104 22098 29132 23122
rect 29196 22642 29224 24142
rect 29184 22636 29236 22642
rect 29184 22578 29236 22584
rect 29288 22166 29316 25350
rect 30104 25356 30156 25362
rect 30104 25298 30156 25304
rect 29828 25288 29880 25294
rect 29828 25230 29880 25236
rect 29368 25152 29420 25158
rect 29368 25094 29420 25100
rect 29380 24818 29408 25094
rect 29368 24812 29420 24818
rect 29368 24754 29420 24760
rect 29840 24410 29868 25230
rect 29828 24404 29880 24410
rect 29828 24346 29880 24352
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 29644 24268 29696 24274
rect 29644 24210 29696 24216
rect 29828 24268 29880 24274
rect 29828 24210 29880 24216
rect 29564 23866 29592 24210
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 29656 23798 29684 24210
rect 29644 23792 29696 23798
rect 29644 23734 29696 23740
rect 29656 22982 29684 23734
rect 29840 23186 29868 24210
rect 29920 24064 29972 24070
rect 29920 24006 29972 24012
rect 29932 23594 29960 24006
rect 29920 23588 29972 23594
rect 29920 23530 29972 23536
rect 29828 23180 29880 23186
rect 29828 23122 29880 23128
rect 29644 22976 29696 22982
rect 29644 22918 29696 22924
rect 29828 22976 29880 22982
rect 29828 22918 29880 22924
rect 29552 22500 29604 22506
rect 29552 22442 29604 22448
rect 29276 22160 29328 22166
rect 29276 22102 29328 22108
rect 29092 22092 29144 22098
rect 29092 22034 29144 22040
rect 29000 21888 29052 21894
rect 29000 21830 29052 21836
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 28172 21072 28224 21078
rect 28172 21014 28224 21020
rect 28356 21072 28408 21078
rect 28356 21014 28408 21020
rect 27816 20862 28028 20890
rect 27620 20596 27672 20602
rect 27620 20538 27672 20544
rect 27712 20596 27764 20602
rect 27712 20538 27764 20544
rect 27528 20392 27580 20398
rect 27528 20334 27580 20340
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27436 20324 27488 20330
rect 27436 20266 27488 20272
rect 27448 20058 27476 20266
rect 27436 20052 27488 20058
rect 27436 19994 27488 20000
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27540 19718 27568 20334
rect 27528 19712 27580 19718
rect 27528 19654 27580 19660
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27252 19236 27304 19242
rect 27252 19178 27304 19184
rect 26884 18080 26936 18086
rect 26884 18022 26936 18028
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 26896 17882 26924 18022
rect 26884 17876 26936 17882
rect 26884 17818 26936 17824
rect 26608 17332 26660 17338
rect 26608 17274 26660 17280
rect 26988 17270 27016 18022
rect 26976 17264 27028 17270
rect 26974 17232 26976 17241
rect 27028 17232 27030 17241
rect 26974 17167 27030 17176
rect 26332 16652 26384 16658
rect 26332 16594 26384 16600
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26608 16652 26660 16658
rect 26608 16594 26660 16600
rect 26332 16516 26384 16522
rect 26332 16458 26384 16464
rect 26344 15978 26372 16458
rect 26332 15972 26384 15978
rect 26332 15914 26384 15920
rect 26436 14618 26464 16594
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26424 14476 26476 14482
rect 26424 14418 26476 14424
rect 26436 14278 26464 14418
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26238 13696 26294 13705
rect 26238 13631 26294 13640
rect 26148 13456 26200 13462
rect 26148 13398 26200 13404
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26240 13388 26292 13394
rect 26240 13330 26292 13336
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 25688 13320 25740 13326
rect 25688 13262 25740 13268
rect 25700 12986 25728 13262
rect 25688 12980 25740 12986
rect 25688 12922 25740 12928
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 25320 12232 25372 12238
rect 25320 12174 25372 12180
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 24964 11694 24992 12174
rect 24952 11688 25004 11694
rect 24952 11630 25004 11636
rect 24860 11144 24912 11150
rect 24860 11086 24912 11092
rect 24872 9994 24900 11086
rect 25332 10810 25360 12174
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 25056 10266 25084 10406
rect 25044 10260 25096 10266
rect 25044 10202 25096 10208
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 25136 9920 25188 9926
rect 25136 9862 25188 9868
rect 25148 9722 25176 9862
rect 25136 9716 25188 9722
rect 25136 9658 25188 9664
rect 25516 9654 25544 12174
rect 26068 11830 26096 13330
rect 26252 12850 26280 13330
rect 26240 12844 26292 12850
rect 26240 12786 26292 12792
rect 26148 12776 26200 12782
rect 26148 12718 26200 12724
rect 26056 11824 26108 11830
rect 26056 11766 26108 11772
rect 26160 11626 26188 12718
rect 26252 12238 26280 12786
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 26148 11620 26200 11626
rect 26148 11562 26200 11568
rect 26252 11150 26280 12174
rect 26344 11354 26372 13330
rect 26436 12442 26464 13806
rect 26528 13530 26556 16594
rect 26620 15434 26648 16594
rect 26700 16040 26752 16046
rect 26700 15982 26752 15988
rect 26712 15638 26740 15982
rect 26700 15632 26752 15638
rect 26700 15574 26752 15580
rect 26608 15428 26660 15434
rect 26608 15370 26660 15376
rect 26976 15428 27028 15434
rect 26976 15370 27028 15376
rect 26700 14952 26752 14958
rect 26700 14894 26752 14900
rect 26712 14618 26740 14894
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26608 14000 26660 14006
rect 26608 13942 26660 13948
rect 26620 13870 26648 13942
rect 26712 13870 26740 14418
rect 26884 14340 26936 14346
rect 26884 14282 26936 14288
rect 26792 14272 26844 14278
rect 26792 14214 26844 14220
rect 26804 13870 26832 14214
rect 26896 14074 26924 14282
rect 26884 14068 26936 14074
rect 26884 14010 26936 14016
rect 26608 13864 26660 13870
rect 26608 13806 26660 13812
rect 26700 13864 26752 13870
rect 26700 13806 26752 13812
rect 26792 13864 26844 13870
rect 26792 13806 26844 13812
rect 26516 13524 26568 13530
rect 26516 13466 26568 13472
rect 26528 12714 26556 13466
rect 26620 13326 26648 13806
rect 26608 13320 26660 13326
rect 26608 13262 26660 13268
rect 26516 12708 26568 12714
rect 26516 12650 26568 12656
rect 26712 12442 26740 13806
rect 26896 12730 26924 14010
rect 26988 13410 27016 15370
rect 27160 15360 27212 15366
rect 27264 15348 27292 19178
rect 27356 18834 27384 19314
rect 27436 19168 27488 19174
rect 27436 19110 27488 19116
rect 27344 18828 27396 18834
rect 27344 18770 27396 18776
rect 27448 18630 27476 19110
rect 27436 18624 27488 18630
rect 27436 18566 27488 18572
rect 27448 18222 27476 18566
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27540 16658 27568 18294
rect 27632 17746 27660 20334
rect 27816 19174 27844 20862
rect 28368 20806 28396 21014
rect 27988 20800 28040 20806
rect 27988 20742 28040 20748
rect 28356 20800 28408 20806
rect 28356 20742 28408 20748
rect 27896 19916 27948 19922
rect 27896 19858 27948 19864
rect 27908 19378 27936 19858
rect 28000 19718 28028 20742
rect 29012 19854 29040 21830
rect 29288 21690 29316 22102
rect 29564 22098 29592 22442
rect 29552 22092 29604 22098
rect 29840 22094 29868 22918
rect 29552 22034 29604 22040
rect 29656 22066 29868 22094
rect 29276 21684 29328 21690
rect 29276 21626 29328 21632
rect 29656 21554 29684 22066
rect 29644 21548 29696 21554
rect 29644 21490 29696 21496
rect 29828 21480 29880 21486
rect 29828 21422 29880 21428
rect 29460 21344 29512 21350
rect 29460 21286 29512 21292
rect 29368 21072 29420 21078
rect 29368 21014 29420 21020
rect 29380 20466 29408 21014
rect 29472 20602 29500 21286
rect 29552 21140 29604 21146
rect 29552 21082 29604 21088
rect 29460 20596 29512 20602
rect 29460 20538 29512 20544
rect 29368 20460 29420 20466
rect 29368 20402 29420 20408
rect 29380 20074 29408 20402
rect 29380 20046 29500 20074
rect 29368 19984 29420 19990
rect 29368 19926 29420 19932
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 29000 19848 29052 19854
rect 29000 19790 29052 19796
rect 27988 19712 28040 19718
rect 27988 19654 28040 19660
rect 28092 19446 28120 19790
rect 29000 19712 29052 19718
rect 29000 19654 29052 19660
rect 28080 19440 28132 19446
rect 27986 19408 28042 19417
rect 27896 19372 27948 19378
rect 28080 19382 28132 19388
rect 28816 19440 28868 19446
rect 28816 19382 28868 19388
rect 27986 19343 28042 19352
rect 27896 19314 27948 19320
rect 27908 19174 27936 19314
rect 27712 19168 27764 19174
rect 27712 19110 27764 19116
rect 27804 19168 27856 19174
rect 27804 19110 27856 19116
rect 27896 19168 27948 19174
rect 27896 19110 27948 19116
rect 27724 18902 27752 19110
rect 27712 18896 27764 18902
rect 27712 18838 27764 18844
rect 27816 18426 27844 19110
rect 27908 18698 27936 19110
rect 28000 18970 28028 19343
rect 28264 19304 28316 19310
rect 28264 19246 28316 19252
rect 27988 18964 28040 18970
rect 27988 18906 28040 18912
rect 27896 18692 27948 18698
rect 27896 18634 27948 18640
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 27804 18420 27856 18426
rect 27804 18362 27856 18368
rect 27620 17740 27672 17746
rect 27620 17682 27672 17688
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27632 16998 27660 17478
rect 27620 16992 27672 16998
rect 27620 16934 27672 16940
rect 27632 16658 27660 16934
rect 27816 16674 27844 18362
rect 28080 18352 28132 18358
rect 28000 18312 28080 18340
rect 28000 18154 28028 18312
rect 28080 18294 28132 18300
rect 27988 18148 28040 18154
rect 27988 18090 28040 18096
rect 27724 16658 27844 16674
rect 27528 16652 27580 16658
rect 27528 16594 27580 16600
rect 27620 16652 27672 16658
rect 27620 16594 27672 16600
rect 27712 16652 27844 16658
rect 27764 16646 27844 16652
rect 27712 16594 27764 16600
rect 27540 16538 27568 16594
rect 27448 16510 27568 16538
rect 27344 16040 27396 16046
rect 27344 15982 27396 15988
rect 27356 15706 27384 15982
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27448 15570 27476 16510
rect 27436 15564 27488 15570
rect 27436 15506 27488 15512
rect 27212 15320 27292 15348
rect 27160 15302 27212 15308
rect 27068 14408 27120 14414
rect 27068 14350 27120 14356
rect 27080 14074 27108 14350
rect 27068 14068 27120 14074
rect 27068 14010 27120 14016
rect 27068 13864 27120 13870
rect 27172 13852 27200 15302
rect 27632 15178 27660 16594
rect 27896 16516 27948 16522
rect 27896 16458 27948 16464
rect 27908 15502 27936 16458
rect 28000 15638 28028 18090
rect 28078 17912 28134 17921
rect 28078 17847 28134 17856
rect 28092 17814 28120 17847
rect 28080 17808 28132 17814
rect 28080 17750 28132 17756
rect 28184 16794 28212 18566
rect 28276 17882 28304 19246
rect 28828 18902 28856 19382
rect 28908 18964 28960 18970
rect 28908 18906 28960 18912
rect 28448 18896 28500 18902
rect 28448 18838 28500 18844
rect 28816 18896 28868 18902
rect 28816 18838 28868 18844
rect 28356 18420 28408 18426
rect 28356 18362 28408 18368
rect 28264 17876 28316 17882
rect 28264 17818 28316 17824
rect 28262 17776 28318 17785
rect 28262 17711 28264 17720
rect 28316 17711 28318 17720
rect 28264 17682 28316 17688
rect 28368 16794 28396 18362
rect 28460 18222 28488 18838
rect 28816 18624 28868 18630
rect 28816 18566 28868 18572
rect 28448 18216 28500 18222
rect 28448 18158 28500 18164
rect 28828 18086 28856 18566
rect 28920 18290 28948 18906
rect 29012 18834 29040 19654
rect 29184 19508 29236 19514
rect 29184 19450 29236 19456
rect 29196 19357 29224 19450
rect 29182 19348 29238 19357
rect 29380 19334 29408 19926
rect 29472 19446 29500 20046
rect 29460 19440 29512 19446
rect 29460 19382 29512 19388
rect 29380 19306 29500 19334
rect 29182 19283 29238 19292
rect 29092 19168 29144 19174
rect 29276 19168 29328 19174
rect 29144 19145 29224 19156
rect 29144 19136 29238 19145
rect 29144 19128 29182 19136
rect 29092 19110 29144 19116
rect 29276 19110 29328 19116
rect 29368 19168 29420 19174
rect 29368 19110 29420 19116
rect 29182 19071 29238 19080
rect 29000 18828 29052 18834
rect 29000 18770 29052 18776
rect 29288 18426 29316 19110
rect 29380 19009 29408 19110
rect 29366 19000 29422 19009
rect 29472 18970 29500 19306
rect 29564 19174 29592 21082
rect 29840 20602 29868 21422
rect 29932 21078 29960 23530
rect 30116 23322 30144 25298
rect 30564 25152 30616 25158
rect 30564 25094 30616 25100
rect 30217 25052 30525 25061
rect 30217 25050 30223 25052
rect 30279 25050 30303 25052
rect 30359 25050 30383 25052
rect 30439 25050 30463 25052
rect 30519 25050 30525 25052
rect 30279 24998 30281 25050
rect 30461 24998 30463 25050
rect 30217 24996 30223 24998
rect 30279 24996 30303 24998
rect 30359 24996 30383 24998
rect 30439 24996 30463 24998
rect 30519 24996 30525 24998
rect 30217 24987 30525 24996
rect 30576 24750 30604 25094
rect 30564 24744 30616 24750
rect 30564 24686 30616 24692
rect 30564 24608 30616 24614
rect 30564 24550 30616 24556
rect 30576 24274 30604 24550
rect 30877 24508 31185 24517
rect 30877 24506 30883 24508
rect 30939 24506 30963 24508
rect 31019 24506 31043 24508
rect 31099 24506 31123 24508
rect 31179 24506 31185 24508
rect 30939 24454 30941 24506
rect 31121 24454 31123 24506
rect 30877 24452 30883 24454
rect 30939 24452 30963 24454
rect 31019 24452 31043 24454
rect 31099 24452 31123 24454
rect 31179 24452 31185 24454
rect 30877 24443 31185 24452
rect 30564 24268 30616 24274
rect 30564 24210 30616 24216
rect 30217 23964 30525 23973
rect 30217 23962 30223 23964
rect 30279 23962 30303 23964
rect 30359 23962 30383 23964
rect 30439 23962 30463 23964
rect 30519 23962 30525 23964
rect 30279 23910 30281 23962
rect 30461 23910 30463 23962
rect 30217 23908 30223 23910
rect 30279 23908 30303 23910
rect 30359 23908 30383 23910
rect 30439 23908 30463 23910
rect 30519 23908 30525 23910
rect 30217 23899 30525 23908
rect 30104 23316 30156 23322
rect 30104 23258 30156 23264
rect 30012 23112 30064 23118
rect 30012 23054 30064 23060
rect 29920 21072 29972 21078
rect 29920 21014 29972 21020
rect 29828 20596 29880 20602
rect 29656 20556 29828 20584
rect 29656 20398 29684 20556
rect 29828 20538 29880 20544
rect 29644 20392 29696 20398
rect 29644 20334 29696 20340
rect 29656 19990 29684 20334
rect 29920 20324 29972 20330
rect 30024 20312 30052 23054
rect 30104 22976 30156 22982
rect 30104 22918 30156 22924
rect 30116 22506 30144 22918
rect 30217 22876 30525 22885
rect 30217 22874 30223 22876
rect 30279 22874 30303 22876
rect 30359 22874 30383 22876
rect 30439 22874 30463 22876
rect 30519 22874 30525 22876
rect 30279 22822 30281 22874
rect 30461 22822 30463 22874
rect 30217 22820 30223 22822
rect 30279 22820 30303 22822
rect 30359 22820 30383 22822
rect 30439 22820 30463 22822
rect 30519 22820 30525 22822
rect 30217 22811 30525 22820
rect 30104 22500 30156 22506
rect 30104 22442 30156 22448
rect 30104 22024 30156 22030
rect 30104 21966 30156 21972
rect 30116 21690 30144 21966
rect 30576 21894 30604 24210
rect 30877 23420 31185 23429
rect 30877 23418 30883 23420
rect 30939 23418 30963 23420
rect 31019 23418 31043 23420
rect 31099 23418 31123 23420
rect 31179 23418 31185 23420
rect 30939 23366 30941 23418
rect 31121 23366 31123 23418
rect 30877 23364 30883 23366
rect 30939 23364 30963 23366
rect 31019 23364 31043 23366
rect 31099 23364 31123 23366
rect 31179 23364 31185 23366
rect 30877 23355 31185 23364
rect 31116 23180 31168 23186
rect 31116 23122 31168 23128
rect 31760 23180 31812 23186
rect 31760 23122 31812 23128
rect 30932 22976 30984 22982
rect 30932 22918 30984 22924
rect 30944 22522 30972 22918
rect 31128 22778 31156 23122
rect 31772 22778 31800 23122
rect 31116 22772 31168 22778
rect 31116 22714 31168 22720
rect 31208 22772 31260 22778
rect 31208 22714 31260 22720
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 30760 22494 30972 22522
rect 30656 22160 30708 22166
rect 30656 22102 30708 22108
rect 30564 21888 30616 21894
rect 30564 21830 30616 21836
rect 30217 21788 30525 21797
rect 30217 21786 30223 21788
rect 30279 21786 30303 21788
rect 30359 21786 30383 21788
rect 30439 21786 30463 21788
rect 30519 21786 30525 21788
rect 30279 21734 30281 21786
rect 30461 21734 30463 21786
rect 30217 21732 30223 21734
rect 30279 21732 30303 21734
rect 30359 21732 30383 21734
rect 30439 21732 30463 21734
rect 30519 21732 30525 21734
rect 30217 21723 30525 21732
rect 30668 21706 30696 22102
rect 30104 21684 30156 21690
rect 30576 21678 30696 21706
rect 30576 21672 30604 21678
rect 30104 21626 30156 21632
rect 30484 21644 30604 21672
rect 30484 20942 30512 21644
rect 30656 21480 30708 21486
rect 30760 21434 30788 22494
rect 30877 22332 31185 22341
rect 30877 22330 30883 22332
rect 30939 22330 30963 22332
rect 31019 22330 31043 22332
rect 31099 22330 31123 22332
rect 31179 22330 31185 22332
rect 30939 22278 30941 22330
rect 31121 22278 31123 22330
rect 30877 22276 30883 22278
rect 30939 22276 30963 22278
rect 31019 22276 31043 22278
rect 31099 22276 31123 22278
rect 31179 22276 31185 22278
rect 30877 22267 31185 22276
rect 30708 21428 30788 21434
rect 30656 21422 30788 21428
rect 31116 21480 31168 21486
rect 31220 21468 31248 22714
rect 31576 22636 31628 22642
rect 31576 22578 31628 22584
rect 31588 22234 31616 22578
rect 31576 22228 31628 22234
rect 31576 22170 31628 22176
rect 31588 22094 31616 22170
rect 31944 22160 31996 22166
rect 31944 22102 31996 22108
rect 31168 21440 31248 21468
rect 31116 21422 31168 21428
rect 30668 21406 30788 21422
rect 30668 21078 30696 21406
rect 30877 21244 31185 21253
rect 30877 21242 30883 21244
rect 30939 21242 30963 21244
rect 31019 21242 31043 21244
rect 31099 21242 31123 21244
rect 31179 21242 31185 21244
rect 30939 21190 30941 21242
rect 31121 21190 31123 21242
rect 30877 21188 30883 21190
rect 30939 21188 30963 21190
rect 31019 21188 31043 21190
rect 31099 21188 31123 21190
rect 31179 21188 31185 21190
rect 30877 21179 31185 21188
rect 30656 21072 30708 21078
rect 30656 21014 30708 21020
rect 30472 20936 30524 20942
rect 30472 20878 30524 20884
rect 30656 20936 30708 20942
rect 30656 20878 30708 20884
rect 31024 20936 31076 20942
rect 31024 20878 31076 20884
rect 30217 20700 30525 20709
rect 30217 20698 30223 20700
rect 30279 20698 30303 20700
rect 30359 20698 30383 20700
rect 30439 20698 30463 20700
rect 30519 20698 30525 20700
rect 30279 20646 30281 20698
rect 30461 20646 30463 20698
rect 30217 20644 30223 20646
rect 30279 20644 30303 20646
rect 30359 20644 30383 20646
rect 30439 20644 30463 20646
rect 30519 20644 30525 20646
rect 30217 20635 30525 20644
rect 30668 20398 30696 20878
rect 30932 20800 30984 20806
rect 30932 20742 30984 20748
rect 30944 20466 30972 20742
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 31036 20398 31064 20878
rect 31220 20806 31248 21440
rect 31404 22066 31616 22094
rect 31300 21412 31352 21418
rect 31300 21354 31352 21360
rect 31312 21146 31340 21354
rect 31300 21140 31352 21146
rect 31300 21082 31352 21088
rect 31208 20800 31260 20806
rect 31208 20742 31260 20748
rect 31404 20398 31432 22066
rect 31956 21690 31984 22102
rect 32324 22094 32352 26206
rect 32508 25702 32536 26726
rect 32496 25696 32548 25702
rect 32496 25638 32548 25644
rect 32232 22066 32352 22094
rect 31944 21684 31996 21690
rect 31944 21626 31996 21632
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 31772 20602 31800 20878
rect 32036 20800 32088 20806
rect 32036 20742 32088 20748
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 31484 20528 31536 20534
rect 31536 20488 31616 20516
rect 31484 20470 31536 20476
rect 30656 20392 30708 20398
rect 30656 20334 30708 20340
rect 30840 20392 30892 20398
rect 30840 20334 30892 20340
rect 31024 20392 31076 20398
rect 31024 20334 31076 20340
rect 31392 20392 31444 20398
rect 31392 20334 31444 20340
rect 29972 20284 30052 20312
rect 29920 20266 29972 20272
rect 29828 20256 29880 20262
rect 29828 20198 29880 20204
rect 30104 20256 30156 20262
rect 30104 20198 30156 20204
rect 30564 20256 30616 20262
rect 30564 20198 30616 20204
rect 29644 19984 29696 19990
rect 29840 19961 29868 20198
rect 29644 19926 29696 19932
rect 29826 19952 29882 19961
rect 29736 19916 29788 19922
rect 29826 19887 29882 19896
rect 29736 19858 29788 19864
rect 29644 19780 29696 19786
rect 29644 19722 29696 19728
rect 29552 19168 29604 19174
rect 29552 19110 29604 19116
rect 29564 18970 29592 19110
rect 29366 18935 29422 18944
rect 29460 18964 29512 18970
rect 29460 18906 29512 18912
rect 29552 18964 29604 18970
rect 29552 18906 29604 18912
rect 29276 18420 29328 18426
rect 29276 18362 29328 18368
rect 29368 18352 29420 18358
rect 29368 18294 29420 18300
rect 28908 18284 28960 18290
rect 28908 18226 28960 18232
rect 29380 18154 29408 18294
rect 29564 18154 29592 18906
rect 29656 18902 29684 19722
rect 29644 18896 29696 18902
rect 29644 18838 29696 18844
rect 29644 18760 29696 18766
rect 29644 18702 29696 18708
rect 29656 18222 29684 18702
rect 29644 18216 29696 18222
rect 29644 18158 29696 18164
rect 29368 18148 29420 18154
rect 29368 18090 29420 18096
rect 29552 18148 29604 18154
rect 29552 18090 29604 18096
rect 28448 18080 28500 18086
rect 28448 18022 28500 18028
rect 28724 18080 28776 18086
rect 28724 18022 28776 18028
rect 28816 18080 28868 18086
rect 28816 18022 28868 18028
rect 28172 16788 28224 16794
rect 28172 16730 28224 16736
rect 28356 16788 28408 16794
rect 28356 16730 28408 16736
rect 28460 16182 28488 18022
rect 28736 17921 28764 18022
rect 28722 17912 28778 17921
rect 28722 17847 28778 17856
rect 28828 17785 28856 18022
rect 29380 17882 29408 18090
rect 29460 18080 29512 18086
rect 29460 18022 29512 18028
rect 29368 17876 29420 17882
rect 29368 17818 29420 17824
rect 28814 17776 28870 17785
rect 28540 17740 28592 17746
rect 28814 17711 28870 17720
rect 29368 17740 29420 17746
rect 28540 17682 28592 17688
rect 28552 17542 28580 17682
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28632 17536 28684 17542
rect 28632 17478 28684 17484
rect 28552 16590 28580 17478
rect 28644 17202 28672 17478
rect 28632 17196 28684 17202
rect 28632 17138 28684 17144
rect 28724 16652 28776 16658
rect 28724 16594 28776 16600
rect 28540 16584 28592 16590
rect 28540 16526 28592 16532
rect 28736 16454 28764 16594
rect 28724 16448 28776 16454
rect 28724 16390 28776 16396
rect 28448 16176 28500 16182
rect 28448 16118 28500 16124
rect 28736 16046 28764 16390
rect 28828 16046 28856 17711
rect 29368 17682 29420 17688
rect 29184 17672 29236 17678
rect 29184 17614 29236 17620
rect 28908 17604 28960 17610
rect 28908 17546 28960 17552
rect 28920 16998 28948 17546
rect 29000 17060 29052 17066
rect 29000 17002 29052 17008
rect 28908 16992 28960 16998
rect 28908 16934 28960 16940
rect 28920 16250 28948 16934
rect 28908 16244 28960 16250
rect 28908 16186 28960 16192
rect 28724 16040 28776 16046
rect 28724 15982 28776 15988
rect 28816 16040 28868 16046
rect 28816 15982 28868 15988
rect 27988 15632 28040 15638
rect 27988 15574 28040 15580
rect 28632 15564 28684 15570
rect 28632 15506 28684 15512
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 28080 15360 28132 15366
rect 28080 15302 28132 15308
rect 27540 15162 27660 15178
rect 27528 15156 27660 15162
rect 27580 15150 27660 15156
rect 27528 15098 27580 15104
rect 27344 14884 27396 14890
rect 27344 14826 27396 14832
rect 27356 14618 27384 14826
rect 27344 14612 27396 14618
rect 27344 14554 27396 14560
rect 27632 14074 27660 15150
rect 28092 14890 28120 15302
rect 28644 14890 28672 15506
rect 28736 15026 28764 15982
rect 28816 15904 28868 15910
rect 28816 15846 28868 15852
rect 28724 15020 28776 15026
rect 28724 14962 28776 14968
rect 28080 14884 28132 14890
rect 28080 14826 28132 14832
rect 28632 14884 28684 14890
rect 28632 14826 28684 14832
rect 27988 14544 28040 14550
rect 27988 14486 28040 14492
rect 27620 14068 27672 14074
rect 27620 14010 27672 14016
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27120 13824 27200 13852
rect 27068 13806 27120 13812
rect 27436 13796 27488 13802
rect 27436 13738 27488 13744
rect 27448 13530 27476 13738
rect 27436 13524 27488 13530
rect 27436 13466 27488 13472
rect 26988 13394 27108 13410
rect 26988 13388 27120 13394
rect 26988 13382 27068 13388
rect 27068 13330 27120 13336
rect 26976 13252 27028 13258
rect 26976 13194 27028 13200
rect 26804 12702 26924 12730
rect 26424 12436 26476 12442
rect 26424 12378 26476 12384
rect 26700 12436 26752 12442
rect 26700 12378 26752 12384
rect 26804 12322 26832 12702
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 26424 12300 26476 12306
rect 26424 12242 26476 12248
rect 26620 12294 26832 12322
rect 26896 12322 26924 12582
rect 26988 12434 27016 13194
rect 27080 12782 27108 13330
rect 27068 12776 27120 12782
rect 27068 12718 27120 12724
rect 27540 12714 27568 13874
rect 27712 13728 27764 13734
rect 27712 13670 27764 13676
rect 27724 12986 27752 13670
rect 27896 13388 27948 13394
rect 27896 13330 27948 13336
rect 27712 12980 27764 12986
rect 27712 12922 27764 12928
rect 27528 12708 27580 12714
rect 27528 12650 27580 12656
rect 27908 12442 27936 13330
rect 28000 12782 28028 14486
rect 28644 14482 28672 14826
rect 28632 14476 28684 14482
rect 28552 14436 28632 14464
rect 28356 13388 28408 13394
rect 28356 13330 28408 13336
rect 28368 12850 28396 13330
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 27988 12776 28040 12782
rect 27988 12718 28040 12724
rect 28080 12708 28132 12714
rect 28080 12650 28132 12656
rect 27896 12436 27948 12442
rect 26988 12406 27108 12434
rect 26896 12306 27016 12322
rect 26896 12300 27028 12306
rect 26896 12294 26976 12300
rect 26436 11830 26464 12242
rect 26424 11824 26476 11830
rect 26424 11766 26476 11772
rect 26620 11694 26648 12294
rect 26976 12242 27028 12248
rect 27080 12238 27108 12406
rect 27896 12378 27948 12384
rect 27068 12232 27120 12238
rect 27068 12174 27120 12180
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 27080 11898 27108 12038
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 27804 11756 27856 11762
rect 27804 11698 27856 11704
rect 26608 11688 26660 11694
rect 26608 11630 26660 11636
rect 26332 11348 26384 11354
rect 26332 11290 26384 11296
rect 27816 11286 27844 11698
rect 27804 11280 27856 11286
rect 27804 11222 27856 11228
rect 26240 11144 26292 11150
rect 26240 11086 26292 11092
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26976 11144 27028 11150
rect 26976 11086 27028 11092
rect 25964 10532 26016 10538
rect 25964 10474 26016 10480
rect 25976 10266 26004 10474
rect 25964 10260 26016 10266
rect 25964 10202 26016 10208
rect 26436 10198 26464 11086
rect 26988 10810 27016 11086
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 26976 10804 27028 10810
rect 26976 10746 27028 10752
rect 27356 10266 27384 10950
rect 27816 10606 27844 11222
rect 28092 10810 28120 12650
rect 28262 11792 28318 11801
rect 28262 11727 28264 11736
rect 28316 11727 28318 11736
rect 28264 11698 28316 11704
rect 28172 11688 28224 11694
rect 28172 11630 28224 11636
rect 28184 11354 28212 11630
rect 28172 11348 28224 11354
rect 28172 11290 28224 11296
rect 28552 11218 28580 14436
rect 28828 14464 28856 15846
rect 29012 15638 29040 17002
rect 29196 16590 29224 17614
rect 29184 16584 29236 16590
rect 29184 16526 29236 16532
rect 29380 15910 29408 17682
rect 29472 17542 29500 18022
rect 29656 17678 29684 18158
rect 29644 17672 29696 17678
rect 29644 17614 29696 17620
rect 29460 17536 29512 17542
rect 29460 17478 29512 17484
rect 29552 17536 29604 17542
rect 29552 17478 29604 17484
rect 29472 16998 29500 17478
rect 29460 16992 29512 16998
rect 29460 16934 29512 16940
rect 29564 16794 29592 17478
rect 29656 17338 29684 17614
rect 29644 17332 29696 17338
rect 29644 17274 29696 17280
rect 29552 16788 29604 16794
rect 29552 16730 29604 16736
rect 29656 16674 29684 17274
rect 29748 17134 29776 19858
rect 30116 19514 30144 20198
rect 30576 19922 30604 20198
rect 30564 19916 30616 19922
rect 30564 19858 30616 19864
rect 30668 19802 30696 20334
rect 30748 20256 30800 20262
rect 30852 20244 30880 20334
rect 31588 20330 31616 20488
rect 32048 20398 32076 20742
rect 32036 20392 32088 20398
rect 32036 20334 32088 20340
rect 31576 20324 31628 20330
rect 31576 20266 31628 20272
rect 31024 20256 31076 20262
rect 30852 20216 31024 20244
rect 30748 20198 30800 20204
rect 31024 20198 31076 20204
rect 30760 20058 30788 20198
rect 30877 20156 31185 20165
rect 30877 20154 30883 20156
rect 30939 20154 30963 20156
rect 31019 20154 31043 20156
rect 31099 20154 31123 20156
rect 31179 20154 31185 20156
rect 30939 20102 30941 20154
rect 31121 20102 31123 20154
rect 30877 20100 30883 20102
rect 30939 20100 30963 20102
rect 31019 20100 31043 20102
rect 31099 20100 31123 20102
rect 31179 20100 31185 20102
rect 30877 20091 31185 20100
rect 30748 20052 30800 20058
rect 30748 19994 30800 20000
rect 30576 19774 30696 19802
rect 30217 19612 30525 19621
rect 30217 19610 30223 19612
rect 30279 19610 30303 19612
rect 30359 19610 30383 19612
rect 30439 19610 30463 19612
rect 30519 19610 30525 19612
rect 30279 19558 30281 19610
rect 30461 19558 30463 19610
rect 30217 19556 30223 19558
rect 30279 19556 30303 19558
rect 30359 19556 30383 19558
rect 30439 19556 30463 19558
rect 30519 19556 30525 19558
rect 30217 19547 30525 19556
rect 30104 19508 30156 19514
rect 30104 19450 30156 19456
rect 29920 19440 29972 19446
rect 29920 19382 29972 19388
rect 29828 19236 29880 19242
rect 29828 19178 29880 19184
rect 29840 19145 29868 19178
rect 29826 19136 29882 19145
rect 29826 19071 29882 19080
rect 29828 18692 29880 18698
rect 29828 18634 29880 18640
rect 29840 18358 29868 18634
rect 29932 18630 29960 19382
rect 30012 19168 30064 19174
rect 30012 19110 30064 19116
rect 30024 18834 30052 19110
rect 30116 18834 30144 19450
rect 30288 19168 30340 19174
rect 30288 19110 30340 19116
rect 30300 18834 30328 19110
rect 30012 18828 30064 18834
rect 30012 18770 30064 18776
rect 30104 18828 30156 18834
rect 30104 18770 30156 18776
rect 30288 18828 30340 18834
rect 30288 18770 30340 18776
rect 29920 18624 29972 18630
rect 29920 18566 29972 18572
rect 29828 18352 29880 18358
rect 29828 18294 29880 18300
rect 29932 18086 29960 18566
rect 30116 18222 30144 18770
rect 30217 18524 30525 18533
rect 30217 18522 30223 18524
rect 30279 18522 30303 18524
rect 30359 18522 30383 18524
rect 30439 18522 30463 18524
rect 30519 18522 30525 18524
rect 30279 18470 30281 18522
rect 30461 18470 30463 18522
rect 30217 18468 30223 18470
rect 30279 18468 30303 18470
rect 30359 18468 30383 18470
rect 30439 18468 30463 18470
rect 30519 18468 30525 18470
rect 30217 18459 30525 18468
rect 30104 18216 30156 18222
rect 30104 18158 30156 18164
rect 30576 18154 30604 19774
rect 30656 19712 30708 19718
rect 30656 19654 30708 19660
rect 30668 19310 30696 19654
rect 30656 19304 30708 19310
rect 30656 19246 30708 19252
rect 31300 19304 31352 19310
rect 31300 19246 31352 19252
rect 30877 19068 31185 19077
rect 30877 19066 30883 19068
rect 30939 19066 30963 19068
rect 31019 19066 31043 19068
rect 31099 19066 31123 19068
rect 31179 19066 31185 19068
rect 30939 19014 30941 19066
rect 31121 19014 31123 19066
rect 30877 19012 30883 19014
rect 30939 19012 30963 19014
rect 31019 19012 31043 19014
rect 31099 19012 31123 19014
rect 31179 19012 31185 19014
rect 30877 19003 31185 19012
rect 30656 18896 30708 18902
rect 30656 18838 30708 18844
rect 30564 18148 30616 18154
rect 30564 18090 30616 18096
rect 29920 18080 29972 18086
rect 29920 18022 29972 18028
rect 30104 18080 30156 18086
rect 30104 18022 30156 18028
rect 30116 17882 30144 18022
rect 30104 17876 30156 17882
rect 30104 17818 30156 17824
rect 29920 17740 29972 17746
rect 29920 17682 29972 17688
rect 29828 17672 29880 17678
rect 29828 17614 29880 17620
rect 29736 17128 29788 17134
rect 29736 17070 29788 17076
rect 29748 16794 29776 17070
rect 29840 16794 29868 17614
rect 29736 16788 29788 16794
rect 29736 16730 29788 16736
rect 29828 16788 29880 16794
rect 29828 16730 29880 16736
rect 29656 16658 29776 16674
rect 29656 16652 29788 16658
rect 29656 16646 29736 16652
rect 29736 16594 29788 16600
rect 29644 16516 29696 16522
rect 29644 16458 29696 16464
rect 29656 16114 29684 16458
rect 29840 16454 29868 16730
rect 29932 16658 29960 17682
rect 30116 16794 30144 17818
rect 30217 17436 30525 17445
rect 30217 17434 30223 17436
rect 30279 17434 30303 17436
rect 30359 17434 30383 17436
rect 30439 17434 30463 17436
rect 30519 17434 30525 17436
rect 30279 17382 30281 17434
rect 30461 17382 30463 17434
rect 30217 17380 30223 17382
rect 30279 17380 30303 17382
rect 30359 17380 30383 17382
rect 30439 17380 30463 17382
rect 30519 17380 30525 17382
rect 30217 17371 30525 17380
rect 30576 17082 30604 18090
rect 30668 17814 30696 18838
rect 30840 18624 30892 18630
rect 30840 18566 30892 18572
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30656 17808 30708 17814
rect 30656 17750 30708 17756
rect 30656 17672 30708 17678
rect 30656 17614 30708 17620
rect 30484 17054 30604 17082
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30196 16720 30248 16726
rect 30196 16662 30248 16668
rect 29920 16652 29972 16658
rect 29920 16594 29972 16600
rect 29828 16448 29880 16454
rect 29828 16390 29880 16396
rect 29932 16250 29960 16594
rect 30208 16522 30236 16662
rect 30484 16590 30512 17054
rect 30564 16992 30616 16998
rect 30564 16934 30616 16940
rect 30576 16726 30604 16934
rect 30668 16794 30696 17614
rect 30760 17542 30788 18362
rect 30852 18222 30880 18566
rect 31208 18352 31260 18358
rect 31208 18294 31260 18300
rect 30840 18216 30892 18222
rect 30840 18158 30892 18164
rect 30877 17980 31185 17989
rect 30877 17978 30883 17980
rect 30939 17978 30963 17980
rect 31019 17978 31043 17980
rect 31099 17978 31123 17980
rect 31179 17978 31185 17980
rect 30939 17926 30941 17978
rect 31121 17926 31123 17978
rect 30877 17924 30883 17926
rect 30939 17924 30963 17926
rect 31019 17924 31043 17926
rect 31099 17924 31123 17926
rect 31179 17924 31185 17926
rect 30877 17915 31185 17924
rect 31220 17746 31248 18294
rect 31312 18222 31340 19246
rect 32036 18624 32088 18630
rect 32036 18566 32088 18572
rect 31300 18216 31352 18222
rect 31300 18158 31352 18164
rect 32048 18154 32076 18566
rect 32036 18148 32088 18154
rect 32036 18090 32088 18096
rect 31208 17740 31260 17746
rect 31208 17682 31260 17688
rect 32128 17672 32180 17678
rect 32128 17614 32180 17620
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 31024 17536 31076 17542
rect 31024 17478 31076 17484
rect 30656 16788 30708 16794
rect 30656 16730 30708 16736
rect 30564 16720 30616 16726
rect 30564 16662 30616 16668
rect 30760 16658 30788 17478
rect 31036 17338 31064 17478
rect 32140 17338 32168 17614
rect 31024 17332 31076 17338
rect 31024 17274 31076 17280
rect 32128 17332 32180 17338
rect 32128 17274 32180 17280
rect 32036 17060 32088 17066
rect 32036 17002 32088 17008
rect 31300 16992 31352 16998
rect 31300 16934 31352 16940
rect 30877 16892 31185 16901
rect 30877 16890 30883 16892
rect 30939 16890 30963 16892
rect 31019 16890 31043 16892
rect 31099 16890 31123 16892
rect 31179 16890 31185 16892
rect 30939 16838 30941 16890
rect 31121 16838 31123 16890
rect 30877 16836 30883 16838
rect 30939 16836 30963 16838
rect 31019 16836 31043 16838
rect 31099 16836 31123 16838
rect 31179 16836 31185 16838
rect 30877 16827 31185 16836
rect 31312 16794 31340 16934
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 30748 16652 30800 16658
rect 30748 16594 30800 16600
rect 30472 16584 30524 16590
rect 30472 16526 30524 16532
rect 30196 16516 30248 16522
rect 30196 16458 30248 16464
rect 30217 16348 30525 16357
rect 30217 16346 30223 16348
rect 30279 16346 30303 16348
rect 30359 16346 30383 16348
rect 30439 16346 30463 16348
rect 30519 16346 30525 16348
rect 30279 16294 30281 16346
rect 30461 16294 30463 16346
rect 30217 16292 30223 16294
rect 30279 16292 30303 16294
rect 30359 16292 30383 16294
rect 30439 16292 30463 16294
rect 30519 16292 30525 16294
rect 30217 16283 30525 16292
rect 32048 16250 32076 17002
rect 29920 16244 29972 16250
rect 29920 16186 29972 16192
rect 32036 16244 32088 16250
rect 32036 16186 32088 16192
rect 29932 16114 29960 16186
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29920 16108 29972 16114
rect 29920 16050 29972 16056
rect 31944 16040 31996 16046
rect 31944 15982 31996 15988
rect 32036 16040 32088 16046
rect 32036 15982 32088 15988
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 30564 15904 30616 15910
rect 30564 15846 30616 15852
rect 30576 15638 30604 15846
rect 30877 15804 31185 15813
rect 30877 15802 30883 15804
rect 30939 15802 30963 15804
rect 31019 15802 31043 15804
rect 31099 15802 31123 15804
rect 31179 15802 31185 15804
rect 30939 15750 30941 15802
rect 31121 15750 31123 15802
rect 30877 15748 30883 15750
rect 30939 15748 30963 15750
rect 31019 15748 31043 15750
rect 31099 15748 31123 15750
rect 31179 15748 31185 15750
rect 30877 15739 31185 15748
rect 29000 15632 29052 15638
rect 29000 15574 29052 15580
rect 30564 15632 30616 15638
rect 30564 15574 30616 15580
rect 31300 15632 31352 15638
rect 31300 15574 31352 15580
rect 29920 15564 29972 15570
rect 29920 15506 29972 15512
rect 28908 15496 28960 15502
rect 28908 15438 28960 15444
rect 28632 14418 28684 14424
rect 28736 14436 28856 14464
rect 28736 11218 28764 14436
rect 28816 14340 28868 14346
rect 28816 14282 28868 14288
rect 28828 13530 28856 14282
rect 28920 14278 28948 15438
rect 29828 14952 29880 14958
rect 29828 14894 29880 14900
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 29000 14544 29052 14550
rect 28998 14512 29000 14521
rect 29052 14512 29054 14521
rect 29472 14482 29500 14758
rect 29840 14618 29868 14894
rect 29828 14612 29880 14618
rect 29828 14554 29880 14560
rect 28998 14447 29054 14456
rect 29184 14476 29236 14482
rect 29184 14418 29236 14424
rect 29460 14476 29512 14482
rect 29460 14418 29512 14424
rect 29828 14476 29880 14482
rect 29828 14418 29880 14424
rect 28908 14272 28960 14278
rect 28908 14214 28960 14220
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 28920 14074 28948 14214
rect 28908 14068 28960 14074
rect 28908 14010 28960 14016
rect 29012 13870 29040 14214
rect 29092 14068 29144 14074
rect 29092 14010 29144 14016
rect 29104 13870 29132 14010
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29092 13864 29144 13870
rect 29092 13806 29144 13812
rect 28908 13728 28960 13734
rect 28908 13670 28960 13676
rect 29092 13728 29144 13734
rect 29092 13670 29144 13676
rect 28816 13524 28868 13530
rect 28816 13466 28868 13472
rect 28920 13394 28948 13670
rect 29104 13394 29132 13670
rect 29196 13530 29224 14418
rect 29840 13870 29868 14418
rect 29932 13870 29960 15506
rect 30217 15260 30525 15269
rect 30217 15258 30223 15260
rect 30279 15258 30303 15260
rect 30359 15258 30383 15260
rect 30439 15258 30463 15260
rect 30519 15258 30525 15260
rect 30279 15206 30281 15258
rect 30461 15206 30463 15258
rect 30217 15204 30223 15206
rect 30279 15204 30303 15206
rect 30359 15204 30383 15206
rect 30439 15204 30463 15206
rect 30519 15204 30525 15206
rect 30217 15195 30525 15204
rect 31312 15162 31340 15574
rect 31956 15434 31984 15982
rect 31944 15428 31996 15434
rect 31944 15370 31996 15376
rect 31852 15360 31904 15366
rect 31852 15302 31904 15308
rect 31300 15156 31352 15162
rect 31300 15098 31352 15104
rect 31864 15026 31892 15302
rect 31852 15020 31904 15026
rect 31852 14962 31904 14968
rect 30012 14952 30064 14958
rect 30012 14894 30064 14900
rect 30024 14618 30052 14894
rect 30656 14816 30708 14822
rect 30656 14758 30708 14764
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 30668 14618 30696 14758
rect 30877 14716 31185 14725
rect 30877 14714 30883 14716
rect 30939 14714 30963 14716
rect 31019 14714 31043 14716
rect 31099 14714 31123 14716
rect 31179 14714 31185 14716
rect 30939 14662 30941 14714
rect 31121 14662 31123 14714
rect 30877 14660 30883 14662
rect 30939 14660 30963 14662
rect 31019 14660 31043 14662
rect 31099 14660 31123 14662
rect 31179 14660 31185 14662
rect 30877 14651 31185 14660
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 31220 14550 31248 14758
rect 31208 14544 31260 14550
rect 31208 14486 31260 14492
rect 31864 14482 31892 14962
rect 32048 14890 32076 15982
rect 32036 14884 32088 14890
rect 32036 14826 32088 14832
rect 32128 14884 32180 14890
rect 32128 14826 32180 14832
rect 31852 14476 31904 14482
rect 31852 14418 31904 14424
rect 30012 14340 30064 14346
rect 30012 14282 30064 14288
rect 30024 13938 30052 14282
rect 30217 14172 30525 14181
rect 30217 14170 30223 14172
rect 30279 14170 30303 14172
rect 30359 14170 30383 14172
rect 30439 14170 30463 14172
rect 30519 14170 30525 14172
rect 30279 14118 30281 14170
rect 30461 14118 30463 14170
rect 30217 14116 30223 14118
rect 30279 14116 30303 14118
rect 30359 14116 30383 14118
rect 30439 14116 30463 14118
rect 30519 14116 30525 14118
rect 30217 14107 30525 14116
rect 32140 14074 32168 14826
rect 32128 14068 32180 14074
rect 32128 14010 32180 14016
rect 30012 13932 30064 13938
rect 30012 13874 30064 13880
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29920 13864 29972 13870
rect 31208 13864 31260 13870
rect 29920 13806 29972 13812
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 29460 13524 29512 13530
rect 29460 13466 29512 13472
rect 28908 13388 28960 13394
rect 28908 13330 28960 13336
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 28816 12980 28868 12986
rect 28816 12922 28868 12928
rect 28828 12850 28856 12922
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 28828 12322 28856 12786
rect 28920 12442 28948 13330
rect 29276 13252 29328 13258
rect 29276 13194 29328 13200
rect 29184 12776 29236 12782
rect 29184 12718 29236 12724
rect 29196 12594 29224 12718
rect 29012 12566 29224 12594
rect 28908 12436 28960 12442
rect 29012 12434 29040 12566
rect 29288 12442 29316 13194
rect 29276 12436 29328 12442
rect 29012 12406 29224 12434
rect 28908 12378 28960 12384
rect 29196 12322 29224 12406
rect 29276 12378 29328 12384
rect 28828 12306 29040 12322
rect 29196 12306 29316 12322
rect 28828 12300 29052 12306
rect 28828 12294 29000 12300
rect 28540 11212 28592 11218
rect 28540 11154 28592 11160
rect 28724 11212 28776 11218
rect 28724 11154 28776 11160
rect 28080 10804 28132 10810
rect 28080 10746 28132 10752
rect 27804 10600 27856 10606
rect 27804 10542 27856 10548
rect 27344 10260 27396 10266
rect 27344 10202 27396 10208
rect 26424 10192 26476 10198
rect 26424 10134 26476 10140
rect 26976 10124 27028 10130
rect 26976 10066 27028 10072
rect 27436 10124 27488 10130
rect 27436 10066 27488 10072
rect 25688 10056 25740 10062
rect 25688 9998 25740 10004
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 25228 9648 25280 9654
rect 25228 9590 25280 9596
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 24858 9480 24914 9489
rect 24858 9415 24914 9424
rect 24766 9208 24822 9217
rect 24766 9143 24822 9152
rect 24872 9042 24900 9415
rect 25240 9194 25268 9590
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25148 9178 25268 9194
rect 25136 9172 25268 9178
rect 25188 9166 25268 9172
rect 25136 9114 25188 9120
rect 25424 9042 25452 9386
rect 25700 9178 25728 9998
rect 26252 9654 26280 9998
rect 26240 9648 26292 9654
rect 26240 9590 26292 9596
rect 26252 9178 26280 9590
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 26344 9178 26372 9318
rect 25688 9172 25740 9178
rect 25688 9114 25740 9120
rect 26240 9172 26292 9178
rect 26240 9114 26292 9120
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 25228 9036 25280 9042
rect 25228 8978 25280 8984
rect 25412 9036 25464 9042
rect 25412 8978 25464 8984
rect 24952 8968 25004 8974
rect 24952 8910 25004 8916
rect 24860 8424 24912 8430
rect 24860 8366 24912 8372
rect 24492 8288 24544 8294
rect 24492 8230 24544 8236
rect 24504 6118 24532 8230
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24780 6662 24808 7822
rect 24872 7546 24900 8366
rect 24964 8090 24992 8910
rect 25240 8430 25268 8978
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25872 8968 25924 8974
rect 25872 8910 25924 8916
rect 26238 8936 26294 8945
rect 25320 8900 25372 8906
rect 25320 8842 25372 8848
rect 25332 8634 25360 8842
rect 25700 8634 25728 8910
rect 25320 8628 25372 8634
rect 25320 8570 25372 8576
rect 25688 8628 25740 8634
rect 25688 8570 25740 8576
rect 25228 8424 25280 8430
rect 25228 8366 25280 8372
rect 24952 8084 25004 8090
rect 24952 8026 25004 8032
rect 24860 7540 24912 7546
rect 24860 7482 24912 7488
rect 24964 7410 24992 8026
rect 24952 7404 25004 7410
rect 24952 7346 25004 7352
rect 25240 7274 25268 8366
rect 25136 7268 25188 7274
rect 25136 7210 25188 7216
rect 25228 7268 25280 7274
rect 25228 7210 25280 7216
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 24872 7002 24900 7142
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24768 6656 24820 6662
rect 24768 6598 24820 6604
rect 24860 6656 24912 6662
rect 24860 6598 24912 6604
rect 24492 6112 24544 6118
rect 24492 6054 24544 6060
rect 24492 5704 24544 5710
rect 24492 5646 24544 5652
rect 24400 3460 24452 3466
rect 24400 3402 24452 3408
rect 24504 3194 24532 5646
rect 24780 4826 24808 6598
rect 24872 6225 24900 6598
rect 25148 6458 25176 7210
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 25240 6254 25268 7210
rect 25332 6458 25360 8570
rect 25688 8356 25740 8362
rect 25688 8298 25740 8304
rect 25412 8016 25464 8022
rect 25412 7958 25464 7964
rect 25424 7546 25452 7958
rect 25504 7948 25556 7954
rect 25504 7890 25556 7896
rect 25412 7540 25464 7546
rect 25412 7482 25464 7488
rect 25516 6984 25544 7890
rect 25424 6956 25544 6984
rect 25424 6866 25452 6956
rect 25412 6860 25464 6866
rect 25412 6802 25464 6808
rect 25504 6860 25556 6866
rect 25504 6802 25556 6808
rect 25320 6452 25372 6458
rect 25320 6394 25372 6400
rect 25228 6248 25280 6254
rect 24858 6216 24914 6225
rect 25228 6190 25280 6196
rect 24858 6151 24914 6160
rect 24872 5710 24900 6151
rect 24952 6112 25004 6118
rect 24952 6054 25004 6060
rect 24860 5704 24912 5710
rect 24860 5646 24912 5652
rect 24964 5234 24992 6054
rect 25332 5846 25360 6394
rect 25516 5914 25544 6802
rect 25700 6798 25728 8298
rect 25780 7200 25832 7206
rect 25780 7142 25832 7148
rect 25792 6934 25820 7142
rect 25780 6928 25832 6934
rect 25780 6870 25832 6876
rect 25688 6792 25740 6798
rect 25688 6734 25740 6740
rect 25792 6186 25820 6870
rect 25780 6180 25832 6186
rect 25780 6122 25832 6128
rect 25688 6112 25740 6118
rect 25688 6054 25740 6060
rect 25504 5908 25556 5914
rect 25504 5850 25556 5856
rect 25320 5840 25372 5846
rect 25320 5782 25372 5788
rect 25410 5808 25466 5817
rect 25410 5743 25466 5752
rect 25424 5710 25452 5743
rect 25700 5710 25728 6054
rect 25228 5704 25280 5710
rect 25228 5646 25280 5652
rect 25412 5704 25464 5710
rect 25412 5646 25464 5652
rect 25688 5704 25740 5710
rect 25688 5646 25740 5652
rect 24952 5228 25004 5234
rect 24952 5170 25004 5176
rect 24768 4820 24820 4826
rect 24768 4762 24820 4768
rect 24952 4616 25004 4622
rect 24952 4558 25004 4564
rect 24964 4282 24992 4558
rect 24952 4276 25004 4282
rect 24952 4218 25004 4224
rect 25240 3194 25268 5646
rect 25424 5114 25452 5646
rect 25424 5086 25544 5114
rect 25412 5024 25464 5030
rect 25412 4966 25464 4972
rect 25424 4826 25452 4966
rect 25412 4820 25464 4826
rect 25412 4762 25464 4768
rect 25516 4146 25544 5086
rect 25596 4616 25648 4622
rect 25596 4558 25648 4564
rect 25608 4282 25636 4558
rect 25596 4276 25648 4282
rect 25596 4218 25648 4224
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 24492 3188 24544 3194
rect 24492 3130 24544 3136
rect 25228 3188 25280 3194
rect 25228 3130 25280 3136
rect 24308 3120 24360 3126
rect 24308 3062 24360 3068
rect 24584 3052 24636 3058
rect 24584 2994 24636 3000
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 22988 2748 23296 2757
rect 22988 2746 22994 2748
rect 23050 2746 23074 2748
rect 23130 2746 23154 2748
rect 23210 2746 23234 2748
rect 23290 2746 23296 2748
rect 23050 2694 23052 2746
rect 23232 2694 23234 2746
rect 22988 2692 22994 2694
rect 23050 2692 23074 2694
rect 23130 2692 23154 2694
rect 23210 2692 23234 2694
rect 23290 2692 23296 2694
rect 22988 2683 23296 2692
rect 23400 1578 23428 2926
rect 21928 1414 22048 1442
rect 23216 1550 23428 1578
rect 21928 800 21956 1414
rect 23216 800 23244 1550
rect 24596 1442 24624 2994
rect 25700 2854 25728 5646
rect 25884 3738 25912 8910
rect 26238 8871 26294 8880
rect 26252 6662 26280 8871
rect 26330 8664 26386 8673
rect 26330 8599 26332 8608
rect 26384 8599 26386 8608
rect 26332 8570 26384 8576
rect 26332 8424 26384 8430
rect 26332 8366 26384 8372
rect 26344 6798 26372 8366
rect 26436 8090 26464 9998
rect 26528 8430 26556 9998
rect 26988 9674 27016 10066
rect 27160 9920 27212 9926
rect 27160 9862 27212 9868
rect 26988 9646 27108 9674
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26804 9042 26832 9318
rect 26792 9036 26844 9042
rect 26792 8978 26844 8984
rect 26608 8968 26660 8974
rect 26608 8910 26660 8916
rect 26884 8968 26936 8974
rect 26884 8910 26936 8916
rect 26620 8650 26648 8910
rect 26620 8622 26832 8650
rect 26700 8560 26752 8566
rect 26700 8502 26752 8508
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26424 8084 26476 8090
rect 26476 8044 26556 8072
rect 26424 8026 26476 8032
rect 26424 7880 26476 7886
rect 26424 7822 26476 7828
rect 26436 7546 26464 7822
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26528 7002 26556 8044
rect 26516 6996 26568 7002
rect 26516 6938 26568 6944
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26240 6656 26292 6662
rect 26240 6598 26292 6604
rect 26252 6236 26280 6598
rect 26424 6248 26476 6254
rect 26252 6208 26424 6236
rect 26424 6190 26476 6196
rect 26712 5778 26740 8502
rect 26700 5772 26752 5778
rect 26700 5714 26752 5720
rect 26608 5296 26660 5302
rect 26608 5238 26660 5244
rect 25964 5228 26016 5234
rect 25964 5170 26016 5176
rect 25976 4622 26004 5170
rect 25964 4616 26016 4622
rect 25964 4558 26016 4564
rect 25976 3738 26004 4558
rect 26620 4146 26648 5238
rect 26712 5234 26740 5714
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 26608 4140 26660 4146
rect 26608 4082 26660 4088
rect 26804 3738 26832 8622
rect 26896 8566 26924 8910
rect 26884 8560 26936 8566
rect 26884 8502 26936 8508
rect 27080 8430 27108 9646
rect 27172 9450 27200 9862
rect 27160 9444 27212 9450
rect 27160 9386 27212 9392
rect 27448 8634 27476 10066
rect 28736 9722 28764 11154
rect 28828 10674 28856 12294
rect 29196 12300 29328 12306
rect 29196 12294 29276 12300
rect 29000 12242 29052 12248
rect 29276 12242 29328 12248
rect 29288 11898 29316 12242
rect 29276 11892 29328 11898
rect 29276 11834 29328 11840
rect 29184 11688 29236 11694
rect 29184 11630 29236 11636
rect 28908 11620 28960 11626
rect 28908 11562 28960 11568
rect 28920 11218 28948 11562
rect 29196 11354 29224 11630
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 28908 11212 28960 11218
rect 28908 11154 28960 11160
rect 29092 11212 29144 11218
rect 29092 11154 29144 11160
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28920 10470 28948 11154
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 28908 10464 28960 10470
rect 28908 10406 28960 10412
rect 29012 10146 29040 10542
rect 29104 10266 29132 11154
rect 29368 10600 29420 10606
rect 29368 10542 29420 10548
rect 29092 10260 29144 10266
rect 29092 10202 29144 10208
rect 28816 10124 28868 10130
rect 29012 10118 29132 10146
rect 28816 10066 28868 10072
rect 28724 9716 28776 9722
rect 28724 9658 28776 9664
rect 27804 9580 27856 9586
rect 27804 9522 27856 9528
rect 27528 8832 27580 8838
rect 27528 8774 27580 8780
rect 27620 8832 27672 8838
rect 27620 8774 27672 8780
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 27540 8430 27568 8774
rect 26884 8424 26936 8430
rect 26884 8366 26936 8372
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 27436 8424 27488 8430
rect 27436 8366 27488 8372
rect 27528 8424 27580 8430
rect 27528 8366 27580 8372
rect 26896 8294 26924 8366
rect 26884 8288 26936 8294
rect 26884 8230 26936 8236
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 27448 8276 27476 8366
rect 27632 8276 27660 8774
rect 27712 8356 27764 8362
rect 27712 8298 27764 8304
rect 27448 8248 27660 8276
rect 26896 6254 26924 8230
rect 26988 7274 27016 8230
rect 26976 7268 27028 7274
rect 26976 7210 27028 7216
rect 27448 7206 27476 8248
rect 27620 7268 27672 7274
rect 27620 7210 27672 7216
rect 27436 7200 27488 7206
rect 27436 7142 27488 7148
rect 26974 6352 27030 6361
rect 26974 6287 27030 6296
rect 26884 6248 26936 6254
rect 26884 6190 26936 6196
rect 26988 6186 27016 6287
rect 26976 6180 27028 6186
rect 26976 6122 27028 6128
rect 27252 6112 27304 6118
rect 27252 6054 27304 6060
rect 27264 5914 27292 6054
rect 27252 5908 27304 5914
rect 27252 5850 27304 5856
rect 27448 5778 27476 7142
rect 27632 7002 27660 7210
rect 27620 6996 27672 7002
rect 27620 6938 27672 6944
rect 27724 6866 27752 8298
rect 27816 7886 27844 9522
rect 28540 9444 28592 9450
rect 28540 9386 28592 9392
rect 28170 9208 28226 9217
rect 27896 9172 27948 9178
rect 28170 9143 28226 9152
rect 27896 9114 27948 9120
rect 27908 8498 27936 9114
rect 28184 8498 28212 9143
rect 28552 8974 28580 9386
rect 28828 9382 28856 10066
rect 29104 9926 29132 10118
rect 29380 10062 29408 10542
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 29092 9920 29144 9926
rect 29092 9862 29144 9868
rect 29000 9716 29052 9722
rect 29000 9658 29052 9664
rect 29012 9586 29040 9658
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 29104 9518 29132 9862
rect 29092 9512 29144 9518
rect 29092 9454 29144 9460
rect 28724 9376 28776 9382
rect 28724 9318 28776 9324
rect 28816 9376 28868 9382
rect 28816 9318 28868 9324
rect 28736 9178 28764 9318
rect 28724 9172 28776 9178
rect 28724 9114 28776 9120
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28460 8634 28488 8910
rect 29472 8634 29500 13466
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29564 12442 29592 12718
rect 29552 12436 29604 12442
rect 29552 12378 29604 12384
rect 29748 12374 29776 13806
rect 29736 12368 29788 12374
rect 29736 12310 29788 12316
rect 29644 11552 29696 11558
rect 29644 11494 29696 11500
rect 29656 11286 29684 11494
rect 29644 11280 29696 11286
rect 29644 11222 29696 11228
rect 29736 10260 29788 10266
rect 29736 10202 29788 10208
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29564 9178 29592 9522
rect 29748 9178 29776 10202
rect 29552 9172 29604 9178
rect 29552 9114 29604 9120
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 28448 8628 28500 8634
rect 28448 8570 28500 8576
rect 29000 8628 29052 8634
rect 29000 8570 29052 8576
rect 29460 8628 29512 8634
rect 29460 8570 29512 8576
rect 27896 8492 27948 8498
rect 27896 8434 27948 8440
rect 28172 8492 28224 8498
rect 28172 8434 28224 8440
rect 27908 8090 27936 8434
rect 29012 8430 29040 8570
rect 29472 8430 29500 8570
rect 28724 8424 28776 8430
rect 29000 8424 29052 8430
rect 28724 8366 28776 8372
rect 28998 8392 29000 8401
rect 29460 8424 29512 8430
rect 29052 8392 29054 8401
rect 28172 8288 28224 8294
rect 28172 8230 28224 8236
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27816 7410 27844 7822
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 28184 7342 28212 8230
rect 28172 7336 28224 7342
rect 28172 7278 28224 7284
rect 28630 6896 28686 6905
rect 27712 6860 27764 6866
rect 27712 6802 27764 6808
rect 27988 6860 28040 6866
rect 28630 6831 28632 6840
rect 27988 6802 28040 6808
rect 28684 6831 28686 6840
rect 28632 6802 28684 6808
rect 27712 6112 27764 6118
rect 27712 6054 27764 6060
rect 27436 5772 27488 5778
rect 27436 5714 27488 5720
rect 26884 4752 26936 4758
rect 26884 4694 26936 4700
rect 26896 4282 26924 4694
rect 27448 4690 27476 5714
rect 27620 5636 27672 5642
rect 27620 5578 27672 5584
rect 27528 5568 27580 5574
rect 27528 5510 27580 5516
rect 27540 5098 27568 5510
rect 27528 5092 27580 5098
rect 27528 5034 27580 5040
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27068 4480 27120 4486
rect 27068 4422 27120 4428
rect 26884 4276 26936 4282
rect 26884 4218 26936 4224
rect 25872 3732 25924 3738
rect 25872 3674 25924 3680
rect 25964 3732 26016 3738
rect 25964 3674 26016 3680
rect 26792 3732 26844 3738
rect 26792 3674 26844 3680
rect 27080 2990 27108 4422
rect 27448 4078 27476 4626
rect 27436 4072 27488 4078
rect 27436 4014 27488 4020
rect 27632 3194 27660 5578
rect 27724 5234 27752 6054
rect 28000 5914 28028 6802
rect 28448 6724 28500 6730
rect 28448 6666 28500 6672
rect 28460 6254 28488 6666
rect 28736 6254 28764 8366
rect 29460 8366 29512 8372
rect 29840 8362 29868 13806
rect 30208 13802 30420 13818
rect 31208 13806 31260 13812
rect 31484 13864 31536 13870
rect 31484 13806 31536 13812
rect 30196 13796 30420 13802
rect 30248 13790 30420 13796
rect 30196 13738 30248 13744
rect 30392 13530 30420 13790
rect 30564 13796 30616 13802
rect 30564 13738 30616 13744
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 30288 13524 30340 13530
rect 30288 13466 30340 13472
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30012 13388 30064 13394
rect 30012 13330 30064 13336
rect 30196 13388 30248 13394
rect 30196 13330 30248 13336
rect 29920 13320 29972 13326
rect 29920 13262 29972 13268
rect 29932 13190 29960 13262
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 29932 12170 29960 13126
rect 30024 12646 30052 13330
rect 30208 13274 30236 13330
rect 30300 13308 30328 13466
rect 30484 13462 30512 13670
rect 30472 13456 30524 13462
rect 30472 13398 30524 13404
rect 30576 13308 30604 13738
rect 30877 13628 31185 13637
rect 30877 13626 30883 13628
rect 30939 13626 30963 13628
rect 31019 13626 31043 13628
rect 31099 13626 31123 13628
rect 31179 13626 31185 13628
rect 30939 13574 30941 13626
rect 31121 13574 31123 13626
rect 30877 13572 30883 13574
rect 30939 13572 30963 13574
rect 31019 13572 31043 13574
rect 31099 13572 31123 13574
rect 31179 13572 31185 13574
rect 30877 13563 31185 13572
rect 30300 13280 30604 13308
rect 30116 13246 30236 13274
rect 30012 12640 30064 12646
rect 30012 12582 30064 12588
rect 30024 12374 30052 12582
rect 30116 12442 30144 13246
rect 30217 13084 30525 13093
rect 30217 13082 30223 13084
rect 30279 13082 30303 13084
rect 30359 13082 30383 13084
rect 30439 13082 30463 13084
rect 30519 13082 30525 13084
rect 30279 13030 30281 13082
rect 30461 13030 30463 13082
rect 30217 13028 30223 13030
rect 30279 13028 30303 13030
rect 30359 13028 30383 13030
rect 30439 13028 30463 13030
rect 30519 13028 30525 13030
rect 30217 13019 30525 13028
rect 30380 12776 30432 12782
rect 30380 12718 30432 12724
rect 30104 12436 30156 12442
rect 30104 12378 30156 12384
rect 30012 12368 30064 12374
rect 30012 12310 30064 12316
rect 30392 12238 30420 12718
rect 30877 12540 31185 12549
rect 30877 12538 30883 12540
rect 30939 12538 30963 12540
rect 31019 12538 31043 12540
rect 31099 12538 31123 12540
rect 31179 12538 31185 12540
rect 30939 12486 30941 12538
rect 31121 12486 31123 12538
rect 30877 12484 30883 12486
rect 30939 12484 30963 12486
rect 31019 12484 31043 12486
rect 31099 12484 31123 12486
rect 31179 12484 31185 12486
rect 30877 12475 31185 12484
rect 31220 12238 31248 13806
rect 31300 13728 31352 13734
rect 31300 13670 31352 13676
rect 31312 12850 31340 13670
rect 31496 13530 31524 13806
rect 31484 13524 31536 13530
rect 31484 13466 31536 13472
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31760 12640 31812 12646
rect 31760 12582 31812 12588
rect 31772 12374 31800 12582
rect 31300 12368 31352 12374
rect 31300 12310 31352 12316
rect 31760 12368 31812 12374
rect 31760 12310 31812 12316
rect 31942 12336 31998 12345
rect 30380 12232 30432 12238
rect 30380 12174 30432 12180
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 30217 11996 30525 12005
rect 30217 11994 30223 11996
rect 30279 11994 30303 11996
rect 30359 11994 30383 11996
rect 30439 11994 30463 11996
rect 30519 11994 30525 11996
rect 30279 11942 30281 11994
rect 30461 11942 30463 11994
rect 30217 11940 30223 11942
rect 30279 11940 30303 11942
rect 30359 11940 30383 11942
rect 30439 11940 30463 11942
rect 30519 11940 30525 11942
rect 30217 11931 30525 11940
rect 31312 11898 31340 12310
rect 31942 12271 31998 12280
rect 31956 11898 31984 12271
rect 32128 12096 32180 12102
rect 32128 12038 32180 12044
rect 31300 11892 31352 11898
rect 31300 11834 31352 11840
rect 31944 11892 31996 11898
rect 31944 11834 31996 11840
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30668 11354 30696 11630
rect 31956 11626 31984 11834
rect 31944 11620 31996 11626
rect 31944 11562 31996 11568
rect 31208 11552 31260 11558
rect 31208 11494 31260 11500
rect 30877 11452 31185 11461
rect 30877 11450 30883 11452
rect 30939 11450 30963 11452
rect 31019 11450 31043 11452
rect 31099 11450 31123 11452
rect 31179 11450 31185 11452
rect 30939 11398 30941 11450
rect 31121 11398 31123 11450
rect 30877 11396 30883 11398
rect 30939 11396 30963 11398
rect 31019 11396 31043 11398
rect 31099 11396 31123 11398
rect 31179 11396 31185 11398
rect 30877 11387 31185 11396
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30932 11348 30984 11354
rect 30932 11290 30984 11296
rect 30217 10908 30525 10917
rect 30217 10906 30223 10908
rect 30279 10906 30303 10908
rect 30359 10906 30383 10908
rect 30439 10906 30463 10908
rect 30519 10906 30525 10908
rect 30279 10854 30281 10906
rect 30461 10854 30463 10906
rect 30217 10852 30223 10854
rect 30279 10852 30303 10854
rect 30359 10852 30383 10854
rect 30439 10852 30463 10854
rect 30519 10852 30525 10854
rect 30217 10843 30525 10852
rect 30944 10606 30972 11290
rect 31220 11218 31248 11494
rect 32140 11286 32168 12038
rect 32128 11280 32180 11286
rect 32128 11222 32180 11228
rect 31208 11212 31260 11218
rect 31208 11154 31260 11160
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 29920 10600 29972 10606
rect 29920 10542 29972 10548
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 30932 10600 30984 10606
rect 30932 10542 30984 10548
rect 29932 9722 29960 10542
rect 30024 10198 30052 10542
rect 30196 10464 30248 10470
rect 30196 10406 30248 10412
rect 30656 10464 30708 10470
rect 30656 10406 30708 10412
rect 30208 10198 30236 10406
rect 30012 10192 30064 10198
rect 30012 10134 30064 10140
rect 30196 10192 30248 10198
rect 30196 10134 30248 10140
rect 30217 9820 30525 9829
rect 30217 9818 30223 9820
rect 30279 9818 30303 9820
rect 30359 9818 30383 9820
rect 30439 9818 30463 9820
rect 30519 9818 30525 9820
rect 30279 9766 30281 9818
rect 30461 9766 30463 9818
rect 30217 9764 30223 9766
rect 30279 9764 30303 9766
rect 30359 9764 30383 9766
rect 30439 9764 30463 9766
rect 30519 9764 30525 9766
rect 30217 9755 30525 9764
rect 29920 9716 29972 9722
rect 29920 9658 29972 9664
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 29932 8634 29960 8910
rect 30668 8838 30696 10406
rect 30877 10364 31185 10373
rect 30877 10362 30883 10364
rect 30939 10362 30963 10364
rect 31019 10362 31043 10364
rect 31099 10362 31123 10364
rect 31179 10362 31185 10364
rect 30939 10310 30941 10362
rect 31121 10310 31123 10362
rect 30877 10308 30883 10310
rect 30939 10308 30963 10310
rect 31019 10308 31043 10310
rect 31099 10308 31123 10310
rect 31179 10308 31185 10310
rect 30877 10299 31185 10308
rect 31680 10266 31708 11086
rect 31208 10260 31260 10266
rect 31208 10202 31260 10208
rect 31668 10260 31720 10266
rect 31668 10202 31720 10208
rect 30877 9276 31185 9285
rect 30877 9274 30883 9276
rect 30939 9274 30963 9276
rect 31019 9274 31043 9276
rect 31099 9274 31123 9276
rect 31179 9274 31185 9276
rect 30939 9222 30941 9274
rect 31121 9222 31123 9274
rect 30877 9220 30883 9222
rect 30939 9220 30963 9222
rect 31019 9220 31043 9222
rect 31099 9220 31123 9222
rect 31179 9220 31185 9222
rect 30877 9211 31185 9220
rect 30656 8832 30708 8838
rect 30656 8774 30708 8780
rect 30217 8732 30525 8741
rect 30217 8730 30223 8732
rect 30279 8730 30303 8732
rect 30359 8730 30383 8732
rect 30439 8730 30463 8732
rect 30519 8730 30525 8732
rect 30279 8678 30281 8730
rect 30461 8678 30463 8730
rect 30217 8676 30223 8678
rect 30279 8676 30303 8678
rect 30359 8676 30383 8678
rect 30439 8676 30463 8678
rect 30519 8676 30525 8678
rect 30217 8667 30525 8676
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 28998 8327 29054 8336
rect 29092 8356 29144 8362
rect 29092 8298 29144 8304
rect 29276 8356 29328 8362
rect 29276 8298 29328 8304
rect 29828 8356 29880 8362
rect 29828 8298 29880 8304
rect 29104 8090 29132 8298
rect 29288 8129 29316 8298
rect 29274 8120 29330 8129
rect 29092 8084 29144 8090
rect 30562 8120 30618 8129
rect 29274 8055 29330 8064
rect 30196 8084 30248 8090
rect 29092 8026 29144 8032
rect 30562 8055 30618 8064
rect 30196 8026 30248 8032
rect 28816 8016 28868 8022
rect 28816 7958 28868 7964
rect 28828 7546 28856 7958
rect 28908 7880 28960 7886
rect 28908 7822 28960 7828
rect 28920 7546 28948 7822
rect 30012 7744 30064 7750
rect 30208 7732 30236 8026
rect 30576 7954 30604 8055
rect 30564 7948 30616 7954
rect 30564 7890 30616 7896
rect 30012 7686 30064 7692
rect 30116 7704 30236 7732
rect 30024 7546 30052 7686
rect 28816 7540 28868 7546
rect 28816 7482 28868 7488
rect 28908 7540 28960 7546
rect 28908 7482 28960 7488
rect 30012 7540 30064 7546
rect 30012 7482 30064 7488
rect 30116 7002 30144 7704
rect 30217 7644 30525 7653
rect 30217 7642 30223 7644
rect 30279 7642 30303 7644
rect 30359 7642 30383 7644
rect 30439 7642 30463 7644
rect 30519 7642 30525 7644
rect 30279 7590 30281 7642
rect 30461 7590 30463 7642
rect 30217 7588 30223 7590
rect 30279 7588 30303 7590
rect 30359 7588 30383 7590
rect 30439 7588 30463 7590
rect 30519 7588 30525 7590
rect 30217 7579 30525 7588
rect 30668 7546 30696 8774
rect 31220 8498 31248 10202
rect 31392 10124 31444 10130
rect 31392 10066 31444 10072
rect 31404 9722 31432 10066
rect 31392 9716 31444 9722
rect 31392 9658 31444 9664
rect 31208 8492 31260 8498
rect 31208 8434 31260 8440
rect 30877 8188 31185 8197
rect 30877 8186 30883 8188
rect 30939 8186 30963 8188
rect 31019 8186 31043 8188
rect 31099 8186 31123 8188
rect 31179 8186 31185 8188
rect 30939 8134 30941 8186
rect 31121 8134 31123 8186
rect 30877 8132 30883 8134
rect 30939 8132 30963 8134
rect 31019 8132 31043 8134
rect 31099 8132 31123 8134
rect 31179 8132 31185 8134
rect 30877 8123 31185 8132
rect 30748 7880 30800 7886
rect 30748 7822 30800 7828
rect 30656 7540 30708 7546
rect 30656 7482 30708 7488
rect 30196 7404 30248 7410
rect 30196 7346 30248 7352
rect 30104 6996 30156 7002
rect 30104 6938 30156 6944
rect 29460 6724 29512 6730
rect 29460 6666 29512 6672
rect 29196 6446 29408 6474
rect 29196 6390 29224 6446
rect 29184 6384 29236 6390
rect 29184 6326 29236 6332
rect 28816 6316 28868 6322
rect 28868 6276 28948 6304
rect 28816 6258 28868 6264
rect 28448 6248 28500 6254
rect 28448 6190 28500 6196
rect 28724 6248 28776 6254
rect 28724 6190 28776 6196
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 27804 5704 27856 5710
rect 28172 5704 28224 5710
rect 27804 5646 27856 5652
rect 28170 5672 28172 5681
rect 28224 5672 28226 5681
rect 27816 5370 27844 5646
rect 28170 5607 28226 5616
rect 27804 5364 27856 5370
rect 27804 5306 27856 5312
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 28184 4826 28212 5607
rect 28448 5228 28500 5234
rect 28448 5170 28500 5176
rect 28172 4820 28224 4826
rect 28172 4762 28224 4768
rect 28460 4282 28488 5170
rect 28632 5160 28684 5166
rect 28632 5102 28684 5108
rect 28540 5024 28592 5030
rect 28540 4966 28592 4972
rect 28448 4276 28500 4282
rect 28448 4218 28500 4224
rect 28552 4146 28580 4966
rect 28644 4826 28672 5102
rect 28632 4820 28684 4826
rect 28632 4762 28684 4768
rect 28736 4554 28764 6190
rect 28920 6118 28948 6276
rect 28908 6112 28960 6118
rect 28908 6054 28960 6060
rect 28920 5302 28948 6054
rect 29276 5908 29328 5914
rect 29276 5850 29328 5856
rect 29184 5840 29236 5846
rect 29184 5782 29236 5788
rect 28908 5296 28960 5302
rect 28908 5238 28960 5244
rect 29196 5234 29224 5782
rect 29184 5228 29236 5234
rect 29184 5170 29236 5176
rect 29288 5114 29316 5850
rect 29380 5710 29408 6446
rect 29472 6390 29500 6666
rect 30208 6662 30236 7346
rect 30760 7002 30788 7822
rect 31220 7410 31248 8434
rect 31208 7404 31260 7410
rect 31208 7346 31260 7352
rect 31208 7200 31260 7206
rect 31208 7142 31260 7148
rect 30877 7100 31185 7109
rect 30877 7098 30883 7100
rect 30939 7098 30963 7100
rect 31019 7098 31043 7100
rect 31099 7098 31123 7100
rect 31179 7098 31185 7100
rect 30939 7046 30941 7098
rect 31121 7046 31123 7098
rect 30877 7044 30883 7046
rect 30939 7044 30963 7046
rect 31019 7044 31043 7046
rect 31099 7044 31123 7046
rect 31179 7044 31185 7046
rect 30877 7035 31185 7044
rect 30748 6996 30800 7002
rect 30748 6938 30800 6944
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30012 6656 30064 6662
rect 30012 6598 30064 6604
rect 30196 6656 30248 6662
rect 30196 6598 30248 6604
rect 30024 6458 30052 6598
rect 30217 6556 30525 6565
rect 30217 6554 30223 6556
rect 30279 6554 30303 6556
rect 30359 6554 30383 6556
rect 30439 6554 30463 6556
rect 30519 6554 30525 6556
rect 30279 6502 30281 6554
rect 30461 6502 30463 6554
rect 30217 6500 30223 6502
rect 30279 6500 30303 6502
rect 30359 6500 30383 6502
rect 30439 6500 30463 6502
rect 30519 6500 30525 6502
rect 30217 6491 30525 6500
rect 30576 6458 30604 6802
rect 31220 6798 31248 7142
rect 31208 6792 31260 6798
rect 31208 6734 31260 6740
rect 30748 6656 30800 6662
rect 30748 6598 30800 6604
rect 30012 6452 30064 6458
rect 30012 6394 30064 6400
rect 30564 6452 30616 6458
rect 30564 6394 30616 6400
rect 29460 6384 29512 6390
rect 29460 6326 29512 6332
rect 30564 6316 30616 6322
rect 30564 6258 30616 6264
rect 30576 5914 30604 6258
rect 30656 6180 30708 6186
rect 30656 6122 30708 6128
rect 30668 5914 30696 6122
rect 30564 5908 30616 5914
rect 30564 5850 30616 5856
rect 30656 5908 30708 5914
rect 30656 5850 30708 5856
rect 30012 5772 30064 5778
rect 30012 5714 30064 5720
rect 30760 5760 30788 6598
rect 30877 6012 31185 6021
rect 30877 6010 30883 6012
rect 30939 6010 30963 6012
rect 31019 6010 31043 6012
rect 31099 6010 31123 6012
rect 31179 6010 31185 6012
rect 30939 5958 30941 6010
rect 31121 5958 31123 6010
rect 30877 5956 30883 5958
rect 30939 5956 30963 5958
rect 31019 5956 31043 5958
rect 31099 5956 31123 5958
rect 31179 5956 31185 5958
rect 30877 5947 31185 5956
rect 30840 5772 30892 5778
rect 30760 5732 30840 5760
rect 29368 5704 29420 5710
rect 29368 5646 29420 5652
rect 29552 5704 29604 5710
rect 29552 5646 29604 5652
rect 29012 5086 29316 5114
rect 29012 4826 29040 5086
rect 29092 5024 29144 5030
rect 29092 4966 29144 4972
rect 29104 4826 29132 4966
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 29092 4820 29144 4826
rect 29092 4762 29144 4768
rect 29564 4758 29592 5646
rect 30024 5370 30052 5714
rect 30217 5468 30525 5477
rect 30217 5466 30223 5468
rect 30279 5466 30303 5468
rect 30359 5466 30383 5468
rect 30439 5466 30463 5468
rect 30519 5466 30525 5468
rect 30279 5414 30281 5466
rect 30461 5414 30463 5466
rect 30217 5412 30223 5414
rect 30279 5412 30303 5414
rect 30359 5412 30383 5414
rect 30439 5412 30463 5414
rect 30519 5412 30525 5414
rect 30217 5403 30525 5412
rect 30012 5364 30064 5370
rect 30012 5306 30064 5312
rect 30760 5234 30788 5732
rect 30840 5714 30892 5720
rect 31220 5302 31248 6734
rect 31404 6458 31432 9658
rect 32036 8832 32088 8838
rect 32036 8774 32088 8780
rect 31576 8424 31628 8430
rect 31576 8366 31628 8372
rect 31484 6656 31536 6662
rect 31484 6598 31536 6604
rect 31392 6452 31444 6458
rect 31392 6394 31444 6400
rect 31496 5710 31524 6598
rect 31484 5704 31536 5710
rect 31484 5646 31536 5652
rect 31208 5296 31260 5302
rect 31208 5238 31260 5244
rect 30748 5228 30800 5234
rect 30748 5170 30800 5176
rect 29828 5160 29880 5166
rect 29828 5102 29880 5108
rect 30012 5160 30064 5166
rect 30012 5102 30064 5108
rect 29552 4752 29604 4758
rect 29552 4694 29604 4700
rect 28908 4616 28960 4622
rect 28908 4558 28960 4564
rect 28724 4548 28776 4554
rect 28724 4490 28776 4496
rect 28540 4140 28592 4146
rect 28540 4082 28592 4088
rect 28724 4140 28776 4146
rect 28724 4082 28776 4088
rect 28736 3738 28764 4082
rect 28920 3942 28948 4558
rect 29552 4480 29604 4486
rect 29552 4422 29604 4428
rect 29564 4078 29592 4422
rect 29840 4282 29868 5102
rect 30024 4690 30052 5102
rect 30012 4684 30064 4690
rect 30012 4626 30064 4632
rect 30760 4622 30788 5170
rect 31208 5024 31260 5030
rect 31208 4966 31260 4972
rect 30877 4924 31185 4933
rect 30877 4922 30883 4924
rect 30939 4922 30963 4924
rect 31019 4922 31043 4924
rect 31099 4922 31123 4924
rect 31179 4922 31185 4924
rect 30939 4870 30941 4922
rect 31121 4870 31123 4922
rect 30877 4868 30883 4870
rect 30939 4868 30963 4870
rect 31019 4868 31043 4870
rect 31099 4868 31123 4870
rect 31179 4868 31185 4870
rect 30877 4859 31185 4868
rect 31220 4826 31248 4966
rect 31208 4820 31260 4826
rect 31208 4762 31260 4768
rect 30748 4616 30800 4622
rect 30748 4558 30800 4564
rect 30217 4380 30525 4389
rect 30217 4378 30223 4380
rect 30279 4378 30303 4380
rect 30359 4378 30383 4380
rect 30439 4378 30463 4380
rect 30519 4378 30525 4380
rect 30279 4326 30281 4378
rect 30461 4326 30463 4378
rect 30217 4324 30223 4326
rect 30279 4324 30303 4326
rect 30359 4324 30383 4326
rect 30439 4324 30463 4326
rect 30519 4324 30525 4326
rect 30217 4315 30525 4324
rect 29828 4276 29880 4282
rect 29828 4218 29880 4224
rect 29552 4072 29604 4078
rect 29552 4014 29604 4020
rect 28908 3936 28960 3942
rect 28908 3878 28960 3884
rect 29000 3936 29052 3942
rect 29000 3878 29052 3884
rect 28920 3738 28948 3878
rect 28724 3732 28776 3738
rect 28724 3674 28776 3680
rect 28908 3732 28960 3738
rect 28908 3674 28960 3680
rect 29012 3670 29040 3878
rect 29000 3664 29052 3670
rect 29000 3606 29052 3612
rect 27620 3188 27672 3194
rect 27620 3130 27672 3136
rect 27160 3052 27212 3058
rect 27160 2994 27212 3000
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 25780 2984 25832 2990
rect 25780 2926 25832 2932
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 25688 2848 25740 2854
rect 25688 2790 25740 2796
rect 24504 1414 24624 1442
rect 24504 800 24532 1414
rect 25792 800 25820 2926
rect 27172 1442 27200 2994
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 27080 1414 27200 1442
rect 27080 800 27108 1414
rect 28368 800 28396 2926
rect 29748 1442 29776 2994
rect 29840 2990 29868 4218
rect 30877 3836 31185 3845
rect 30877 3834 30883 3836
rect 30939 3834 30963 3836
rect 31019 3834 31043 3836
rect 31099 3834 31123 3836
rect 31179 3834 31185 3836
rect 30939 3782 30941 3834
rect 31121 3782 31123 3834
rect 30877 3780 30883 3782
rect 30939 3780 30963 3782
rect 31019 3780 31043 3782
rect 31099 3780 31123 3782
rect 31179 3780 31185 3782
rect 30877 3771 31185 3780
rect 30217 3292 30525 3301
rect 30217 3290 30223 3292
rect 30279 3290 30303 3292
rect 30359 3290 30383 3292
rect 30439 3290 30463 3292
rect 30519 3290 30525 3292
rect 30279 3238 30281 3290
rect 30461 3238 30463 3290
rect 30217 3236 30223 3238
rect 30279 3236 30303 3238
rect 30359 3236 30383 3238
rect 30439 3236 30463 3238
rect 30519 3236 30525 3238
rect 30217 3227 30525 3236
rect 31588 3194 31616 8366
rect 31852 8288 31904 8294
rect 31852 8230 31904 8236
rect 31864 7546 31892 8230
rect 31852 7540 31904 7546
rect 31852 7482 31904 7488
rect 32048 7410 32076 8774
rect 32036 7404 32088 7410
rect 32036 7346 32088 7352
rect 32036 6724 32088 6730
rect 32036 6666 32088 6672
rect 32048 6322 32076 6666
rect 32036 6316 32088 6322
rect 32036 6258 32088 6264
rect 31760 5908 31812 5914
rect 31760 5850 31812 5856
rect 31772 5234 31800 5850
rect 31944 5840 31996 5846
rect 31944 5782 31996 5788
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 31956 4826 31984 5782
rect 32232 5681 32260 22066
rect 32404 21888 32456 21894
rect 32404 21830 32456 21836
rect 32416 21690 32444 21830
rect 32404 21684 32456 21690
rect 32404 21626 32456 21632
rect 32588 21480 32640 21486
rect 32588 21422 32640 21428
rect 32600 21146 32628 21422
rect 32588 21140 32640 21146
rect 32588 21082 32640 21088
rect 32312 20936 32364 20942
rect 32312 20878 32364 20884
rect 32324 20058 32352 20878
rect 32588 20800 32640 20806
rect 32588 20742 32640 20748
rect 32600 20466 32628 20742
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32312 20052 32364 20058
rect 32312 19994 32364 20000
rect 32404 20052 32456 20058
rect 32404 19994 32456 20000
rect 32324 19854 32352 19994
rect 32416 19961 32444 19994
rect 32402 19952 32458 19961
rect 32402 19887 32458 19896
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32508 18970 32536 19110
rect 32496 18964 32548 18970
rect 32496 18906 32548 18912
rect 32404 18148 32456 18154
rect 32404 18090 32456 18096
rect 32416 17882 32444 18090
rect 32404 17876 32456 17882
rect 32404 17818 32456 17824
rect 32404 15904 32456 15910
rect 32404 15846 32456 15852
rect 32416 15706 32444 15846
rect 32404 15700 32456 15706
rect 32404 15642 32456 15648
rect 32312 14476 32364 14482
rect 32312 14418 32364 14424
rect 32324 13462 32352 14418
rect 32404 14272 32456 14278
rect 32404 14214 32456 14220
rect 32416 14074 32444 14214
rect 32404 14068 32456 14074
rect 32404 14010 32456 14016
rect 32312 13456 32364 13462
rect 32312 13398 32364 13404
rect 32588 13388 32640 13394
rect 32588 13330 32640 13336
rect 32312 13320 32364 13326
rect 32312 13262 32364 13268
rect 32324 12986 32352 13262
rect 32312 12980 32364 12986
rect 32312 12922 32364 12928
rect 32600 12306 32628 13330
rect 32692 12345 32720 26982
rect 33416 26920 33468 26926
rect 33416 26862 33468 26868
rect 33048 26376 33100 26382
rect 33048 26318 33100 26324
rect 33060 25945 33088 26318
rect 33046 25936 33102 25945
rect 33046 25871 33102 25880
rect 33048 25696 33100 25702
rect 33048 25638 33100 25644
rect 32772 22500 32824 22506
rect 32772 22442 32824 22448
rect 32784 22234 32812 22442
rect 32772 22228 32824 22234
rect 32772 22170 32824 22176
rect 32772 19984 32824 19990
rect 32772 19926 32824 19932
rect 32784 19310 32812 19926
rect 33060 19854 33088 25638
rect 33428 22642 33456 26862
rect 33796 23662 33824 27270
rect 33784 23656 33836 23662
rect 33784 23598 33836 23604
rect 33416 22636 33468 22642
rect 33416 22578 33468 22584
rect 33428 21010 33456 22578
rect 33784 22432 33836 22438
rect 33784 22374 33836 22380
rect 33796 22094 33824 22374
rect 33796 22066 34008 22094
rect 33416 21004 33468 21010
rect 33416 20946 33468 20952
rect 33140 20936 33192 20942
rect 33140 20878 33192 20884
rect 33324 20936 33376 20942
rect 33324 20878 33376 20884
rect 33152 19922 33180 20878
rect 33140 19916 33192 19922
rect 33140 19858 33192 19864
rect 33336 19854 33364 20878
rect 33876 20800 33928 20806
rect 33876 20742 33928 20748
rect 33888 20398 33916 20742
rect 33876 20392 33928 20398
rect 33876 20334 33928 20340
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33324 19848 33376 19854
rect 33324 19790 33376 19796
rect 33782 19816 33838 19825
rect 32772 19304 32824 19310
rect 32772 19246 32824 19252
rect 33060 19174 33088 19790
rect 33782 19751 33838 19760
rect 33796 19378 33824 19751
rect 33784 19372 33836 19378
rect 33784 19314 33836 19320
rect 33048 19168 33100 19174
rect 33048 19110 33100 19116
rect 33692 19168 33744 19174
rect 33692 19110 33744 19116
rect 32956 18828 33008 18834
rect 32956 18770 33008 18776
rect 33508 18828 33560 18834
rect 33508 18770 33560 18776
rect 32968 18306 32996 18770
rect 32968 18278 33088 18306
rect 33520 18290 33548 18770
rect 33704 18290 33732 19110
rect 32956 18216 33008 18222
rect 32956 18158 33008 18164
rect 32968 17202 32996 18158
rect 33060 17762 33088 18278
rect 33508 18284 33560 18290
rect 33508 18226 33560 18232
rect 33692 18284 33744 18290
rect 33692 18226 33744 18232
rect 33520 17882 33548 18226
rect 33600 18080 33652 18086
rect 33600 18022 33652 18028
rect 33508 17876 33560 17882
rect 33508 17818 33560 17824
rect 33060 17746 33180 17762
rect 33060 17740 33192 17746
rect 33060 17734 33140 17740
rect 33140 17682 33192 17688
rect 32956 17196 33008 17202
rect 32956 17138 33008 17144
rect 32968 15706 32996 17138
rect 33046 17096 33102 17105
rect 33046 17031 33102 17040
rect 33060 16590 33088 17031
rect 33048 16584 33100 16590
rect 33048 16526 33100 16532
rect 33152 16114 33180 17682
rect 33612 17202 33640 18022
rect 33600 17196 33652 17202
rect 33600 17138 33652 17144
rect 33140 16108 33192 16114
rect 33140 16050 33192 16056
rect 32956 15700 33008 15706
rect 32956 15642 33008 15648
rect 33152 15570 33180 16050
rect 33600 16040 33652 16046
rect 33600 15982 33652 15988
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 33152 15314 33180 15506
rect 33060 15286 33180 15314
rect 32864 14408 32916 14414
rect 32864 14350 32916 14356
rect 32876 14074 32904 14350
rect 32864 14068 32916 14074
rect 32864 14010 32916 14016
rect 33060 13530 33088 15286
rect 33612 15162 33640 15982
rect 33600 15156 33652 15162
rect 33600 15098 33652 15104
rect 33508 14272 33560 14278
rect 33508 14214 33560 14220
rect 33048 13524 33100 13530
rect 33048 13466 33100 13472
rect 33520 12442 33548 14214
rect 33612 13938 33640 15098
rect 33704 14414 33732 18226
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33888 14958 33916 15302
rect 33876 14952 33928 14958
rect 33876 14894 33928 14900
rect 33692 14408 33744 14414
rect 33692 14350 33744 14356
rect 33600 13932 33652 13938
rect 33600 13874 33652 13880
rect 33508 12436 33560 12442
rect 33508 12378 33560 12384
rect 32678 12336 32734 12345
rect 32588 12300 32640 12306
rect 32678 12271 32734 12280
rect 32588 12242 32640 12248
rect 32680 12232 32732 12238
rect 32680 12174 32732 12180
rect 32692 11898 32720 12174
rect 33048 12096 33100 12102
rect 33048 12038 33100 12044
rect 32680 11892 32732 11898
rect 32680 11834 32732 11840
rect 33060 11694 33088 12038
rect 33520 11762 33548 12378
rect 33508 11756 33560 11762
rect 33508 11698 33560 11704
rect 33048 11688 33100 11694
rect 33048 11630 33100 11636
rect 32588 11552 32640 11558
rect 32588 11494 32640 11500
rect 32600 11150 32628 11494
rect 32588 11144 32640 11150
rect 32588 11086 32640 11092
rect 32600 10606 32628 11086
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32588 8968 32640 8974
rect 32588 8910 32640 8916
rect 32600 8090 32628 8910
rect 33416 8900 33468 8906
rect 33416 8842 33468 8848
rect 32588 8084 32640 8090
rect 32588 8026 32640 8032
rect 33428 7954 33456 8842
rect 33520 8634 33548 11698
rect 33784 9920 33836 9926
rect 33784 9862 33836 9868
rect 33796 9081 33824 9862
rect 33980 9654 34008 22066
rect 33968 9648 34020 9654
rect 33968 9590 34020 9596
rect 33782 9072 33838 9081
rect 33782 9007 33838 9016
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 32588 7948 32640 7954
rect 32588 7890 32640 7896
rect 33416 7948 33468 7954
rect 33416 7890 33468 7896
rect 32312 7880 32364 7886
rect 32312 7822 32364 7828
rect 32324 7274 32352 7822
rect 32312 7268 32364 7274
rect 32312 7210 32364 7216
rect 32324 6866 32352 7210
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 32600 6254 32628 7890
rect 33520 7886 33548 8570
rect 33784 8560 33836 8566
rect 33782 8528 33784 8537
rect 33836 8528 33838 8537
rect 33782 8463 33838 8472
rect 32680 7880 32732 7886
rect 32680 7822 32732 7828
rect 33508 7880 33560 7886
rect 33508 7822 33560 7828
rect 32692 7002 32720 7822
rect 33692 7268 33744 7274
rect 33692 7210 33744 7216
rect 32680 6996 32732 7002
rect 32680 6938 32732 6944
rect 33704 6458 33732 7210
rect 33692 6452 33744 6458
rect 33692 6394 33744 6400
rect 32588 6248 32640 6254
rect 32588 6190 32640 6196
rect 32312 6112 32364 6118
rect 32312 6054 32364 6060
rect 32864 6112 32916 6118
rect 32864 6054 32916 6060
rect 33784 6112 33836 6118
rect 33784 6054 33836 6060
rect 32218 5672 32274 5681
rect 32218 5607 32274 5616
rect 32324 5522 32352 6054
rect 32876 5914 32904 6054
rect 32864 5908 32916 5914
rect 32864 5850 32916 5856
rect 33796 5778 33824 6054
rect 34072 5817 34100 30058
rect 35176 30025 35204 30126
rect 35162 30016 35218 30025
rect 35162 29951 35218 29960
rect 35164 27396 35216 27402
rect 35164 27338 35216 27344
rect 35176 27305 35204 27338
rect 35162 27296 35218 27305
rect 35162 27231 35218 27240
rect 34704 24200 34756 24206
rect 34704 24142 34756 24148
rect 34716 23905 34744 24142
rect 34702 23896 34758 23905
rect 34702 23831 34758 23840
rect 35164 22568 35216 22574
rect 35162 22536 35164 22545
rect 35216 22536 35218 22545
rect 35162 22471 35218 22480
rect 34888 21412 34940 21418
rect 34888 21354 34940 21360
rect 34900 21185 34928 21354
rect 34886 21176 34942 21185
rect 34886 21111 34942 21120
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34532 18465 34560 18702
rect 34518 18456 34574 18465
rect 34518 18391 34574 18400
rect 34888 15972 34940 15978
rect 34888 15914 34940 15920
rect 34900 15745 34928 15914
rect 34886 15736 34942 15745
rect 34886 15671 34942 15680
rect 35162 13696 35218 13705
rect 35162 13631 35218 13640
rect 35176 13530 35204 13631
rect 35164 13524 35216 13530
rect 35164 13466 35216 13472
rect 34428 12776 34480 12782
rect 34428 12718 34480 12724
rect 34440 12345 34468 12718
rect 34426 12336 34482 12345
rect 34426 12271 34482 12280
rect 34886 10976 34942 10985
rect 34886 10911 34942 10920
rect 34900 10674 34928 10911
rect 34888 10668 34940 10674
rect 34888 10610 34940 10616
rect 34428 10056 34480 10062
rect 34428 9998 34480 10004
rect 34440 9625 34468 9998
rect 34426 9616 34482 9625
rect 34426 9551 34482 9560
rect 34428 8356 34480 8362
rect 34428 8298 34480 8304
rect 34440 8265 34468 8298
rect 34426 8256 34482 8265
rect 34426 8191 34482 8200
rect 34702 6896 34758 6905
rect 34702 6831 34704 6840
rect 34756 6831 34758 6840
rect 34704 6802 34756 6808
rect 34058 5808 34114 5817
rect 33784 5772 33836 5778
rect 34058 5743 34114 5752
rect 33784 5714 33836 5720
rect 33140 5636 33192 5642
rect 33140 5578 33192 5584
rect 32404 5568 32456 5574
rect 32324 5516 32404 5522
rect 32324 5510 32456 5516
rect 32324 5494 32444 5510
rect 32036 5024 32088 5030
rect 32036 4966 32088 4972
rect 32220 5024 32272 5030
rect 32220 4966 32272 4972
rect 31944 4820 31996 4826
rect 31944 4762 31996 4768
rect 31576 3188 31628 3194
rect 31576 3130 31628 3136
rect 31956 2990 31984 4762
rect 32048 4758 32076 4966
rect 32036 4752 32088 4758
rect 32036 4694 32088 4700
rect 32232 4690 32260 4966
rect 32220 4684 32272 4690
rect 32220 4626 32272 4632
rect 32324 3602 32352 5494
rect 33152 5098 33180 5578
rect 34886 5536 34942 5545
rect 34886 5471 34942 5480
rect 34900 5234 34928 5471
rect 34888 5228 34940 5234
rect 34888 5170 34940 5176
rect 33140 5092 33192 5098
rect 33140 5034 33192 5040
rect 34704 4616 34756 4622
rect 34704 4558 34756 4564
rect 34716 4185 34744 4558
rect 34702 4176 34758 4185
rect 34702 4111 34758 4120
rect 33968 4072 34020 4078
rect 33968 4014 34020 4020
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 32312 3596 32364 3602
rect 32312 3538 32364 3544
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 32864 3052 32916 3058
rect 32864 2994 32916 3000
rect 29828 2984 29880 2990
rect 29828 2926 29880 2932
rect 31576 2984 31628 2990
rect 31576 2926 31628 2932
rect 31944 2984 31996 2990
rect 31944 2926 31996 2932
rect 30877 2748 31185 2757
rect 30877 2746 30883 2748
rect 30939 2746 30963 2748
rect 31019 2746 31043 2748
rect 31099 2746 31123 2748
rect 31179 2746 31185 2748
rect 30939 2694 30941 2746
rect 31121 2694 31123 2746
rect 30877 2692 30883 2694
rect 30939 2692 30963 2694
rect 31019 2692 31043 2694
rect 31099 2692 31123 2694
rect 31179 2692 31185 2694
rect 30877 2683 31185 2692
rect 29656 1414 29776 1442
rect 29656 800 29684 1414
rect 31588 800 31616 2926
rect 32876 800 32904 2994
rect 33060 921 33088 3470
rect 33980 2122 34008 4014
rect 34440 2145 34468 4014
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 34426 2136 34482 2145
rect 33980 2094 34192 2122
rect 33046 912 33102 921
rect 33046 847 33102 856
rect 34164 800 34192 2094
rect 34426 2071 34482 2080
rect 35452 800 35480 3538
rect 36728 2984 36780 2990
rect 36728 2926 36780 2932
rect 36740 800 36768 2926
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 6458 0 6514 800
rect 7746 0 7802 800
rect 9034 0 9090 800
rect 10966 0 11022 800
rect 12254 0 12310 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 16118 0 16174 800
rect 17406 0 17462 800
rect 18694 0 18750 800
rect 20626 0 20682 800
rect 21914 0 21970 800
rect 23202 0 23258 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 36726 0 36782 800
<< via2 >>
rect 3790 36080 3846 36136
rect 3054 34720 3110 34776
rect 3238 33360 3294 33416
rect 7216 34298 7272 34300
rect 7296 34298 7352 34300
rect 7376 34298 7432 34300
rect 7456 34298 7512 34300
rect 7216 34246 7262 34298
rect 7262 34246 7272 34298
rect 7296 34246 7326 34298
rect 7326 34246 7338 34298
rect 7338 34246 7352 34298
rect 7376 34246 7390 34298
rect 7390 34246 7402 34298
rect 7402 34246 7432 34298
rect 7456 34246 7466 34298
rect 7466 34246 7512 34298
rect 7216 34244 7272 34246
rect 7296 34244 7352 34246
rect 7376 34244 7432 34246
rect 7456 34244 7512 34246
rect 4434 32308 4436 32328
rect 4436 32308 4488 32328
rect 4488 32308 4490 32328
rect 4434 32272 4490 32308
rect 3238 31320 3294 31376
rect 1306 29960 1362 30016
rect 1306 28620 1362 28656
rect 1306 28600 1308 28620
rect 1308 28600 1360 28620
rect 1360 28600 1362 28620
rect 1306 27240 1362 27296
rect 6556 33754 6612 33756
rect 6636 33754 6692 33756
rect 6716 33754 6772 33756
rect 6796 33754 6852 33756
rect 6556 33702 6602 33754
rect 6602 33702 6612 33754
rect 6636 33702 6666 33754
rect 6666 33702 6678 33754
rect 6678 33702 6692 33754
rect 6716 33702 6730 33754
rect 6730 33702 6742 33754
rect 6742 33702 6772 33754
rect 6796 33702 6806 33754
rect 6806 33702 6852 33754
rect 6556 33700 6612 33702
rect 6636 33700 6692 33702
rect 6716 33700 6772 33702
rect 6796 33700 6852 33702
rect 7216 33210 7272 33212
rect 7296 33210 7352 33212
rect 7376 33210 7432 33212
rect 7456 33210 7512 33212
rect 7216 33158 7262 33210
rect 7262 33158 7272 33210
rect 7296 33158 7326 33210
rect 7326 33158 7338 33210
rect 7338 33158 7352 33210
rect 7376 33158 7390 33210
rect 7390 33158 7402 33210
rect 7402 33158 7432 33210
rect 7456 33158 7466 33210
rect 7466 33158 7512 33210
rect 7216 33156 7272 33158
rect 7296 33156 7352 33158
rect 7376 33156 7432 33158
rect 7456 33156 7512 33158
rect 6556 32666 6612 32668
rect 6636 32666 6692 32668
rect 6716 32666 6772 32668
rect 6796 32666 6852 32668
rect 6556 32614 6602 32666
rect 6602 32614 6612 32666
rect 6636 32614 6666 32666
rect 6666 32614 6678 32666
rect 6678 32614 6692 32666
rect 6716 32614 6730 32666
rect 6730 32614 6742 32666
rect 6742 32614 6772 32666
rect 6796 32614 6806 32666
rect 6806 32614 6852 32666
rect 6556 32612 6612 32614
rect 6636 32612 6692 32614
rect 6716 32612 6772 32614
rect 6796 32612 6852 32614
rect 1306 24520 1362 24576
rect 1306 21120 1362 21176
rect 1306 18400 1362 18456
rect 1306 17060 1362 17096
rect 1306 17040 1308 17060
rect 1308 17040 1360 17060
rect 1360 17040 1362 17060
rect 1306 15680 1362 15736
rect 1306 14320 1362 14376
rect 1306 12960 1362 13016
rect 1306 11600 1362 11656
rect 1306 9580 1362 9616
rect 1306 9560 1308 9580
rect 1308 9560 1360 9580
rect 1360 9560 1362 9580
rect 3238 25880 3294 25936
rect 3514 23160 3570 23216
rect 3238 19760 3294 19816
rect 4342 24792 4398 24848
rect 6556 31578 6612 31580
rect 6636 31578 6692 31580
rect 6716 31578 6772 31580
rect 6796 31578 6852 31580
rect 6556 31526 6602 31578
rect 6602 31526 6612 31578
rect 6636 31526 6666 31578
rect 6666 31526 6678 31578
rect 6678 31526 6692 31578
rect 6716 31526 6730 31578
rect 6730 31526 6742 31578
rect 6742 31526 6772 31578
rect 6796 31526 6806 31578
rect 6806 31526 6852 31578
rect 6556 31524 6612 31526
rect 6636 31524 6692 31526
rect 6716 31524 6772 31526
rect 6796 31524 6852 31526
rect 7216 32122 7272 32124
rect 7296 32122 7352 32124
rect 7376 32122 7432 32124
rect 7456 32122 7512 32124
rect 7216 32070 7262 32122
rect 7262 32070 7272 32122
rect 7296 32070 7326 32122
rect 7326 32070 7338 32122
rect 7338 32070 7352 32122
rect 7376 32070 7390 32122
rect 7390 32070 7402 32122
rect 7402 32070 7432 32122
rect 7456 32070 7466 32122
rect 7466 32070 7512 32122
rect 7216 32068 7272 32070
rect 7296 32068 7352 32070
rect 7376 32068 7432 32070
rect 7456 32068 7512 32070
rect 6556 30490 6612 30492
rect 6636 30490 6692 30492
rect 6716 30490 6772 30492
rect 6796 30490 6852 30492
rect 6556 30438 6602 30490
rect 6602 30438 6612 30490
rect 6636 30438 6666 30490
rect 6666 30438 6678 30490
rect 6678 30438 6692 30490
rect 6716 30438 6730 30490
rect 6730 30438 6742 30490
rect 6742 30438 6772 30490
rect 6796 30438 6806 30490
rect 6806 30438 6852 30490
rect 6556 30436 6612 30438
rect 6636 30436 6692 30438
rect 6716 30436 6772 30438
rect 6796 30436 6852 30438
rect 7216 31034 7272 31036
rect 7296 31034 7352 31036
rect 7376 31034 7432 31036
rect 7456 31034 7512 31036
rect 7216 30982 7262 31034
rect 7262 30982 7272 31034
rect 7296 30982 7326 31034
rect 7326 30982 7338 31034
rect 7338 30982 7352 31034
rect 7376 30982 7390 31034
rect 7390 30982 7402 31034
rect 7402 30982 7432 31034
rect 7456 30982 7466 31034
rect 7466 30982 7512 31034
rect 7216 30980 7272 30982
rect 7296 30980 7352 30982
rect 7376 30980 7432 30982
rect 7456 30980 7512 30982
rect 6556 29402 6612 29404
rect 6636 29402 6692 29404
rect 6716 29402 6772 29404
rect 6796 29402 6852 29404
rect 6556 29350 6602 29402
rect 6602 29350 6612 29402
rect 6636 29350 6666 29402
rect 6666 29350 6678 29402
rect 6678 29350 6692 29402
rect 6716 29350 6730 29402
rect 6730 29350 6742 29402
rect 6742 29350 6772 29402
rect 6796 29350 6806 29402
rect 6806 29350 6852 29402
rect 6556 29348 6612 29350
rect 6636 29348 6692 29350
rect 6716 29348 6772 29350
rect 6796 29348 6852 29350
rect 5906 24928 5962 24984
rect 7216 29946 7272 29948
rect 7296 29946 7352 29948
rect 7376 29946 7432 29948
rect 7456 29946 7512 29948
rect 7216 29894 7262 29946
rect 7262 29894 7272 29946
rect 7296 29894 7326 29946
rect 7326 29894 7338 29946
rect 7338 29894 7352 29946
rect 7376 29894 7390 29946
rect 7390 29894 7402 29946
rect 7402 29894 7432 29946
rect 7456 29894 7466 29946
rect 7466 29894 7512 29946
rect 7216 29892 7272 29894
rect 7296 29892 7352 29894
rect 7376 29892 7432 29894
rect 7456 29892 7512 29894
rect 7216 28858 7272 28860
rect 7296 28858 7352 28860
rect 7376 28858 7432 28860
rect 7456 28858 7512 28860
rect 7216 28806 7262 28858
rect 7262 28806 7272 28858
rect 7296 28806 7326 28858
rect 7326 28806 7338 28858
rect 7338 28806 7352 28858
rect 7376 28806 7390 28858
rect 7390 28806 7402 28858
rect 7402 28806 7432 28858
rect 7456 28806 7466 28858
rect 7466 28806 7512 28858
rect 7216 28804 7272 28806
rect 7296 28804 7352 28806
rect 7376 28804 7432 28806
rect 7456 28804 7512 28806
rect 6556 28314 6612 28316
rect 6636 28314 6692 28316
rect 6716 28314 6772 28316
rect 6796 28314 6852 28316
rect 6556 28262 6602 28314
rect 6602 28262 6612 28314
rect 6636 28262 6666 28314
rect 6666 28262 6678 28314
rect 6678 28262 6692 28314
rect 6716 28262 6730 28314
rect 6730 28262 6742 28314
rect 6742 28262 6772 28314
rect 6796 28262 6806 28314
rect 6806 28262 6852 28314
rect 6556 28260 6612 28262
rect 6636 28260 6692 28262
rect 6716 28260 6772 28262
rect 6796 28260 6852 28262
rect 7216 27770 7272 27772
rect 7296 27770 7352 27772
rect 7376 27770 7432 27772
rect 7456 27770 7512 27772
rect 7216 27718 7262 27770
rect 7262 27718 7272 27770
rect 7296 27718 7326 27770
rect 7326 27718 7338 27770
rect 7338 27718 7352 27770
rect 7376 27718 7390 27770
rect 7390 27718 7402 27770
rect 7402 27718 7432 27770
rect 7456 27718 7466 27770
rect 7466 27718 7512 27770
rect 7216 27716 7272 27718
rect 7296 27716 7352 27718
rect 7376 27716 7432 27718
rect 7456 27716 7512 27718
rect 6556 27226 6612 27228
rect 6636 27226 6692 27228
rect 6716 27226 6772 27228
rect 6796 27226 6852 27228
rect 6556 27174 6602 27226
rect 6602 27174 6612 27226
rect 6636 27174 6666 27226
rect 6666 27174 6678 27226
rect 6678 27174 6692 27226
rect 6716 27174 6730 27226
rect 6730 27174 6742 27226
rect 6742 27174 6772 27226
rect 6796 27174 6806 27226
rect 6806 27174 6852 27226
rect 6556 27172 6612 27174
rect 6636 27172 6692 27174
rect 6716 27172 6772 27174
rect 6796 27172 6852 27174
rect 6556 26138 6612 26140
rect 6636 26138 6692 26140
rect 6716 26138 6772 26140
rect 6796 26138 6852 26140
rect 6556 26086 6602 26138
rect 6602 26086 6612 26138
rect 6636 26086 6666 26138
rect 6666 26086 6678 26138
rect 6678 26086 6692 26138
rect 6716 26086 6730 26138
rect 6730 26086 6742 26138
rect 6742 26086 6772 26138
rect 6796 26086 6806 26138
rect 6806 26086 6852 26138
rect 6556 26084 6612 26086
rect 6636 26084 6692 26086
rect 6716 26084 6772 26086
rect 6796 26084 6852 26086
rect 5814 23468 5816 23488
rect 5816 23468 5868 23488
rect 5868 23468 5870 23488
rect 5814 23432 5870 23468
rect 5170 19352 5226 19408
rect 5538 21004 5594 21040
rect 5538 20984 5540 21004
rect 5540 20984 5592 21004
rect 5592 20984 5594 21004
rect 6556 25050 6612 25052
rect 6636 25050 6692 25052
rect 6716 25050 6772 25052
rect 6796 25050 6852 25052
rect 6556 24998 6602 25050
rect 6602 24998 6612 25050
rect 6636 24998 6666 25050
rect 6666 24998 6678 25050
rect 6678 24998 6692 25050
rect 6716 24998 6730 25050
rect 6730 24998 6742 25050
rect 6742 24998 6772 25050
rect 6796 24998 6806 25050
rect 6806 24998 6852 25050
rect 6556 24996 6612 24998
rect 6636 24996 6692 24998
rect 6716 24996 6772 24998
rect 6796 24996 6852 24998
rect 6556 23962 6612 23964
rect 6636 23962 6692 23964
rect 6716 23962 6772 23964
rect 6796 23962 6852 23964
rect 6556 23910 6602 23962
rect 6602 23910 6612 23962
rect 6636 23910 6666 23962
rect 6666 23910 6678 23962
rect 6678 23910 6692 23962
rect 6716 23910 6730 23962
rect 6730 23910 6742 23962
rect 6742 23910 6772 23962
rect 6796 23910 6806 23962
rect 6806 23910 6852 23962
rect 6556 23908 6612 23910
rect 6636 23908 6692 23910
rect 6716 23908 6772 23910
rect 6796 23908 6852 23910
rect 6182 23568 6238 23624
rect 6556 22874 6612 22876
rect 6636 22874 6692 22876
rect 6716 22874 6772 22876
rect 6796 22874 6852 22876
rect 6556 22822 6602 22874
rect 6602 22822 6612 22874
rect 6636 22822 6666 22874
rect 6666 22822 6678 22874
rect 6678 22822 6692 22874
rect 6716 22822 6730 22874
rect 6730 22822 6742 22874
rect 6742 22822 6772 22874
rect 6796 22822 6806 22874
rect 6806 22822 6852 22874
rect 6556 22820 6612 22822
rect 6636 22820 6692 22822
rect 6716 22820 6772 22822
rect 6796 22820 6852 22822
rect 6556 21786 6612 21788
rect 6636 21786 6692 21788
rect 6716 21786 6772 21788
rect 6796 21786 6852 21788
rect 6556 21734 6602 21786
rect 6602 21734 6612 21786
rect 6636 21734 6666 21786
rect 6666 21734 6678 21786
rect 6678 21734 6692 21786
rect 6716 21734 6730 21786
rect 6730 21734 6742 21786
rect 6742 21734 6772 21786
rect 6796 21734 6806 21786
rect 6806 21734 6852 21786
rect 6556 21732 6612 21734
rect 6636 21732 6692 21734
rect 6716 21732 6772 21734
rect 6796 21732 6852 21734
rect 5814 20168 5870 20224
rect 1306 8200 1362 8256
rect 3514 6840 3570 6896
rect 5722 18284 5778 18320
rect 5722 18264 5724 18284
rect 5724 18264 5776 18284
rect 5776 18264 5778 18284
rect 7216 26682 7272 26684
rect 7296 26682 7352 26684
rect 7376 26682 7432 26684
rect 7456 26682 7512 26684
rect 7216 26630 7262 26682
rect 7262 26630 7272 26682
rect 7296 26630 7326 26682
rect 7326 26630 7338 26682
rect 7338 26630 7352 26682
rect 7376 26630 7390 26682
rect 7390 26630 7402 26682
rect 7402 26630 7432 26682
rect 7456 26630 7466 26682
rect 7466 26630 7512 26682
rect 7216 26628 7272 26630
rect 7296 26628 7352 26630
rect 7376 26628 7432 26630
rect 7456 26628 7512 26630
rect 7216 25594 7272 25596
rect 7296 25594 7352 25596
rect 7376 25594 7432 25596
rect 7456 25594 7512 25596
rect 7216 25542 7262 25594
rect 7262 25542 7272 25594
rect 7296 25542 7326 25594
rect 7326 25542 7338 25594
rect 7338 25542 7352 25594
rect 7376 25542 7390 25594
rect 7390 25542 7402 25594
rect 7402 25542 7432 25594
rect 7456 25542 7466 25594
rect 7466 25542 7512 25594
rect 7216 25540 7272 25542
rect 7296 25540 7352 25542
rect 7376 25540 7432 25542
rect 7456 25540 7512 25542
rect 7216 24506 7272 24508
rect 7296 24506 7352 24508
rect 7376 24506 7432 24508
rect 7456 24506 7512 24508
rect 7216 24454 7262 24506
rect 7262 24454 7272 24506
rect 7296 24454 7326 24506
rect 7326 24454 7338 24506
rect 7338 24454 7352 24506
rect 7376 24454 7390 24506
rect 7390 24454 7402 24506
rect 7402 24454 7432 24506
rect 7456 24454 7466 24506
rect 7466 24454 7512 24506
rect 7216 24452 7272 24454
rect 7296 24452 7352 24454
rect 7376 24452 7432 24454
rect 7456 24452 7512 24454
rect 7216 23418 7272 23420
rect 7296 23418 7352 23420
rect 7376 23418 7432 23420
rect 7456 23418 7512 23420
rect 7216 23366 7262 23418
rect 7262 23366 7272 23418
rect 7296 23366 7326 23418
rect 7326 23366 7338 23418
rect 7338 23366 7352 23418
rect 7376 23366 7390 23418
rect 7390 23366 7402 23418
rect 7402 23366 7432 23418
rect 7456 23366 7466 23418
rect 7466 23366 7512 23418
rect 7216 23364 7272 23366
rect 7296 23364 7352 23366
rect 7376 23364 7432 23366
rect 7456 23364 7512 23366
rect 7216 22330 7272 22332
rect 7296 22330 7352 22332
rect 7376 22330 7432 22332
rect 7456 22330 7512 22332
rect 7216 22278 7262 22330
rect 7262 22278 7272 22330
rect 7296 22278 7326 22330
rect 7326 22278 7338 22330
rect 7338 22278 7352 22330
rect 7376 22278 7390 22330
rect 7390 22278 7402 22330
rect 7402 22278 7432 22330
rect 7456 22278 7466 22330
rect 7466 22278 7512 22330
rect 7216 22276 7272 22278
rect 7296 22276 7352 22278
rect 7376 22276 7432 22278
rect 7456 22276 7512 22278
rect 10874 33224 10930 33280
rect 11426 33224 11482 33280
rect 15105 34298 15161 34300
rect 15185 34298 15241 34300
rect 15265 34298 15321 34300
rect 15345 34298 15401 34300
rect 15105 34246 15151 34298
rect 15151 34246 15161 34298
rect 15185 34246 15215 34298
rect 15215 34246 15227 34298
rect 15227 34246 15241 34298
rect 15265 34246 15279 34298
rect 15279 34246 15291 34298
rect 15291 34246 15321 34298
rect 15345 34246 15355 34298
rect 15355 34246 15401 34298
rect 15105 34244 15161 34246
rect 15185 34244 15241 34246
rect 15265 34244 15321 34246
rect 15345 34244 15401 34246
rect 11610 33088 11666 33144
rect 11058 32816 11114 32872
rect 12070 32952 12126 33008
rect 12070 32816 12126 32872
rect 14445 33754 14501 33756
rect 14525 33754 14581 33756
rect 14605 33754 14661 33756
rect 14685 33754 14741 33756
rect 14445 33702 14491 33754
rect 14491 33702 14501 33754
rect 14525 33702 14555 33754
rect 14555 33702 14567 33754
rect 14567 33702 14581 33754
rect 14605 33702 14619 33754
rect 14619 33702 14631 33754
rect 14631 33702 14661 33754
rect 14685 33702 14695 33754
rect 14695 33702 14741 33754
rect 14445 33700 14501 33702
rect 14525 33700 14581 33702
rect 14605 33700 14661 33702
rect 14685 33700 14741 33702
rect 13082 33224 13138 33280
rect 13266 32408 13322 32464
rect 15105 33210 15161 33212
rect 15185 33210 15241 33212
rect 15265 33210 15321 33212
rect 15345 33210 15401 33212
rect 15105 33158 15151 33210
rect 15151 33158 15161 33210
rect 15185 33158 15215 33210
rect 15215 33158 15227 33210
rect 15227 33158 15241 33210
rect 15265 33158 15279 33210
rect 15279 33158 15291 33210
rect 15291 33158 15321 33210
rect 15345 33158 15355 33210
rect 15355 33158 15401 33210
rect 15105 33156 15161 33158
rect 15185 33156 15241 33158
rect 15265 33156 15321 33158
rect 15345 33156 15401 33158
rect 14002 32972 14058 33008
rect 14002 32952 14004 32972
rect 14004 32952 14056 32972
rect 14056 32952 14058 32972
rect 8114 24656 8170 24712
rect 7216 21242 7272 21244
rect 7296 21242 7352 21244
rect 7376 21242 7432 21244
rect 7456 21242 7512 21244
rect 7216 21190 7262 21242
rect 7262 21190 7272 21242
rect 7296 21190 7326 21242
rect 7326 21190 7338 21242
rect 7338 21190 7352 21242
rect 7376 21190 7390 21242
rect 7390 21190 7402 21242
rect 7402 21190 7432 21242
rect 7456 21190 7466 21242
rect 7466 21190 7512 21242
rect 7216 21188 7272 21190
rect 7296 21188 7352 21190
rect 7376 21188 7432 21190
rect 7456 21188 7512 21190
rect 5722 15136 5778 15192
rect 4066 7828 4068 7848
rect 4068 7828 4120 7848
rect 4120 7828 4122 7848
rect 4066 7792 4122 7828
rect 5722 9560 5778 9616
rect 6366 19352 6422 19408
rect 6556 20698 6612 20700
rect 6636 20698 6692 20700
rect 6716 20698 6772 20700
rect 6796 20698 6852 20700
rect 6556 20646 6602 20698
rect 6602 20646 6612 20698
rect 6636 20646 6666 20698
rect 6666 20646 6678 20698
rect 6678 20646 6692 20698
rect 6716 20646 6730 20698
rect 6730 20646 6742 20698
rect 6742 20646 6772 20698
rect 6796 20646 6806 20698
rect 6806 20646 6852 20698
rect 6556 20644 6612 20646
rect 6636 20644 6692 20646
rect 6716 20644 6772 20646
rect 6796 20644 6852 20646
rect 6556 19610 6612 19612
rect 6636 19610 6692 19612
rect 6716 19610 6772 19612
rect 6796 19610 6852 19612
rect 6556 19558 6602 19610
rect 6602 19558 6612 19610
rect 6636 19558 6666 19610
rect 6666 19558 6678 19610
rect 6678 19558 6692 19610
rect 6716 19558 6730 19610
rect 6730 19558 6742 19610
rect 6742 19558 6772 19610
rect 6796 19558 6806 19610
rect 6806 19558 6852 19610
rect 6556 19556 6612 19558
rect 6636 19556 6692 19558
rect 6716 19556 6772 19558
rect 6796 19556 6852 19558
rect 6734 19216 6790 19272
rect 6556 18522 6612 18524
rect 6636 18522 6692 18524
rect 6716 18522 6772 18524
rect 6796 18522 6852 18524
rect 6556 18470 6602 18522
rect 6602 18470 6612 18522
rect 6636 18470 6666 18522
rect 6666 18470 6678 18522
rect 6678 18470 6692 18522
rect 6716 18470 6730 18522
rect 6730 18470 6742 18522
rect 6742 18470 6772 18522
rect 6796 18470 6806 18522
rect 6806 18470 6852 18522
rect 6556 18468 6612 18470
rect 6636 18468 6692 18470
rect 6716 18468 6772 18470
rect 6796 18468 6852 18470
rect 7216 20154 7272 20156
rect 7296 20154 7352 20156
rect 7376 20154 7432 20156
rect 7456 20154 7512 20156
rect 7216 20102 7262 20154
rect 7262 20102 7272 20154
rect 7296 20102 7326 20154
rect 7326 20102 7338 20154
rect 7338 20102 7352 20154
rect 7376 20102 7390 20154
rect 7390 20102 7402 20154
rect 7402 20102 7432 20154
rect 7456 20102 7466 20154
rect 7466 20102 7512 20154
rect 7216 20100 7272 20102
rect 7296 20100 7352 20102
rect 7376 20100 7432 20102
rect 7456 20100 7512 20102
rect 7216 19066 7272 19068
rect 7296 19066 7352 19068
rect 7376 19066 7432 19068
rect 7456 19066 7512 19068
rect 7216 19014 7262 19066
rect 7262 19014 7272 19066
rect 7296 19014 7326 19066
rect 7326 19014 7338 19066
rect 7338 19014 7352 19066
rect 7376 19014 7390 19066
rect 7390 19014 7402 19066
rect 7402 19014 7432 19066
rect 7456 19014 7466 19066
rect 7466 19014 7512 19066
rect 7216 19012 7272 19014
rect 7296 19012 7352 19014
rect 7376 19012 7432 19014
rect 7456 19012 7512 19014
rect 7216 17978 7272 17980
rect 7296 17978 7352 17980
rect 7376 17978 7432 17980
rect 7456 17978 7512 17980
rect 7216 17926 7262 17978
rect 7262 17926 7272 17978
rect 7296 17926 7326 17978
rect 7326 17926 7338 17978
rect 7338 17926 7352 17978
rect 7376 17926 7390 17978
rect 7390 17926 7402 17978
rect 7402 17926 7432 17978
rect 7456 17926 7466 17978
rect 7466 17926 7512 17978
rect 7216 17924 7272 17926
rect 7296 17924 7352 17926
rect 7376 17924 7432 17926
rect 7456 17924 7512 17926
rect 6556 17434 6612 17436
rect 6636 17434 6692 17436
rect 6716 17434 6772 17436
rect 6796 17434 6852 17436
rect 6556 17382 6602 17434
rect 6602 17382 6612 17434
rect 6636 17382 6666 17434
rect 6666 17382 6678 17434
rect 6678 17382 6692 17434
rect 6716 17382 6730 17434
rect 6730 17382 6742 17434
rect 6742 17382 6772 17434
rect 6796 17382 6806 17434
rect 6806 17382 6852 17434
rect 6556 17380 6612 17382
rect 6636 17380 6692 17382
rect 6716 17380 6772 17382
rect 6796 17380 6852 17382
rect 6556 16346 6612 16348
rect 6636 16346 6692 16348
rect 6716 16346 6772 16348
rect 6796 16346 6852 16348
rect 6556 16294 6602 16346
rect 6602 16294 6612 16346
rect 6636 16294 6666 16346
rect 6666 16294 6678 16346
rect 6678 16294 6692 16346
rect 6716 16294 6730 16346
rect 6730 16294 6742 16346
rect 6742 16294 6772 16346
rect 6796 16294 6806 16346
rect 6806 16294 6852 16346
rect 6556 16292 6612 16294
rect 6636 16292 6692 16294
rect 6716 16292 6772 16294
rect 6796 16292 6852 16294
rect 6556 15258 6612 15260
rect 6636 15258 6692 15260
rect 6716 15258 6772 15260
rect 6796 15258 6852 15260
rect 6556 15206 6602 15258
rect 6602 15206 6612 15258
rect 6636 15206 6666 15258
rect 6666 15206 6678 15258
rect 6678 15206 6692 15258
rect 6716 15206 6730 15258
rect 6730 15206 6742 15258
rect 6742 15206 6772 15258
rect 6796 15206 6806 15258
rect 6806 15206 6852 15258
rect 6556 15204 6612 15206
rect 6636 15204 6692 15206
rect 6716 15204 6772 15206
rect 6796 15204 6852 15206
rect 6556 14170 6612 14172
rect 6636 14170 6692 14172
rect 6716 14170 6772 14172
rect 6796 14170 6852 14172
rect 6556 14118 6602 14170
rect 6602 14118 6612 14170
rect 6636 14118 6666 14170
rect 6666 14118 6678 14170
rect 6678 14118 6692 14170
rect 6716 14118 6730 14170
rect 6730 14118 6742 14170
rect 6742 14118 6772 14170
rect 6796 14118 6806 14170
rect 6806 14118 6852 14170
rect 6556 14116 6612 14118
rect 6636 14116 6692 14118
rect 6716 14116 6772 14118
rect 6796 14116 6852 14118
rect 7216 16890 7272 16892
rect 7296 16890 7352 16892
rect 7376 16890 7432 16892
rect 7456 16890 7512 16892
rect 7216 16838 7262 16890
rect 7262 16838 7272 16890
rect 7296 16838 7326 16890
rect 7326 16838 7338 16890
rect 7338 16838 7352 16890
rect 7376 16838 7390 16890
rect 7390 16838 7402 16890
rect 7402 16838 7432 16890
rect 7456 16838 7466 16890
rect 7466 16838 7512 16890
rect 7216 16836 7272 16838
rect 7296 16836 7352 16838
rect 7376 16836 7432 16838
rect 7456 16836 7512 16838
rect 7216 15802 7272 15804
rect 7296 15802 7352 15804
rect 7376 15802 7432 15804
rect 7456 15802 7512 15804
rect 7216 15750 7262 15802
rect 7262 15750 7272 15802
rect 7296 15750 7326 15802
rect 7326 15750 7338 15802
rect 7338 15750 7352 15802
rect 7376 15750 7390 15802
rect 7390 15750 7402 15802
rect 7402 15750 7432 15802
rect 7456 15750 7466 15802
rect 7466 15750 7512 15802
rect 7216 15748 7272 15750
rect 7296 15748 7352 15750
rect 7376 15748 7432 15750
rect 7456 15748 7512 15750
rect 7746 17720 7802 17776
rect 7216 14714 7272 14716
rect 7296 14714 7352 14716
rect 7376 14714 7432 14716
rect 7456 14714 7512 14716
rect 7216 14662 7262 14714
rect 7262 14662 7272 14714
rect 7296 14662 7326 14714
rect 7326 14662 7338 14714
rect 7338 14662 7352 14714
rect 7376 14662 7390 14714
rect 7390 14662 7402 14714
rect 7402 14662 7432 14714
rect 7456 14662 7466 14714
rect 7466 14662 7512 14714
rect 7216 14660 7272 14662
rect 7296 14660 7352 14662
rect 7376 14660 7432 14662
rect 7456 14660 7512 14662
rect 7216 13626 7272 13628
rect 7296 13626 7352 13628
rect 7376 13626 7432 13628
rect 7456 13626 7512 13628
rect 7216 13574 7262 13626
rect 7262 13574 7272 13626
rect 7296 13574 7326 13626
rect 7326 13574 7338 13626
rect 7338 13574 7352 13626
rect 7376 13574 7390 13626
rect 7390 13574 7402 13626
rect 7402 13574 7432 13626
rect 7456 13574 7466 13626
rect 7466 13574 7512 13626
rect 7216 13572 7272 13574
rect 7296 13572 7352 13574
rect 7376 13572 7432 13574
rect 7456 13572 7512 13574
rect 6556 13082 6612 13084
rect 6636 13082 6692 13084
rect 6716 13082 6772 13084
rect 6796 13082 6852 13084
rect 6556 13030 6602 13082
rect 6602 13030 6612 13082
rect 6636 13030 6666 13082
rect 6666 13030 6678 13082
rect 6678 13030 6692 13082
rect 6716 13030 6730 13082
rect 6730 13030 6742 13082
rect 6742 13030 6772 13082
rect 6796 13030 6806 13082
rect 6806 13030 6852 13082
rect 6556 13028 6612 13030
rect 6636 13028 6692 13030
rect 6716 13028 6772 13030
rect 6796 13028 6852 13030
rect 7216 12538 7272 12540
rect 7296 12538 7352 12540
rect 7376 12538 7432 12540
rect 7456 12538 7512 12540
rect 7216 12486 7262 12538
rect 7262 12486 7272 12538
rect 7296 12486 7326 12538
rect 7326 12486 7338 12538
rect 7338 12486 7352 12538
rect 7376 12486 7390 12538
rect 7390 12486 7402 12538
rect 7402 12486 7432 12538
rect 7456 12486 7466 12538
rect 7466 12486 7512 12538
rect 7216 12484 7272 12486
rect 7296 12484 7352 12486
rect 7376 12484 7432 12486
rect 7456 12484 7512 12486
rect 6556 11994 6612 11996
rect 6636 11994 6692 11996
rect 6716 11994 6772 11996
rect 6796 11994 6852 11996
rect 6556 11942 6602 11994
rect 6602 11942 6612 11994
rect 6636 11942 6666 11994
rect 6666 11942 6678 11994
rect 6678 11942 6692 11994
rect 6716 11942 6730 11994
rect 6730 11942 6742 11994
rect 6742 11942 6772 11994
rect 6796 11942 6806 11994
rect 6806 11942 6852 11994
rect 6556 11940 6612 11942
rect 6636 11940 6692 11942
rect 6716 11940 6772 11942
rect 6796 11940 6852 11942
rect 7216 11450 7272 11452
rect 7296 11450 7352 11452
rect 7376 11450 7432 11452
rect 7456 11450 7512 11452
rect 7216 11398 7262 11450
rect 7262 11398 7272 11450
rect 7296 11398 7326 11450
rect 7326 11398 7338 11450
rect 7338 11398 7352 11450
rect 7376 11398 7390 11450
rect 7390 11398 7402 11450
rect 7402 11398 7432 11450
rect 7456 11398 7466 11450
rect 7466 11398 7512 11450
rect 7216 11396 7272 11398
rect 7296 11396 7352 11398
rect 7376 11396 7432 11398
rect 7456 11396 7512 11398
rect 6556 10906 6612 10908
rect 6636 10906 6692 10908
rect 6716 10906 6772 10908
rect 6796 10906 6852 10908
rect 6556 10854 6602 10906
rect 6602 10854 6612 10906
rect 6636 10854 6666 10906
rect 6666 10854 6678 10906
rect 6678 10854 6692 10906
rect 6716 10854 6730 10906
rect 6730 10854 6742 10906
rect 6742 10854 6772 10906
rect 6796 10854 6806 10906
rect 6806 10854 6852 10906
rect 6556 10852 6612 10854
rect 6636 10852 6692 10854
rect 6716 10852 6772 10854
rect 6796 10852 6852 10854
rect 4066 6160 4122 6216
rect 3054 5480 3110 5536
rect 1306 4120 1362 4176
rect 1306 2760 1362 2816
rect 3054 1400 3110 1456
rect 6556 9818 6612 9820
rect 6636 9818 6692 9820
rect 6716 9818 6772 9820
rect 6796 9818 6852 9820
rect 6556 9766 6602 9818
rect 6602 9766 6612 9818
rect 6636 9766 6666 9818
rect 6666 9766 6678 9818
rect 6678 9766 6692 9818
rect 6716 9766 6730 9818
rect 6730 9766 6742 9818
rect 6742 9766 6772 9818
rect 6796 9766 6806 9818
rect 6806 9766 6852 9818
rect 6556 9764 6612 9766
rect 6636 9764 6692 9766
rect 6716 9764 6772 9766
rect 6796 9764 6852 9766
rect 7216 10362 7272 10364
rect 7296 10362 7352 10364
rect 7376 10362 7432 10364
rect 7456 10362 7512 10364
rect 7216 10310 7262 10362
rect 7262 10310 7272 10362
rect 7296 10310 7326 10362
rect 7326 10310 7338 10362
rect 7338 10310 7352 10362
rect 7376 10310 7390 10362
rect 7390 10310 7402 10362
rect 7402 10310 7432 10362
rect 7456 10310 7466 10362
rect 7466 10310 7512 10362
rect 7216 10308 7272 10310
rect 7296 10308 7352 10310
rect 7376 10308 7432 10310
rect 7456 10308 7512 10310
rect 8666 18264 8722 18320
rect 10046 23604 10048 23624
rect 10048 23604 10100 23624
rect 10100 23604 10102 23624
rect 10046 23568 10102 23604
rect 9862 21548 9918 21584
rect 9862 21528 9864 21548
rect 9864 21528 9916 21548
rect 9916 21528 9918 21548
rect 9034 19796 9036 19816
rect 9036 19796 9088 19816
rect 9088 19796 9090 19816
rect 9034 19760 9090 19796
rect 10046 20848 10102 20904
rect 13082 29144 13138 29200
rect 11610 24792 11666 24848
rect 14445 32666 14501 32668
rect 14525 32666 14581 32668
rect 14605 32666 14661 32668
rect 14685 32666 14741 32668
rect 14445 32614 14491 32666
rect 14491 32614 14501 32666
rect 14525 32614 14555 32666
rect 14555 32614 14567 32666
rect 14567 32614 14581 32666
rect 14605 32614 14619 32666
rect 14619 32614 14631 32666
rect 14631 32614 14661 32666
rect 14685 32614 14695 32666
rect 14695 32614 14741 32666
rect 14445 32612 14501 32614
rect 14525 32612 14581 32614
rect 14605 32612 14661 32614
rect 14685 32612 14741 32614
rect 15014 32408 15070 32464
rect 15566 32816 15622 32872
rect 11610 23160 11666 23216
rect 10506 20304 10562 20360
rect 10874 20032 10930 20088
rect 11058 19896 11114 19952
rect 10690 19488 10746 19544
rect 9954 18944 10010 19000
rect 7216 9274 7272 9276
rect 7296 9274 7352 9276
rect 7376 9274 7432 9276
rect 7456 9274 7512 9276
rect 7216 9222 7262 9274
rect 7262 9222 7272 9274
rect 7296 9222 7326 9274
rect 7326 9222 7338 9274
rect 7338 9222 7352 9274
rect 7376 9222 7390 9274
rect 7390 9222 7402 9274
rect 7402 9222 7432 9274
rect 7456 9222 7466 9274
rect 7466 9222 7512 9274
rect 7216 9220 7272 9222
rect 7296 9220 7352 9222
rect 7376 9220 7432 9222
rect 7456 9220 7512 9222
rect 6556 8730 6612 8732
rect 6636 8730 6692 8732
rect 6716 8730 6772 8732
rect 6796 8730 6852 8732
rect 6556 8678 6602 8730
rect 6602 8678 6612 8730
rect 6636 8678 6666 8730
rect 6666 8678 6678 8730
rect 6678 8678 6692 8730
rect 6716 8678 6730 8730
rect 6730 8678 6742 8730
rect 6742 8678 6772 8730
rect 6796 8678 6806 8730
rect 6806 8678 6852 8730
rect 6556 8676 6612 8678
rect 6636 8676 6692 8678
rect 6716 8676 6772 8678
rect 6796 8676 6852 8678
rect 7216 8186 7272 8188
rect 7296 8186 7352 8188
rect 7376 8186 7432 8188
rect 7456 8186 7512 8188
rect 7216 8134 7262 8186
rect 7262 8134 7272 8186
rect 7296 8134 7326 8186
rect 7326 8134 7338 8186
rect 7338 8134 7352 8186
rect 7376 8134 7390 8186
rect 7390 8134 7402 8186
rect 7402 8134 7432 8186
rect 7456 8134 7466 8186
rect 7466 8134 7512 8186
rect 7216 8132 7272 8134
rect 7296 8132 7352 8134
rect 7376 8132 7432 8134
rect 7456 8132 7512 8134
rect 6556 7642 6612 7644
rect 6636 7642 6692 7644
rect 6716 7642 6772 7644
rect 6796 7642 6852 7644
rect 6556 7590 6602 7642
rect 6602 7590 6612 7642
rect 6636 7590 6666 7642
rect 6666 7590 6678 7642
rect 6678 7590 6692 7642
rect 6716 7590 6730 7642
rect 6730 7590 6742 7642
rect 6742 7590 6772 7642
rect 6796 7590 6806 7642
rect 6806 7590 6852 7642
rect 6556 7588 6612 7590
rect 6636 7588 6692 7590
rect 6716 7588 6772 7590
rect 6796 7588 6852 7590
rect 7216 7098 7272 7100
rect 7296 7098 7352 7100
rect 7376 7098 7432 7100
rect 7456 7098 7512 7100
rect 7216 7046 7262 7098
rect 7262 7046 7272 7098
rect 7296 7046 7326 7098
rect 7326 7046 7338 7098
rect 7338 7046 7352 7098
rect 7376 7046 7390 7098
rect 7390 7046 7402 7098
rect 7402 7046 7432 7098
rect 7456 7046 7466 7098
rect 7466 7046 7512 7098
rect 7216 7044 7272 7046
rect 7296 7044 7352 7046
rect 7376 7044 7432 7046
rect 7456 7044 7512 7046
rect 6556 6554 6612 6556
rect 6636 6554 6692 6556
rect 6716 6554 6772 6556
rect 6796 6554 6852 6556
rect 6556 6502 6602 6554
rect 6602 6502 6612 6554
rect 6636 6502 6666 6554
rect 6666 6502 6678 6554
rect 6678 6502 6692 6554
rect 6716 6502 6730 6554
rect 6730 6502 6742 6554
rect 6742 6502 6772 6554
rect 6796 6502 6806 6554
rect 6806 6502 6852 6554
rect 6556 6500 6612 6502
rect 6636 6500 6692 6502
rect 6716 6500 6772 6502
rect 6796 6500 6852 6502
rect 7216 6010 7272 6012
rect 7296 6010 7352 6012
rect 7376 6010 7432 6012
rect 7456 6010 7512 6012
rect 7216 5958 7262 6010
rect 7262 5958 7272 6010
rect 7296 5958 7326 6010
rect 7326 5958 7338 6010
rect 7338 5958 7352 6010
rect 7376 5958 7390 6010
rect 7390 5958 7402 6010
rect 7402 5958 7432 6010
rect 7456 5958 7466 6010
rect 7466 5958 7512 6010
rect 7216 5956 7272 5958
rect 7296 5956 7352 5958
rect 7376 5956 7432 5958
rect 7456 5956 7512 5958
rect 6556 5466 6612 5468
rect 6636 5466 6692 5468
rect 6716 5466 6772 5468
rect 6796 5466 6852 5468
rect 6556 5414 6602 5466
rect 6602 5414 6612 5466
rect 6636 5414 6666 5466
rect 6666 5414 6678 5466
rect 6678 5414 6692 5466
rect 6716 5414 6730 5466
rect 6730 5414 6742 5466
rect 6742 5414 6772 5466
rect 6796 5414 6806 5466
rect 6806 5414 6852 5466
rect 6556 5412 6612 5414
rect 6636 5412 6692 5414
rect 6716 5412 6772 5414
rect 6796 5412 6852 5414
rect 7216 4922 7272 4924
rect 7296 4922 7352 4924
rect 7376 4922 7432 4924
rect 7456 4922 7512 4924
rect 7216 4870 7262 4922
rect 7262 4870 7272 4922
rect 7296 4870 7326 4922
rect 7326 4870 7338 4922
rect 7338 4870 7352 4922
rect 7376 4870 7390 4922
rect 7390 4870 7402 4922
rect 7402 4870 7432 4922
rect 7456 4870 7466 4922
rect 7466 4870 7512 4922
rect 7216 4868 7272 4870
rect 7296 4868 7352 4870
rect 7376 4868 7432 4870
rect 7456 4868 7512 4870
rect 6556 4378 6612 4380
rect 6636 4378 6692 4380
rect 6716 4378 6772 4380
rect 6796 4378 6852 4380
rect 6556 4326 6602 4378
rect 6602 4326 6612 4378
rect 6636 4326 6666 4378
rect 6666 4326 6678 4378
rect 6678 4326 6692 4378
rect 6716 4326 6730 4378
rect 6730 4326 6742 4378
rect 6742 4326 6772 4378
rect 6796 4326 6806 4378
rect 6806 4326 6852 4378
rect 6556 4324 6612 4326
rect 6636 4324 6692 4326
rect 6716 4324 6772 4326
rect 6796 4324 6852 4326
rect 7216 3834 7272 3836
rect 7296 3834 7352 3836
rect 7376 3834 7432 3836
rect 7456 3834 7512 3836
rect 7216 3782 7262 3834
rect 7262 3782 7272 3834
rect 7296 3782 7326 3834
rect 7326 3782 7338 3834
rect 7338 3782 7352 3834
rect 7376 3782 7390 3834
rect 7390 3782 7402 3834
rect 7402 3782 7432 3834
rect 7456 3782 7466 3834
rect 7466 3782 7512 3834
rect 7216 3780 7272 3782
rect 7296 3780 7352 3782
rect 7376 3780 7432 3782
rect 7456 3780 7512 3782
rect 6556 3290 6612 3292
rect 6636 3290 6692 3292
rect 6716 3290 6772 3292
rect 6796 3290 6852 3292
rect 6556 3238 6602 3290
rect 6602 3238 6612 3290
rect 6636 3238 6666 3290
rect 6666 3238 6678 3290
rect 6678 3238 6692 3290
rect 6716 3238 6730 3290
rect 6730 3238 6742 3290
rect 6742 3238 6772 3290
rect 6796 3238 6806 3290
rect 6806 3238 6852 3290
rect 6556 3236 6612 3238
rect 6636 3236 6692 3238
rect 6716 3236 6772 3238
rect 6796 3236 6852 3238
rect 5722 3052 5778 3088
rect 5722 3032 5724 3052
rect 5724 3032 5776 3052
rect 5776 3032 5778 3052
rect 7216 2746 7272 2748
rect 7296 2746 7352 2748
rect 7376 2746 7432 2748
rect 7456 2746 7512 2748
rect 7216 2694 7262 2746
rect 7262 2694 7272 2746
rect 7296 2694 7326 2746
rect 7326 2694 7338 2746
rect 7338 2694 7352 2746
rect 7376 2694 7390 2746
rect 7390 2694 7402 2746
rect 7402 2694 7432 2746
rect 7456 2694 7466 2746
rect 7466 2694 7512 2746
rect 7216 2692 7272 2694
rect 7296 2692 7352 2694
rect 7376 2692 7432 2694
rect 7456 2692 7512 2694
rect 12622 23568 12678 23624
rect 11702 21664 11758 21720
rect 11518 20884 11520 20904
rect 11520 20884 11572 20904
rect 11572 20884 11574 20904
rect 11518 20848 11574 20884
rect 12714 20984 12770 21040
rect 11886 20440 11942 20496
rect 11334 19760 11390 19816
rect 11242 19488 11298 19544
rect 8666 7792 8722 7848
rect 9218 7948 9274 7984
rect 9218 7928 9220 7948
rect 9220 7928 9272 7948
rect 9272 7928 9274 7948
rect 12806 19216 12862 19272
rect 12806 17060 12862 17096
rect 12806 17040 12808 17060
rect 12808 17040 12860 17060
rect 12860 17040 12862 17060
rect 14002 26968 14058 27024
rect 15105 32122 15161 32124
rect 15185 32122 15241 32124
rect 15265 32122 15321 32124
rect 15345 32122 15401 32124
rect 15105 32070 15151 32122
rect 15151 32070 15161 32122
rect 15185 32070 15215 32122
rect 15215 32070 15227 32122
rect 15227 32070 15241 32122
rect 15265 32070 15279 32122
rect 15279 32070 15291 32122
rect 15291 32070 15321 32122
rect 15345 32070 15355 32122
rect 15355 32070 15401 32122
rect 15105 32068 15161 32070
rect 15185 32068 15241 32070
rect 15265 32068 15321 32070
rect 15345 32068 15401 32070
rect 14445 31578 14501 31580
rect 14525 31578 14581 31580
rect 14605 31578 14661 31580
rect 14685 31578 14741 31580
rect 14445 31526 14491 31578
rect 14491 31526 14501 31578
rect 14525 31526 14555 31578
rect 14555 31526 14567 31578
rect 14567 31526 14581 31578
rect 14605 31526 14619 31578
rect 14619 31526 14631 31578
rect 14631 31526 14661 31578
rect 14685 31526 14695 31578
rect 14695 31526 14741 31578
rect 14445 31524 14501 31526
rect 14525 31524 14581 31526
rect 14605 31524 14661 31526
rect 14685 31524 14741 31526
rect 14445 30490 14501 30492
rect 14525 30490 14581 30492
rect 14605 30490 14661 30492
rect 14685 30490 14741 30492
rect 14445 30438 14491 30490
rect 14491 30438 14501 30490
rect 14525 30438 14555 30490
rect 14555 30438 14567 30490
rect 14567 30438 14581 30490
rect 14605 30438 14619 30490
rect 14619 30438 14631 30490
rect 14631 30438 14661 30490
rect 14685 30438 14695 30490
rect 14695 30438 14741 30490
rect 14445 30436 14501 30438
rect 14525 30436 14581 30438
rect 14605 30436 14661 30438
rect 14685 30436 14741 30438
rect 14445 29402 14501 29404
rect 14525 29402 14581 29404
rect 14605 29402 14661 29404
rect 14685 29402 14741 29404
rect 14445 29350 14491 29402
rect 14491 29350 14501 29402
rect 14525 29350 14555 29402
rect 14555 29350 14567 29402
rect 14567 29350 14581 29402
rect 14605 29350 14619 29402
rect 14619 29350 14631 29402
rect 14631 29350 14661 29402
rect 14685 29350 14695 29402
rect 14695 29350 14741 29402
rect 14445 29348 14501 29350
rect 14525 29348 14581 29350
rect 14605 29348 14661 29350
rect 14685 29348 14741 29350
rect 15105 31034 15161 31036
rect 15185 31034 15241 31036
rect 15265 31034 15321 31036
rect 15345 31034 15401 31036
rect 15105 30982 15151 31034
rect 15151 30982 15161 31034
rect 15185 30982 15215 31034
rect 15215 30982 15227 31034
rect 15227 30982 15241 31034
rect 15265 30982 15279 31034
rect 15279 30982 15291 31034
rect 15291 30982 15321 31034
rect 15345 30982 15355 31034
rect 15355 30982 15401 31034
rect 15105 30980 15161 30982
rect 15185 30980 15241 30982
rect 15265 30980 15321 30982
rect 15345 30980 15401 30982
rect 15105 29946 15161 29948
rect 15185 29946 15241 29948
rect 15265 29946 15321 29948
rect 15345 29946 15401 29948
rect 15105 29894 15151 29946
rect 15151 29894 15161 29946
rect 15185 29894 15215 29946
rect 15215 29894 15227 29946
rect 15227 29894 15241 29946
rect 15265 29894 15279 29946
rect 15279 29894 15291 29946
rect 15291 29894 15321 29946
rect 15345 29894 15355 29946
rect 15355 29894 15401 29946
rect 15105 29892 15161 29894
rect 15185 29892 15241 29894
rect 15265 29892 15321 29894
rect 15345 29892 15401 29894
rect 14445 28314 14501 28316
rect 14525 28314 14581 28316
rect 14605 28314 14661 28316
rect 14685 28314 14741 28316
rect 14445 28262 14491 28314
rect 14491 28262 14501 28314
rect 14525 28262 14555 28314
rect 14555 28262 14567 28314
rect 14567 28262 14581 28314
rect 14605 28262 14619 28314
rect 14619 28262 14631 28314
rect 14631 28262 14661 28314
rect 14685 28262 14695 28314
rect 14695 28262 14741 28314
rect 14445 28260 14501 28262
rect 14525 28260 14581 28262
rect 14605 28260 14661 28262
rect 14685 28260 14741 28262
rect 14445 27226 14501 27228
rect 14525 27226 14581 27228
rect 14605 27226 14661 27228
rect 14685 27226 14741 27228
rect 14445 27174 14491 27226
rect 14491 27174 14501 27226
rect 14525 27174 14555 27226
rect 14555 27174 14567 27226
rect 14567 27174 14581 27226
rect 14605 27174 14619 27226
rect 14619 27174 14631 27226
rect 14631 27174 14661 27226
rect 14685 27174 14695 27226
rect 14695 27174 14741 27226
rect 14445 27172 14501 27174
rect 14525 27172 14581 27174
rect 14605 27172 14661 27174
rect 14685 27172 14741 27174
rect 15105 28858 15161 28860
rect 15185 28858 15241 28860
rect 15265 28858 15321 28860
rect 15345 28858 15401 28860
rect 15105 28806 15151 28858
rect 15151 28806 15161 28858
rect 15185 28806 15215 28858
rect 15215 28806 15227 28858
rect 15227 28806 15241 28858
rect 15265 28806 15279 28858
rect 15279 28806 15291 28858
rect 15291 28806 15321 28858
rect 15345 28806 15355 28858
rect 15355 28806 15401 28858
rect 15105 28804 15161 28806
rect 15185 28804 15241 28806
rect 15265 28804 15321 28806
rect 15345 28804 15401 28806
rect 15105 27770 15161 27772
rect 15185 27770 15241 27772
rect 15265 27770 15321 27772
rect 15345 27770 15401 27772
rect 15105 27718 15151 27770
rect 15151 27718 15161 27770
rect 15185 27718 15215 27770
rect 15215 27718 15227 27770
rect 15227 27718 15241 27770
rect 15265 27718 15279 27770
rect 15279 27718 15291 27770
rect 15291 27718 15321 27770
rect 15345 27718 15355 27770
rect 15355 27718 15401 27770
rect 15105 27716 15161 27718
rect 15185 27716 15241 27718
rect 15265 27716 15321 27718
rect 15345 27716 15401 27718
rect 15105 26682 15161 26684
rect 15185 26682 15241 26684
rect 15265 26682 15321 26684
rect 15345 26682 15401 26684
rect 15105 26630 15151 26682
rect 15151 26630 15161 26682
rect 15185 26630 15215 26682
rect 15215 26630 15227 26682
rect 15227 26630 15241 26682
rect 15265 26630 15279 26682
rect 15279 26630 15291 26682
rect 15291 26630 15321 26682
rect 15345 26630 15355 26682
rect 15355 26630 15401 26682
rect 15105 26628 15161 26630
rect 15185 26628 15241 26630
rect 15265 26628 15321 26630
rect 15345 26628 15401 26630
rect 14445 26138 14501 26140
rect 14525 26138 14581 26140
rect 14605 26138 14661 26140
rect 14685 26138 14741 26140
rect 14445 26086 14491 26138
rect 14491 26086 14501 26138
rect 14525 26086 14555 26138
rect 14555 26086 14567 26138
rect 14567 26086 14581 26138
rect 14605 26086 14619 26138
rect 14619 26086 14631 26138
rect 14631 26086 14661 26138
rect 14685 26086 14695 26138
rect 14695 26086 14741 26138
rect 14445 26084 14501 26086
rect 14525 26084 14581 26086
rect 14605 26084 14661 26086
rect 14685 26084 14741 26086
rect 15105 25594 15161 25596
rect 15185 25594 15241 25596
rect 15265 25594 15321 25596
rect 15345 25594 15401 25596
rect 15105 25542 15151 25594
rect 15151 25542 15161 25594
rect 15185 25542 15215 25594
rect 15215 25542 15227 25594
rect 15227 25542 15241 25594
rect 15265 25542 15279 25594
rect 15279 25542 15291 25594
rect 15291 25542 15321 25594
rect 15345 25542 15355 25594
rect 15355 25542 15401 25594
rect 15105 25540 15161 25542
rect 15185 25540 15241 25542
rect 15265 25540 15321 25542
rect 15345 25540 15401 25542
rect 14445 25050 14501 25052
rect 14525 25050 14581 25052
rect 14605 25050 14661 25052
rect 14685 25050 14741 25052
rect 14445 24998 14491 25050
rect 14491 24998 14501 25050
rect 14525 24998 14555 25050
rect 14555 24998 14567 25050
rect 14567 24998 14581 25050
rect 14605 24998 14619 25050
rect 14619 24998 14631 25050
rect 14631 24998 14661 25050
rect 14685 24998 14695 25050
rect 14695 24998 14741 25050
rect 14445 24996 14501 24998
rect 14525 24996 14581 24998
rect 14605 24996 14661 24998
rect 14685 24996 14741 24998
rect 14445 23962 14501 23964
rect 14525 23962 14581 23964
rect 14605 23962 14661 23964
rect 14685 23962 14741 23964
rect 14445 23910 14491 23962
rect 14491 23910 14501 23962
rect 14525 23910 14555 23962
rect 14555 23910 14567 23962
rect 14567 23910 14581 23962
rect 14605 23910 14619 23962
rect 14619 23910 14631 23962
rect 14631 23910 14661 23962
rect 14685 23910 14695 23962
rect 14695 23910 14741 23962
rect 14445 23908 14501 23910
rect 14525 23908 14581 23910
rect 14605 23908 14661 23910
rect 14685 23908 14741 23910
rect 13818 20032 13874 20088
rect 13634 17584 13690 17640
rect 12162 11056 12218 11112
rect 14445 22874 14501 22876
rect 14525 22874 14581 22876
rect 14605 22874 14661 22876
rect 14685 22874 14741 22876
rect 14445 22822 14491 22874
rect 14491 22822 14501 22874
rect 14525 22822 14555 22874
rect 14555 22822 14567 22874
rect 14567 22822 14581 22874
rect 14605 22822 14619 22874
rect 14619 22822 14631 22874
rect 14631 22822 14661 22874
rect 14685 22822 14695 22874
rect 14695 22822 14741 22874
rect 14445 22820 14501 22822
rect 14525 22820 14581 22822
rect 14605 22820 14661 22822
rect 14685 22820 14741 22822
rect 15105 24506 15161 24508
rect 15185 24506 15241 24508
rect 15265 24506 15321 24508
rect 15345 24506 15401 24508
rect 15105 24454 15151 24506
rect 15151 24454 15161 24506
rect 15185 24454 15215 24506
rect 15215 24454 15227 24506
rect 15227 24454 15241 24506
rect 15265 24454 15279 24506
rect 15279 24454 15291 24506
rect 15291 24454 15321 24506
rect 15345 24454 15355 24506
rect 15355 24454 15401 24506
rect 15105 24452 15161 24454
rect 15185 24452 15241 24454
rect 15265 24452 15321 24454
rect 15345 24452 15401 24454
rect 15105 23418 15161 23420
rect 15185 23418 15241 23420
rect 15265 23418 15321 23420
rect 15345 23418 15401 23420
rect 15105 23366 15151 23418
rect 15151 23366 15161 23418
rect 15185 23366 15215 23418
rect 15215 23366 15227 23418
rect 15227 23366 15241 23418
rect 15265 23366 15279 23418
rect 15279 23366 15291 23418
rect 15291 23366 15321 23418
rect 15345 23366 15355 23418
rect 15355 23366 15401 23418
rect 15105 23364 15161 23366
rect 15185 23364 15241 23366
rect 15265 23364 15321 23366
rect 15345 23364 15401 23366
rect 14445 21786 14501 21788
rect 14525 21786 14581 21788
rect 14605 21786 14661 21788
rect 14685 21786 14741 21788
rect 14445 21734 14491 21786
rect 14491 21734 14501 21786
rect 14525 21734 14555 21786
rect 14555 21734 14567 21786
rect 14567 21734 14581 21786
rect 14605 21734 14619 21786
rect 14619 21734 14631 21786
rect 14631 21734 14661 21786
rect 14685 21734 14695 21786
rect 14695 21734 14741 21786
rect 14445 21732 14501 21734
rect 14525 21732 14581 21734
rect 14605 21732 14661 21734
rect 14685 21732 14741 21734
rect 14445 20698 14501 20700
rect 14525 20698 14581 20700
rect 14605 20698 14661 20700
rect 14685 20698 14741 20700
rect 14445 20646 14491 20698
rect 14491 20646 14501 20698
rect 14525 20646 14555 20698
rect 14555 20646 14567 20698
rect 14567 20646 14581 20698
rect 14605 20646 14619 20698
rect 14619 20646 14631 20698
rect 14631 20646 14661 20698
rect 14685 20646 14695 20698
rect 14695 20646 14741 20698
rect 14445 20644 14501 20646
rect 14525 20644 14581 20646
rect 14605 20644 14661 20646
rect 14685 20644 14741 20646
rect 15105 22330 15161 22332
rect 15185 22330 15241 22332
rect 15265 22330 15321 22332
rect 15345 22330 15401 22332
rect 15105 22278 15151 22330
rect 15151 22278 15161 22330
rect 15185 22278 15215 22330
rect 15215 22278 15227 22330
rect 15227 22278 15241 22330
rect 15265 22278 15279 22330
rect 15279 22278 15291 22330
rect 15291 22278 15321 22330
rect 15345 22278 15355 22330
rect 15355 22278 15401 22330
rect 15105 22276 15161 22278
rect 15185 22276 15241 22278
rect 15265 22276 15321 22278
rect 15345 22276 15401 22278
rect 14186 19932 14188 19952
rect 14188 19932 14240 19952
rect 14240 19932 14242 19952
rect 14186 19896 14242 19932
rect 14445 19610 14501 19612
rect 14525 19610 14581 19612
rect 14605 19610 14661 19612
rect 14685 19610 14741 19612
rect 14445 19558 14491 19610
rect 14491 19558 14501 19610
rect 14525 19558 14555 19610
rect 14555 19558 14567 19610
rect 14567 19558 14581 19610
rect 14605 19558 14619 19610
rect 14619 19558 14631 19610
rect 14631 19558 14661 19610
rect 14685 19558 14695 19610
rect 14695 19558 14741 19610
rect 14445 19556 14501 19558
rect 14525 19556 14581 19558
rect 14605 19556 14661 19558
rect 14685 19556 14741 19558
rect 14370 19216 14426 19272
rect 14445 18522 14501 18524
rect 14525 18522 14581 18524
rect 14605 18522 14661 18524
rect 14685 18522 14741 18524
rect 14445 18470 14491 18522
rect 14491 18470 14501 18522
rect 14525 18470 14555 18522
rect 14555 18470 14567 18522
rect 14567 18470 14581 18522
rect 14605 18470 14619 18522
rect 14619 18470 14631 18522
rect 14631 18470 14661 18522
rect 14685 18470 14695 18522
rect 14695 18470 14741 18522
rect 14445 18468 14501 18470
rect 14525 18468 14581 18470
rect 14605 18468 14661 18470
rect 14685 18468 14741 18470
rect 14922 18264 14978 18320
rect 14278 18128 14334 18184
rect 14445 17434 14501 17436
rect 14525 17434 14581 17436
rect 14605 17434 14661 17436
rect 14685 17434 14741 17436
rect 14445 17382 14491 17434
rect 14491 17382 14501 17434
rect 14525 17382 14555 17434
rect 14555 17382 14567 17434
rect 14567 17382 14581 17434
rect 14605 17382 14619 17434
rect 14619 17382 14631 17434
rect 14631 17382 14661 17434
rect 14685 17382 14695 17434
rect 14695 17382 14741 17434
rect 14445 17380 14501 17382
rect 14525 17380 14581 17382
rect 14605 17380 14661 17382
rect 14685 17380 14741 17382
rect 15105 21242 15161 21244
rect 15185 21242 15241 21244
rect 15265 21242 15321 21244
rect 15345 21242 15401 21244
rect 15105 21190 15151 21242
rect 15151 21190 15161 21242
rect 15185 21190 15215 21242
rect 15215 21190 15227 21242
rect 15227 21190 15241 21242
rect 15265 21190 15279 21242
rect 15279 21190 15291 21242
rect 15291 21190 15321 21242
rect 15345 21190 15355 21242
rect 15355 21190 15401 21242
rect 15105 21188 15161 21190
rect 15185 21188 15241 21190
rect 15265 21188 15321 21190
rect 15345 21188 15401 21190
rect 15934 26968 15990 27024
rect 15566 23704 15622 23760
rect 15105 20154 15161 20156
rect 15185 20154 15241 20156
rect 15265 20154 15321 20156
rect 15345 20154 15401 20156
rect 15105 20102 15151 20154
rect 15151 20102 15161 20154
rect 15185 20102 15215 20154
rect 15215 20102 15227 20154
rect 15227 20102 15241 20154
rect 15265 20102 15279 20154
rect 15279 20102 15291 20154
rect 15291 20102 15321 20154
rect 15345 20102 15355 20154
rect 15355 20102 15401 20154
rect 15105 20100 15161 20102
rect 15185 20100 15241 20102
rect 15265 20100 15321 20102
rect 15345 20100 15401 20102
rect 15105 19066 15161 19068
rect 15185 19066 15241 19068
rect 15265 19066 15321 19068
rect 15345 19066 15401 19068
rect 15105 19014 15151 19066
rect 15151 19014 15161 19066
rect 15185 19014 15215 19066
rect 15215 19014 15227 19066
rect 15227 19014 15241 19066
rect 15265 19014 15279 19066
rect 15279 19014 15291 19066
rect 15291 19014 15321 19066
rect 15345 19014 15355 19066
rect 15355 19014 15401 19066
rect 15105 19012 15161 19014
rect 15185 19012 15241 19014
rect 15265 19012 15321 19014
rect 15345 19012 15401 19014
rect 15105 17978 15161 17980
rect 15185 17978 15241 17980
rect 15265 17978 15321 17980
rect 15345 17978 15401 17980
rect 15105 17926 15151 17978
rect 15151 17926 15161 17978
rect 15185 17926 15215 17978
rect 15215 17926 15227 17978
rect 15227 17926 15241 17978
rect 15265 17926 15279 17978
rect 15279 17926 15291 17978
rect 15291 17926 15321 17978
rect 15345 17926 15355 17978
rect 15355 17926 15401 17978
rect 15105 17924 15161 17926
rect 15185 17924 15241 17926
rect 15265 17924 15321 17926
rect 15345 17924 15401 17926
rect 15105 16890 15161 16892
rect 15185 16890 15241 16892
rect 15265 16890 15321 16892
rect 15345 16890 15401 16892
rect 15105 16838 15151 16890
rect 15151 16838 15161 16890
rect 15185 16838 15215 16890
rect 15215 16838 15227 16890
rect 15227 16838 15241 16890
rect 15265 16838 15279 16890
rect 15279 16838 15291 16890
rect 15291 16838 15321 16890
rect 15345 16838 15355 16890
rect 15355 16838 15401 16890
rect 15105 16836 15161 16838
rect 15185 16836 15241 16838
rect 15265 16836 15321 16838
rect 15345 16836 15401 16838
rect 14445 16346 14501 16348
rect 14525 16346 14581 16348
rect 14605 16346 14661 16348
rect 14685 16346 14741 16348
rect 14445 16294 14491 16346
rect 14491 16294 14501 16346
rect 14525 16294 14555 16346
rect 14555 16294 14567 16346
rect 14567 16294 14581 16346
rect 14605 16294 14619 16346
rect 14619 16294 14631 16346
rect 14631 16294 14661 16346
rect 14685 16294 14695 16346
rect 14695 16294 14741 16346
rect 14445 16292 14501 16294
rect 14525 16292 14581 16294
rect 14605 16292 14661 16294
rect 14685 16292 14741 16294
rect 13910 11736 13966 11792
rect 14445 15258 14501 15260
rect 14525 15258 14581 15260
rect 14605 15258 14661 15260
rect 14685 15258 14741 15260
rect 14445 15206 14491 15258
rect 14491 15206 14501 15258
rect 14525 15206 14555 15258
rect 14555 15206 14567 15258
rect 14567 15206 14581 15258
rect 14605 15206 14619 15258
rect 14619 15206 14631 15258
rect 14631 15206 14661 15258
rect 14685 15206 14695 15258
rect 14695 15206 14741 15258
rect 14445 15204 14501 15206
rect 14525 15204 14581 15206
rect 14605 15204 14661 15206
rect 14685 15204 14741 15206
rect 14445 14170 14501 14172
rect 14525 14170 14581 14172
rect 14605 14170 14661 14172
rect 14685 14170 14741 14172
rect 14445 14118 14491 14170
rect 14491 14118 14501 14170
rect 14525 14118 14555 14170
rect 14555 14118 14567 14170
rect 14567 14118 14581 14170
rect 14605 14118 14619 14170
rect 14619 14118 14631 14170
rect 14631 14118 14661 14170
rect 14685 14118 14695 14170
rect 14695 14118 14741 14170
rect 14445 14116 14501 14118
rect 14525 14116 14581 14118
rect 14605 14116 14661 14118
rect 14685 14116 14741 14118
rect 15105 15802 15161 15804
rect 15185 15802 15241 15804
rect 15265 15802 15321 15804
rect 15345 15802 15401 15804
rect 15105 15750 15151 15802
rect 15151 15750 15161 15802
rect 15185 15750 15215 15802
rect 15215 15750 15227 15802
rect 15227 15750 15241 15802
rect 15265 15750 15279 15802
rect 15279 15750 15291 15802
rect 15291 15750 15321 15802
rect 15345 15750 15355 15802
rect 15355 15750 15401 15802
rect 15105 15748 15161 15750
rect 15185 15748 15241 15750
rect 15265 15748 15321 15750
rect 15345 15748 15401 15750
rect 16486 29164 16542 29200
rect 16486 29144 16488 29164
rect 16488 29144 16540 29164
rect 16540 29144 16542 29164
rect 16670 24812 16726 24848
rect 16670 24792 16672 24812
rect 16672 24792 16724 24812
rect 16724 24792 16726 24812
rect 16486 23196 16488 23216
rect 16488 23196 16540 23216
rect 16540 23196 16542 23216
rect 16486 23160 16542 23196
rect 16026 17856 16082 17912
rect 15105 14714 15161 14716
rect 15185 14714 15241 14716
rect 15265 14714 15321 14716
rect 15345 14714 15401 14716
rect 15105 14662 15151 14714
rect 15151 14662 15161 14714
rect 15185 14662 15215 14714
rect 15215 14662 15227 14714
rect 15227 14662 15241 14714
rect 15265 14662 15279 14714
rect 15279 14662 15291 14714
rect 15291 14662 15321 14714
rect 15345 14662 15355 14714
rect 15355 14662 15401 14714
rect 15105 14660 15161 14662
rect 15185 14660 15241 14662
rect 15265 14660 15321 14662
rect 15345 14660 15401 14662
rect 14738 13776 14794 13832
rect 14445 13082 14501 13084
rect 14525 13082 14581 13084
rect 14605 13082 14661 13084
rect 14685 13082 14741 13084
rect 14445 13030 14491 13082
rect 14491 13030 14501 13082
rect 14525 13030 14555 13082
rect 14555 13030 14567 13082
rect 14567 13030 14581 13082
rect 14605 13030 14619 13082
rect 14619 13030 14631 13082
rect 14631 13030 14661 13082
rect 14685 13030 14695 13082
rect 14695 13030 14741 13082
rect 14445 13028 14501 13030
rect 14525 13028 14581 13030
rect 14605 13028 14661 13030
rect 14685 13028 14741 13030
rect 15474 14048 15530 14104
rect 15566 13776 15622 13832
rect 15566 13640 15622 13696
rect 15105 13626 15161 13628
rect 15185 13626 15241 13628
rect 15265 13626 15321 13628
rect 15345 13626 15401 13628
rect 15105 13574 15151 13626
rect 15151 13574 15161 13626
rect 15185 13574 15215 13626
rect 15215 13574 15227 13626
rect 15227 13574 15241 13626
rect 15265 13574 15279 13626
rect 15279 13574 15291 13626
rect 15291 13574 15321 13626
rect 15345 13574 15355 13626
rect 15355 13574 15401 13626
rect 15105 13572 15161 13574
rect 15185 13572 15241 13574
rect 15265 13572 15321 13574
rect 15345 13572 15401 13574
rect 15198 13232 15254 13288
rect 15474 12844 15530 12880
rect 15474 12824 15476 12844
rect 15476 12824 15528 12844
rect 15528 12824 15530 12844
rect 15105 12538 15161 12540
rect 15185 12538 15241 12540
rect 15265 12538 15321 12540
rect 15345 12538 15401 12540
rect 15105 12486 15151 12538
rect 15151 12486 15161 12538
rect 15185 12486 15215 12538
rect 15215 12486 15227 12538
rect 15227 12486 15241 12538
rect 15265 12486 15279 12538
rect 15279 12486 15291 12538
rect 15291 12486 15321 12538
rect 15345 12486 15355 12538
rect 15355 12486 15401 12538
rect 15105 12484 15161 12486
rect 15185 12484 15241 12486
rect 15265 12484 15321 12486
rect 15345 12484 15401 12486
rect 14445 11994 14501 11996
rect 14525 11994 14581 11996
rect 14605 11994 14661 11996
rect 14685 11994 14741 11996
rect 14445 11942 14491 11994
rect 14491 11942 14501 11994
rect 14525 11942 14555 11994
rect 14555 11942 14567 11994
rect 14567 11942 14581 11994
rect 14605 11942 14619 11994
rect 14619 11942 14631 11994
rect 14631 11942 14661 11994
rect 14685 11942 14695 11994
rect 14695 11942 14741 11994
rect 14445 11940 14501 11942
rect 14525 11940 14581 11942
rect 14605 11940 14661 11942
rect 14685 11940 14741 11942
rect 14738 11056 14794 11112
rect 14445 10906 14501 10908
rect 14525 10906 14581 10908
rect 14605 10906 14661 10908
rect 14685 10906 14741 10908
rect 14445 10854 14491 10906
rect 14491 10854 14501 10906
rect 14525 10854 14555 10906
rect 14555 10854 14567 10906
rect 14567 10854 14581 10906
rect 14605 10854 14619 10906
rect 14619 10854 14631 10906
rect 14631 10854 14661 10906
rect 14685 10854 14695 10906
rect 14695 10854 14741 10906
rect 14445 10852 14501 10854
rect 14525 10852 14581 10854
rect 14605 10852 14661 10854
rect 14685 10852 14741 10854
rect 15474 12180 15476 12200
rect 15476 12180 15528 12200
rect 15528 12180 15530 12200
rect 15474 12144 15530 12180
rect 15105 11450 15161 11452
rect 15185 11450 15241 11452
rect 15265 11450 15321 11452
rect 15345 11450 15401 11452
rect 15105 11398 15151 11450
rect 15151 11398 15161 11450
rect 15185 11398 15215 11450
rect 15215 11398 15227 11450
rect 15227 11398 15241 11450
rect 15265 11398 15279 11450
rect 15279 11398 15291 11450
rect 15291 11398 15321 11450
rect 15345 11398 15355 11450
rect 15355 11398 15401 11450
rect 15105 11396 15161 11398
rect 15185 11396 15241 11398
rect 15265 11396 15321 11398
rect 15345 11396 15401 11398
rect 15105 10362 15161 10364
rect 15185 10362 15241 10364
rect 15265 10362 15321 10364
rect 15345 10362 15401 10364
rect 15105 10310 15151 10362
rect 15151 10310 15161 10362
rect 15185 10310 15215 10362
rect 15215 10310 15227 10362
rect 15227 10310 15241 10362
rect 15265 10310 15279 10362
rect 15279 10310 15291 10362
rect 15291 10310 15321 10362
rect 15345 10310 15355 10362
rect 15355 10310 15401 10362
rect 15105 10308 15161 10310
rect 15185 10308 15241 10310
rect 15265 10308 15321 10310
rect 15345 10308 15401 10310
rect 14445 9818 14501 9820
rect 14525 9818 14581 9820
rect 14605 9818 14661 9820
rect 14685 9818 14741 9820
rect 14445 9766 14491 9818
rect 14491 9766 14501 9818
rect 14525 9766 14555 9818
rect 14555 9766 14567 9818
rect 14567 9766 14581 9818
rect 14605 9766 14619 9818
rect 14619 9766 14631 9818
rect 14631 9766 14661 9818
rect 14685 9766 14695 9818
rect 14695 9766 14741 9818
rect 14445 9764 14501 9766
rect 14525 9764 14581 9766
rect 14605 9764 14661 9766
rect 14685 9764 14741 9766
rect 15105 9274 15161 9276
rect 15185 9274 15241 9276
rect 15265 9274 15321 9276
rect 15345 9274 15401 9276
rect 15105 9222 15151 9274
rect 15151 9222 15161 9274
rect 15185 9222 15215 9274
rect 15215 9222 15227 9274
rect 15227 9222 15241 9274
rect 15265 9222 15279 9274
rect 15279 9222 15291 9274
rect 15291 9222 15321 9274
rect 15345 9222 15355 9274
rect 15355 9222 15401 9274
rect 15105 9220 15161 9222
rect 15185 9220 15241 9222
rect 15265 9220 15321 9222
rect 15345 9220 15401 9222
rect 14554 9016 14610 9072
rect 14445 8730 14501 8732
rect 14525 8730 14581 8732
rect 14605 8730 14661 8732
rect 14685 8730 14741 8732
rect 14445 8678 14491 8730
rect 14491 8678 14501 8730
rect 14525 8678 14555 8730
rect 14555 8678 14567 8730
rect 14567 8678 14581 8730
rect 14605 8678 14619 8730
rect 14619 8678 14631 8730
rect 14631 8678 14661 8730
rect 14685 8678 14695 8730
rect 14695 8678 14741 8730
rect 14445 8676 14501 8678
rect 14525 8676 14581 8678
rect 14605 8676 14661 8678
rect 14685 8676 14741 8678
rect 12162 5652 12164 5672
rect 12164 5652 12216 5672
rect 12216 5652 12218 5672
rect 12162 5616 12218 5652
rect 15105 8186 15161 8188
rect 15185 8186 15241 8188
rect 15265 8186 15321 8188
rect 15345 8186 15401 8188
rect 15105 8134 15151 8186
rect 15151 8134 15161 8186
rect 15185 8134 15215 8186
rect 15215 8134 15227 8186
rect 15227 8134 15241 8186
rect 15265 8134 15279 8186
rect 15279 8134 15291 8186
rect 15291 8134 15321 8186
rect 15345 8134 15355 8186
rect 15355 8134 15401 8186
rect 15105 8132 15161 8134
rect 15185 8132 15241 8134
rect 15265 8132 15321 8134
rect 15345 8132 15401 8134
rect 14445 7642 14501 7644
rect 14525 7642 14581 7644
rect 14605 7642 14661 7644
rect 14685 7642 14741 7644
rect 14445 7590 14491 7642
rect 14491 7590 14501 7642
rect 14525 7590 14555 7642
rect 14555 7590 14567 7642
rect 14567 7590 14581 7642
rect 14605 7590 14619 7642
rect 14619 7590 14631 7642
rect 14631 7590 14661 7642
rect 14685 7590 14695 7642
rect 14695 7590 14741 7642
rect 14445 7588 14501 7590
rect 14525 7588 14581 7590
rect 14605 7588 14661 7590
rect 14685 7588 14741 7590
rect 14445 6554 14501 6556
rect 14525 6554 14581 6556
rect 14605 6554 14661 6556
rect 14685 6554 14741 6556
rect 14445 6502 14491 6554
rect 14491 6502 14501 6554
rect 14525 6502 14555 6554
rect 14555 6502 14567 6554
rect 14567 6502 14581 6554
rect 14605 6502 14619 6554
rect 14619 6502 14631 6554
rect 14631 6502 14661 6554
rect 14685 6502 14695 6554
rect 14695 6502 14741 6554
rect 14445 6500 14501 6502
rect 14525 6500 14581 6502
rect 14605 6500 14661 6502
rect 14685 6500 14741 6502
rect 14445 5466 14501 5468
rect 14525 5466 14581 5468
rect 14605 5466 14661 5468
rect 14685 5466 14741 5468
rect 14445 5414 14491 5466
rect 14491 5414 14501 5466
rect 14525 5414 14555 5466
rect 14555 5414 14567 5466
rect 14567 5414 14581 5466
rect 14605 5414 14619 5466
rect 14619 5414 14631 5466
rect 14631 5414 14661 5466
rect 14685 5414 14695 5466
rect 14695 5414 14741 5466
rect 14445 5412 14501 5414
rect 14525 5412 14581 5414
rect 14605 5412 14661 5414
rect 14685 5412 14741 5414
rect 15105 7098 15161 7100
rect 15185 7098 15241 7100
rect 15265 7098 15321 7100
rect 15345 7098 15401 7100
rect 15105 7046 15151 7098
rect 15151 7046 15161 7098
rect 15185 7046 15215 7098
rect 15215 7046 15227 7098
rect 15227 7046 15241 7098
rect 15265 7046 15279 7098
rect 15279 7046 15291 7098
rect 15291 7046 15321 7098
rect 15345 7046 15355 7098
rect 15355 7046 15401 7098
rect 15105 7044 15161 7046
rect 15185 7044 15241 7046
rect 15265 7044 15321 7046
rect 15345 7044 15401 7046
rect 15934 11228 15936 11248
rect 15936 11228 15988 11248
rect 15988 11228 15990 11248
rect 15934 11192 15990 11228
rect 19062 33260 19064 33280
rect 19064 33260 19116 33280
rect 19116 33260 19118 33280
rect 19062 33224 19118 33260
rect 18786 32272 18842 32328
rect 22994 34298 23050 34300
rect 23074 34298 23130 34300
rect 23154 34298 23210 34300
rect 23234 34298 23290 34300
rect 22994 34246 23040 34298
rect 23040 34246 23050 34298
rect 23074 34246 23104 34298
rect 23104 34246 23116 34298
rect 23116 34246 23130 34298
rect 23154 34246 23168 34298
rect 23168 34246 23180 34298
rect 23180 34246 23210 34298
rect 23234 34246 23244 34298
rect 23244 34246 23290 34298
rect 22994 34244 23050 34246
rect 23074 34244 23130 34246
rect 23154 34244 23210 34246
rect 23234 34244 23290 34246
rect 21546 33260 21548 33280
rect 21548 33260 21600 33280
rect 21600 33260 21602 33280
rect 21546 33224 21602 33260
rect 17406 26308 17462 26344
rect 17406 26288 17408 26308
rect 17408 26288 17460 26308
rect 17460 26288 17462 26308
rect 17130 21548 17186 21584
rect 17130 21528 17132 21548
rect 17132 21528 17184 21548
rect 17184 21528 17186 21548
rect 17130 20440 17186 20496
rect 16302 13368 16358 13424
rect 18970 25764 19026 25800
rect 18970 25744 18972 25764
rect 18972 25744 19024 25764
rect 19024 25744 19026 25764
rect 16578 13132 16580 13152
rect 16580 13132 16632 13152
rect 16632 13132 16634 13152
rect 16578 13096 16634 13132
rect 16854 12980 16910 13016
rect 16854 12960 16856 12980
rect 16856 12960 16908 12980
rect 16908 12960 16910 12980
rect 17130 13096 17186 13152
rect 18142 17584 18198 17640
rect 19614 28056 19670 28112
rect 20074 27956 20076 27976
rect 20076 27956 20128 27976
rect 20128 27956 20130 27976
rect 20074 27920 20130 27956
rect 19062 20304 19118 20360
rect 18786 18300 18788 18320
rect 18788 18300 18840 18320
rect 18840 18300 18842 18320
rect 18786 18264 18842 18300
rect 18142 17040 18198 17096
rect 19706 20712 19762 20768
rect 19522 18808 19578 18864
rect 17682 14048 17738 14104
rect 17590 13640 17646 13696
rect 17314 13368 17370 13424
rect 17406 12688 17462 12744
rect 17406 11872 17462 11928
rect 17958 12960 18014 13016
rect 17590 11212 17646 11248
rect 17590 11192 17592 11212
rect 17592 11192 17644 11212
rect 17644 11192 17646 11212
rect 16946 10920 17002 10976
rect 17498 9424 17554 9480
rect 17866 9424 17922 9480
rect 18050 12280 18106 12336
rect 18050 11736 18106 11792
rect 18050 9016 18106 9072
rect 15105 6010 15161 6012
rect 15185 6010 15241 6012
rect 15265 6010 15321 6012
rect 15345 6010 15401 6012
rect 15105 5958 15151 6010
rect 15151 5958 15161 6010
rect 15185 5958 15215 6010
rect 15215 5958 15227 6010
rect 15227 5958 15241 6010
rect 15265 5958 15279 6010
rect 15279 5958 15291 6010
rect 15291 5958 15321 6010
rect 15345 5958 15355 6010
rect 15355 5958 15401 6010
rect 15105 5956 15161 5958
rect 15185 5956 15241 5958
rect 15265 5956 15321 5958
rect 15345 5956 15401 5958
rect 16670 5616 16726 5672
rect 14445 4378 14501 4380
rect 14525 4378 14581 4380
rect 14605 4378 14661 4380
rect 14685 4378 14741 4380
rect 14445 4326 14491 4378
rect 14491 4326 14501 4378
rect 14525 4326 14555 4378
rect 14555 4326 14567 4378
rect 14567 4326 14581 4378
rect 14605 4326 14619 4378
rect 14619 4326 14631 4378
rect 14631 4326 14661 4378
rect 14685 4326 14695 4378
rect 14695 4326 14741 4378
rect 14445 4324 14501 4326
rect 14525 4324 14581 4326
rect 14605 4324 14661 4326
rect 14685 4324 14741 4326
rect 15105 4922 15161 4924
rect 15185 4922 15241 4924
rect 15265 4922 15321 4924
rect 15345 4922 15401 4924
rect 15105 4870 15151 4922
rect 15151 4870 15161 4922
rect 15185 4870 15215 4922
rect 15215 4870 15227 4922
rect 15227 4870 15241 4922
rect 15265 4870 15279 4922
rect 15279 4870 15291 4922
rect 15291 4870 15321 4922
rect 15345 4870 15355 4922
rect 15355 4870 15401 4922
rect 15105 4868 15161 4870
rect 15185 4868 15241 4870
rect 15265 4868 15321 4870
rect 15345 4868 15401 4870
rect 15105 3834 15161 3836
rect 15185 3834 15241 3836
rect 15265 3834 15321 3836
rect 15345 3834 15401 3836
rect 15105 3782 15151 3834
rect 15151 3782 15161 3834
rect 15185 3782 15215 3834
rect 15215 3782 15227 3834
rect 15227 3782 15241 3834
rect 15265 3782 15279 3834
rect 15279 3782 15291 3834
rect 15291 3782 15321 3834
rect 15345 3782 15355 3834
rect 15355 3782 15401 3834
rect 15105 3780 15161 3782
rect 15185 3780 15241 3782
rect 15265 3780 15321 3782
rect 15345 3780 15401 3782
rect 14445 3290 14501 3292
rect 14525 3290 14581 3292
rect 14605 3290 14661 3292
rect 14685 3290 14741 3292
rect 14445 3238 14491 3290
rect 14491 3238 14501 3290
rect 14525 3238 14555 3290
rect 14555 3238 14567 3290
rect 14567 3238 14581 3290
rect 14605 3238 14619 3290
rect 14619 3238 14631 3290
rect 14631 3238 14661 3290
rect 14685 3238 14695 3290
rect 14695 3238 14741 3290
rect 14445 3236 14501 3238
rect 14525 3236 14581 3238
rect 14605 3236 14661 3238
rect 14685 3236 14741 3238
rect 15105 2746 15161 2748
rect 15185 2746 15241 2748
rect 15265 2746 15321 2748
rect 15345 2746 15401 2748
rect 15105 2694 15151 2746
rect 15151 2694 15161 2746
rect 15185 2694 15215 2746
rect 15215 2694 15227 2746
rect 15227 2694 15241 2746
rect 15265 2694 15279 2746
rect 15279 2694 15291 2746
rect 15291 2694 15321 2746
rect 15345 2694 15355 2746
rect 15355 2694 15401 2746
rect 15105 2692 15161 2694
rect 15185 2692 15241 2694
rect 15265 2692 15321 2694
rect 15345 2692 15401 2694
rect 18418 12280 18474 12336
rect 18786 13776 18842 13832
rect 18694 12688 18750 12744
rect 19522 17992 19578 18048
rect 19522 17740 19578 17776
rect 19522 17720 19524 17740
rect 19524 17720 19576 17740
rect 19576 17720 19578 17740
rect 19246 15272 19302 15328
rect 18970 13640 19026 13696
rect 18786 9036 18842 9072
rect 18786 9016 18788 9036
rect 18788 9016 18840 9036
rect 18840 9016 18842 9036
rect 18786 8200 18842 8256
rect 18602 8064 18658 8120
rect 19706 17856 19762 17912
rect 19246 11892 19302 11928
rect 19522 12300 19578 12336
rect 19522 12280 19524 12300
rect 19524 12280 19576 12300
rect 19576 12280 19578 12300
rect 19246 11872 19248 11892
rect 19248 11872 19300 11892
rect 19300 11872 19302 11892
rect 19338 11620 19394 11656
rect 19338 11600 19340 11620
rect 19340 11600 19392 11620
rect 19392 11600 19394 11620
rect 19614 9560 19670 9616
rect 19338 6296 19394 6352
rect 20074 19352 20130 19408
rect 20534 20304 20590 20360
rect 20350 18828 20406 18864
rect 20350 18808 20352 18828
rect 20352 18808 20404 18828
rect 20404 18808 20406 18828
rect 20534 17176 20590 17232
rect 20166 15952 20222 16008
rect 20074 15136 20130 15192
rect 20074 13676 20076 13696
rect 20076 13676 20128 13696
rect 20128 13676 20130 13696
rect 20074 13640 20130 13676
rect 22334 33754 22390 33756
rect 22414 33754 22470 33756
rect 22494 33754 22550 33756
rect 22574 33754 22630 33756
rect 22334 33702 22380 33754
rect 22380 33702 22390 33754
rect 22414 33702 22444 33754
rect 22444 33702 22456 33754
rect 22456 33702 22470 33754
rect 22494 33702 22508 33754
rect 22508 33702 22520 33754
rect 22520 33702 22550 33754
rect 22574 33702 22584 33754
rect 22584 33702 22630 33754
rect 22334 33700 22390 33702
rect 22414 33700 22470 33702
rect 22494 33700 22550 33702
rect 22574 33700 22630 33702
rect 22334 32666 22390 32668
rect 22414 32666 22470 32668
rect 22494 32666 22550 32668
rect 22574 32666 22630 32668
rect 22334 32614 22380 32666
rect 22380 32614 22390 32666
rect 22414 32614 22444 32666
rect 22444 32614 22456 32666
rect 22456 32614 22470 32666
rect 22494 32614 22508 32666
rect 22508 32614 22520 32666
rect 22520 32614 22550 32666
rect 22574 32614 22584 32666
rect 22584 32614 22630 32666
rect 22334 32612 22390 32614
rect 22414 32612 22470 32614
rect 22494 32612 22550 32614
rect 22574 32612 22630 32614
rect 22994 33210 23050 33212
rect 23074 33210 23130 33212
rect 23154 33210 23210 33212
rect 23234 33210 23290 33212
rect 22994 33158 23040 33210
rect 23040 33158 23050 33210
rect 23074 33158 23104 33210
rect 23104 33158 23116 33210
rect 23116 33158 23130 33210
rect 23154 33158 23168 33210
rect 23168 33158 23180 33210
rect 23180 33158 23210 33210
rect 23234 33158 23244 33210
rect 23244 33158 23290 33210
rect 22994 33156 23050 33158
rect 23074 33156 23130 33158
rect 23154 33156 23210 33158
rect 23234 33156 23290 33158
rect 22994 32122 23050 32124
rect 23074 32122 23130 32124
rect 23154 32122 23210 32124
rect 23234 32122 23290 32124
rect 22994 32070 23040 32122
rect 23040 32070 23050 32122
rect 23074 32070 23104 32122
rect 23104 32070 23116 32122
rect 23116 32070 23130 32122
rect 23154 32070 23168 32122
rect 23168 32070 23180 32122
rect 23180 32070 23210 32122
rect 23234 32070 23244 32122
rect 23244 32070 23290 32122
rect 22994 32068 23050 32070
rect 23074 32068 23130 32070
rect 23154 32068 23210 32070
rect 23234 32068 23290 32070
rect 22334 31578 22390 31580
rect 22414 31578 22470 31580
rect 22494 31578 22550 31580
rect 22574 31578 22630 31580
rect 22334 31526 22380 31578
rect 22380 31526 22390 31578
rect 22414 31526 22444 31578
rect 22444 31526 22456 31578
rect 22456 31526 22470 31578
rect 22494 31526 22508 31578
rect 22508 31526 22520 31578
rect 22520 31526 22550 31578
rect 22574 31526 22584 31578
rect 22584 31526 22630 31578
rect 22334 31524 22390 31526
rect 22414 31524 22470 31526
rect 22494 31524 22550 31526
rect 22574 31524 22630 31526
rect 22334 30490 22390 30492
rect 22414 30490 22470 30492
rect 22494 30490 22550 30492
rect 22574 30490 22630 30492
rect 22334 30438 22380 30490
rect 22380 30438 22390 30490
rect 22414 30438 22444 30490
rect 22444 30438 22456 30490
rect 22456 30438 22470 30490
rect 22494 30438 22508 30490
rect 22508 30438 22520 30490
rect 22520 30438 22550 30490
rect 22574 30438 22584 30490
rect 22584 30438 22630 30490
rect 22334 30436 22390 30438
rect 22414 30436 22470 30438
rect 22494 30436 22550 30438
rect 22574 30436 22630 30438
rect 22334 29402 22390 29404
rect 22414 29402 22470 29404
rect 22494 29402 22550 29404
rect 22574 29402 22630 29404
rect 22334 29350 22380 29402
rect 22380 29350 22390 29402
rect 22414 29350 22444 29402
rect 22444 29350 22456 29402
rect 22456 29350 22470 29402
rect 22494 29350 22508 29402
rect 22508 29350 22520 29402
rect 22520 29350 22550 29402
rect 22574 29350 22584 29402
rect 22584 29350 22630 29402
rect 22334 29348 22390 29350
rect 22414 29348 22470 29350
rect 22494 29348 22550 29350
rect 22574 29348 22630 29350
rect 22334 28314 22390 28316
rect 22414 28314 22470 28316
rect 22494 28314 22550 28316
rect 22574 28314 22630 28316
rect 22334 28262 22380 28314
rect 22380 28262 22390 28314
rect 22414 28262 22444 28314
rect 22444 28262 22456 28314
rect 22456 28262 22470 28314
rect 22494 28262 22508 28314
rect 22508 28262 22520 28314
rect 22520 28262 22550 28314
rect 22574 28262 22584 28314
rect 22584 28262 22630 28314
rect 22334 28260 22390 28262
rect 22414 28260 22470 28262
rect 22494 28260 22550 28262
rect 22574 28260 22630 28262
rect 22334 27226 22390 27228
rect 22414 27226 22470 27228
rect 22494 27226 22550 27228
rect 22574 27226 22630 27228
rect 22334 27174 22380 27226
rect 22380 27174 22390 27226
rect 22414 27174 22444 27226
rect 22444 27174 22456 27226
rect 22456 27174 22470 27226
rect 22494 27174 22508 27226
rect 22508 27174 22520 27226
rect 22520 27174 22550 27226
rect 22574 27174 22584 27226
rect 22584 27174 22630 27226
rect 22334 27172 22390 27174
rect 22414 27172 22470 27174
rect 22494 27172 22550 27174
rect 22574 27172 22630 27174
rect 22334 26138 22390 26140
rect 22414 26138 22470 26140
rect 22494 26138 22550 26140
rect 22574 26138 22630 26140
rect 22334 26086 22380 26138
rect 22380 26086 22390 26138
rect 22414 26086 22444 26138
rect 22444 26086 22456 26138
rect 22456 26086 22470 26138
rect 22494 26086 22508 26138
rect 22508 26086 22520 26138
rect 22520 26086 22550 26138
rect 22574 26086 22584 26138
rect 22584 26086 22630 26138
rect 22334 26084 22390 26086
rect 22414 26084 22470 26086
rect 22494 26084 22550 26086
rect 22574 26084 22630 26086
rect 22334 25050 22390 25052
rect 22414 25050 22470 25052
rect 22494 25050 22550 25052
rect 22574 25050 22630 25052
rect 22334 24998 22380 25050
rect 22380 24998 22390 25050
rect 22414 24998 22444 25050
rect 22444 24998 22456 25050
rect 22456 24998 22470 25050
rect 22494 24998 22508 25050
rect 22508 24998 22520 25050
rect 22520 24998 22550 25050
rect 22574 24998 22584 25050
rect 22584 24998 22630 25050
rect 22334 24996 22390 24998
rect 22414 24996 22470 24998
rect 22494 24996 22550 24998
rect 22574 24996 22630 24998
rect 22334 23962 22390 23964
rect 22414 23962 22470 23964
rect 22494 23962 22550 23964
rect 22574 23962 22630 23964
rect 22334 23910 22380 23962
rect 22380 23910 22390 23962
rect 22414 23910 22444 23962
rect 22444 23910 22456 23962
rect 22456 23910 22470 23962
rect 22494 23910 22508 23962
rect 22508 23910 22520 23962
rect 22520 23910 22550 23962
rect 22574 23910 22584 23962
rect 22584 23910 22630 23962
rect 22334 23908 22390 23910
rect 22414 23908 22470 23910
rect 22494 23908 22550 23910
rect 22574 23908 22630 23910
rect 22334 22874 22390 22876
rect 22414 22874 22470 22876
rect 22494 22874 22550 22876
rect 22574 22874 22630 22876
rect 22334 22822 22380 22874
rect 22380 22822 22390 22874
rect 22414 22822 22444 22874
rect 22444 22822 22456 22874
rect 22456 22822 22470 22874
rect 22494 22822 22508 22874
rect 22508 22822 22520 22874
rect 22520 22822 22550 22874
rect 22574 22822 22584 22874
rect 22584 22822 22630 22874
rect 22334 22820 22390 22822
rect 22414 22820 22470 22822
rect 22494 22820 22550 22822
rect 22574 22820 22630 22822
rect 22994 31034 23050 31036
rect 23074 31034 23130 31036
rect 23154 31034 23210 31036
rect 23234 31034 23290 31036
rect 22994 30982 23040 31034
rect 23040 30982 23050 31034
rect 23074 30982 23104 31034
rect 23104 30982 23116 31034
rect 23116 30982 23130 31034
rect 23154 30982 23168 31034
rect 23168 30982 23180 31034
rect 23180 30982 23210 31034
rect 23234 30982 23244 31034
rect 23244 30982 23290 31034
rect 22994 30980 23050 30982
rect 23074 30980 23130 30982
rect 23154 30980 23210 30982
rect 23234 30980 23290 30982
rect 22994 29946 23050 29948
rect 23074 29946 23130 29948
rect 23154 29946 23210 29948
rect 23234 29946 23290 29948
rect 22994 29894 23040 29946
rect 23040 29894 23050 29946
rect 23074 29894 23104 29946
rect 23104 29894 23116 29946
rect 23116 29894 23130 29946
rect 23154 29894 23168 29946
rect 23168 29894 23180 29946
rect 23180 29894 23210 29946
rect 23234 29894 23244 29946
rect 23244 29894 23290 29946
rect 22994 29892 23050 29894
rect 23074 29892 23130 29894
rect 23154 29892 23210 29894
rect 23234 29892 23290 29894
rect 22994 28858 23050 28860
rect 23074 28858 23130 28860
rect 23154 28858 23210 28860
rect 23234 28858 23290 28860
rect 22994 28806 23040 28858
rect 23040 28806 23050 28858
rect 23074 28806 23104 28858
rect 23104 28806 23116 28858
rect 23116 28806 23130 28858
rect 23154 28806 23168 28858
rect 23168 28806 23180 28858
rect 23180 28806 23210 28858
rect 23234 28806 23244 28858
rect 23244 28806 23290 28858
rect 22994 28804 23050 28806
rect 23074 28804 23130 28806
rect 23154 28804 23210 28806
rect 23234 28804 23290 28806
rect 22994 27770 23050 27772
rect 23074 27770 23130 27772
rect 23154 27770 23210 27772
rect 23234 27770 23290 27772
rect 22994 27718 23040 27770
rect 23040 27718 23050 27770
rect 23074 27718 23104 27770
rect 23104 27718 23116 27770
rect 23116 27718 23130 27770
rect 23154 27718 23168 27770
rect 23168 27718 23180 27770
rect 23180 27718 23210 27770
rect 23234 27718 23244 27770
rect 23244 27718 23290 27770
rect 22994 27716 23050 27718
rect 23074 27716 23130 27718
rect 23154 27716 23210 27718
rect 23234 27716 23290 27718
rect 22994 26682 23050 26684
rect 23074 26682 23130 26684
rect 23154 26682 23210 26684
rect 23234 26682 23290 26684
rect 22994 26630 23040 26682
rect 23040 26630 23050 26682
rect 23074 26630 23104 26682
rect 23104 26630 23116 26682
rect 23116 26630 23130 26682
rect 23154 26630 23168 26682
rect 23168 26630 23180 26682
rect 23180 26630 23210 26682
rect 23234 26630 23244 26682
rect 23244 26630 23290 26682
rect 22994 26628 23050 26630
rect 23074 26628 23130 26630
rect 23154 26628 23210 26630
rect 23234 26628 23290 26630
rect 30883 34298 30939 34300
rect 30963 34298 31019 34300
rect 31043 34298 31099 34300
rect 31123 34298 31179 34300
rect 30883 34246 30929 34298
rect 30929 34246 30939 34298
rect 30963 34246 30993 34298
rect 30993 34246 31005 34298
rect 31005 34246 31019 34298
rect 31043 34246 31057 34298
rect 31057 34246 31069 34298
rect 31069 34246 31099 34298
rect 31123 34246 31133 34298
rect 31133 34246 31179 34298
rect 30883 34244 30939 34246
rect 30963 34244 31019 34246
rect 31043 34244 31099 34246
rect 31123 34244 31179 34246
rect 22994 25594 23050 25596
rect 23074 25594 23130 25596
rect 23154 25594 23210 25596
rect 23234 25594 23290 25596
rect 22994 25542 23040 25594
rect 23040 25542 23050 25594
rect 23074 25542 23104 25594
rect 23104 25542 23116 25594
rect 23116 25542 23130 25594
rect 23154 25542 23168 25594
rect 23168 25542 23180 25594
rect 23180 25542 23210 25594
rect 23234 25542 23244 25594
rect 23244 25542 23290 25594
rect 22994 25540 23050 25542
rect 23074 25540 23130 25542
rect 23154 25540 23210 25542
rect 23234 25540 23290 25542
rect 22994 24506 23050 24508
rect 23074 24506 23130 24508
rect 23154 24506 23210 24508
rect 23234 24506 23290 24508
rect 22994 24454 23040 24506
rect 23040 24454 23050 24506
rect 23074 24454 23104 24506
rect 23104 24454 23116 24506
rect 23116 24454 23130 24506
rect 23154 24454 23168 24506
rect 23168 24454 23180 24506
rect 23180 24454 23210 24506
rect 23234 24454 23244 24506
rect 23244 24454 23290 24506
rect 22994 24452 23050 24454
rect 23074 24452 23130 24454
rect 23154 24452 23210 24454
rect 23234 24452 23290 24454
rect 22994 23418 23050 23420
rect 23074 23418 23130 23420
rect 23154 23418 23210 23420
rect 23234 23418 23290 23420
rect 22994 23366 23040 23418
rect 23040 23366 23050 23418
rect 23074 23366 23104 23418
rect 23104 23366 23116 23418
rect 23116 23366 23130 23418
rect 23154 23366 23168 23418
rect 23168 23366 23180 23418
rect 23180 23366 23210 23418
rect 23234 23366 23244 23418
rect 23244 23366 23290 23418
rect 22994 23364 23050 23366
rect 23074 23364 23130 23366
rect 23154 23364 23210 23366
rect 23234 23364 23290 23366
rect 22994 22330 23050 22332
rect 23074 22330 23130 22332
rect 23154 22330 23210 22332
rect 23234 22330 23290 22332
rect 22994 22278 23040 22330
rect 23040 22278 23050 22330
rect 23074 22278 23104 22330
rect 23104 22278 23116 22330
rect 23116 22278 23130 22330
rect 23154 22278 23168 22330
rect 23168 22278 23180 22330
rect 23180 22278 23210 22330
rect 23234 22278 23244 22330
rect 23244 22278 23290 22330
rect 22994 22276 23050 22278
rect 23074 22276 23130 22278
rect 23154 22276 23210 22278
rect 23234 22276 23290 22278
rect 21914 20340 21916 20360
rect 21916 20340 21968 20360
rect 21968 20340 21970 20360
rect 20902 15816 20958 15872
rect 21270 11736 21326 11792
rect 21914 20304 21970 20340
rect 22334 21786 22390 21788
rect 22414 21786 22470 21788
rect 22494 21786 22550 21788
rect 22574 21786 22630 21788
rect 22334 21734 22380 21786
rect 22380 21734 22390 21786
rect 22414 21734 22444 21786
rect 22444 21734 22456 21786
rect 22456 21734 22470 21786
rect 22494 21734 22508 21786
rect 22508 21734 22520 21786
rect 22520 21734 22550 21786
rect 22574 21734 22584 21786
rect 22584 21734 22630 21786
rect 22334 21732 22390 21734
rect 22414 21732 22470 21734
rect 22494 21732 22550 21734
rect 22574 21732 22630 21734
rect 22334 20698 22390 20700
rect 22414 20698 22470 20700
rect 22494 20698 22550 20700
rect 22574 20698 22630 20700
rect 22334 20646 22380 20698
rect 22380 20646 22390 20698
rect 22414 20646 22444 20698
rect 22444 20646 22456 20698
rect 22456 20646 22470 20698
rect 22494 20646 22508 20698
rect 22508 20646 22520 20698
rect 22520 20646 22550 20698
rect 22574 20646 22584 20698
rect 22584 20646 22630 20698
rect 22334 20644 22390 20646
rect 22414 20644 22470 20646
rect 22494 20644 22550 20646
rect 22574 20644 22630 20646
rect 22334 19610 22390 19612
rect 22414 19610 22470 19612
rect 22494 19610 22550 19612
rect 22574 19610 22630 19612
rect 22334 19558 22380 19610
rect 22380 19558 22390 19610
rect 22414 19558 22444 19610
rect 22444 19558 22456 19610
rect 22456 19558 22470 19610
rect 22494 19558 22508 19610
rect 22508 19558 22520 19610
rect 22520 19558 22550 19610
rect 22574 19558 22584 19610
rect 22584 19558 22630 19610
rect 22334 19556 22390 19558
rect 22414 19556 22470 19558
rect 22494 19556 22550 19558
rect 22574 19556 22630 19558
rect 21822 14728 21878 14784
rect 22334 18522 22390 18524
rect 22414 18522 22470 18524
rect 22494 18522 22550 18524
rect 22574 18522 22630 18524
rect 22334 18470 22380 18522
rect 22380 18470 22390 18522
rect 22414 18470 22444 18522
rect 22444 18470 22456 18522
rect 22456 18470 22470 18522
rect 22494 18470 22508 18522
rect 22508 18470 22520 18522
rect 22520 18470 22550 18522
rect 22574 18470 22584 18522
rect 22584 18470 22630 18522
rect 22334 18468 22390 18470
rect 22414 18468 22470 18470
rect 22494 18468 22550 18470
rect 22574 18468 22630 18470
rect 23202 22072 23258 22128
rect 22994 21242 23050 21244
rect 23074 21242 23130 21244
rect 23154 21242 23210 21244
rect 23234 21242 23290 21244
rect 22994 21190 23040 21242
rect 23040 21190 23050 21242
rect 23074 21190 23104 21242
rect 23104 21190 23116 21242
rect 23116 21190 23130 21242
rect 23154 21190 23168 21242
rect 23168 21190 23180 21242
rect 23180 21190 23210 21242
rect 23234 21190 23244 21242
rect 23244 21190 23290 21242
rect 22994 21188 23050 21190
rect 23074 21188 23130 21190
rect 23154 21188 23210 21190
rect 23234 21188 23290 21190
rect 22994 20154 23050 20156
rect 23074 20154 23130 20156
rect 23154 20154 23210 20156
rect 23234 20154 23290 20156
rect 22994 20102 23040 20154
rect 23040 20102 23050 20154
rect 23074 20102 23104 20154
rect 23104 20102 23116 20154
rect 23116 20102 23130 20154
rect 23154 20102 23168 20154
rect 23168 20102 23180 20154
rect 23180 20102 23210 20154
rect 23234 20102 23244 20154
rect 23244 20102 23290 20154
rect 22994 20100 23050 20102
rect 23074 20100 23130 20102
rect 23154 20100 23210 20102
rect 23234 20100 23290 20102
rect 22994 19066 23050 19068
rect 23074 19066 23130 19068
rect 23154 19066 23210 19068
rect 23234 19066 23290 19068
rect 22994 19014 23040 19066
rect 23040 19014 23050 19066
rect 23074 19014 23104 19066
rect 23104 19014 23116 19066
rect 23116 19014 23130 19066
rect 23154 19014 23168 19066
rect 23168 19014 23180 19066
rect 23180 19014 23210 19066
rect 23234 19014 23244 19066
rect 23244 19014 23290 19066
rect 22994 19012 23050 19014
rect 23074 19012 23130 19014
rect 23154 19012 23210 19014
rect 23234 19012 23290 19014
rect 23662 24112 23718 24168
rect 25042 28076 25098 28112
rect 25042 28056 25044 28076
rect 25044 28056 25096 28076
rect 25096 28056 25098 28076
rect 27710 29008 27766 29064
rect 26698 25744 26754 25800
rect 26606 24012 26608 24032
rect 26608 24012 26660 24032
rect 26660 24012 26662 24032
rect 26606 23976 26662 24012
rect 26054 22072 26110 22128
rect 22994 17978 23050 17980
rect 23074 17978 23130 17980
rect 23154 17978 23210 17980
rect 23234 17978 23290 17980
rect 22994 17926 23040 17978
rect 23040 17926 23050 17978
rect 23074 17926 23104 17978
rect 23104 17926 23116 17978
rect 23116 17926 23130 17978
rect 23154 17926 23168 17978
rect 23168 17926 23180 17978
rect 23180 17926 23210 17978
rect 23234 17926 23244 17978
rect 23244 17926 23290 17978
rect 22994 17924 23050 17926
rect 23074 17924 23130 17926
rect 23154 17924 23210 17926
rect 23234 17924 23290 17926
rect 22650 17720 22706 17776
rect 22334 17434 22390 17436
rect 22414 17434 22470 17436
rect 22494 17434 22550 17436
rect 22574 17434 22630 17436
rect 22334 17382 22380 17434
rect 22380 17382 22390 17434
rect 22414 17382 22444 17434
rect 22444 17382 22456 17434
rect 22456 17382 22470 17434
rect 22494 17382 22508 17434
rect 22508 17382 22520 17434
rect 22520 17382 22550 17434
rect 22574 17382 22584 17434
rect 22584 17382 22630 17434
rect 22334 17380 22390 17382
rect 22414 17380 22470 17382
rect 22494 17380 22550 17382
rect 22574 17380 22630 17382
rect 22334 16346 22390 16348
rect 22414 16346 22470 16348
rect 22494 16346 22550 16348
rect 22574 16346 22630 16348
rect 22334 16294 22380 16346
rect 22380 16294 22390 16346
rect 22414 16294 22444 16346
rect 22444 16294 22456 16346
rect 22456 16294 22470 16346
rect 22494 16294 22508 16346
rect 22508 16294 22520 16346
rect 22520 16294 22550 16346
rect 22574 16294 22584 16346
rect 22584 16294 22630 16346
rect 22334 16292 22390 16294
rect 22414 16292 22470 16294
rect 22494 16292 22550 16294
rect 22574 16292 22630 16294
rect 22334 15258 22390 15260
rect 22414 15258 22470 15260
rect 22494 15258 22550 15260
rect 22574 15258 22630 15260
rect 22334 15206 22380 15258
rect 22380 15206 22390 15258
rect 22414 15206 22444 15258
rect 22444 15206 22456 15258
rect 22456 15206 22470 15258
rect 22494 15206 22508 15258
rect 22508 15206 22520 15258
rect 22520 15206 22550 15258
rect 22574 15206 22584 15258
rect 22584 15206 22630 15258
rect 22334 15204 22390 15206
rect 22414 15204 22470 15206
rect 22494 15204 22550 15206
rect 22574 15204 22630 15206
rect 22190 14728 22246 14784
rect 22994 16890 23050 16892
rect 23074 16890 23130 16892
rect 23154 16890 23210 16892
rect 23234 16890 23290 16892
rect 22994 16838 23040 16890
rect 23040 16838 23050 16890
rect 23074 16838 23104 16890
rect 23104 16838 23116 16890
rect 23116 16838 23130 16890
rect 23154 16838 23168 16890
rect 23168 16838 23180 16890
rect 23180 16838 23210 16890
rect 23234 16838 23244 16890
rect 23244 16838 23290 16890
rect 22994 16836 23050 16838
rect 23074 16836 23130 16838
rect 23154 16836 23210 16838
rect 23234 16836 23290 16838
rect 22006 13676 22008 13696
rect 22008 13676 22060 13696
rect 22060 13676 22062 13696
rect 22006 13640 22062 13676
rect 22334 14170 22390 14172
rect 22414 14170 22470 14172
rect 22494 14170 22550 14172
rect 22574 14170 22630 14172
rect 22334 14118 22380 14170
rect 22380 14118 22390 14170
rect 22414 14118 22444 14170
rect 22444 14118 22456 14170
rect 22456 14118 22470 14170
rect 22494 14118 22508 14170
rect 22508 14118 22520 14170
rect 22520 14118 22550 14170
rect 22574 14118 22584 14170
rect 22584 14118 22630 14170
rect 22334 14116 22390 14118
rect 22414 14116 22470 14118
rect 22494 14116 22550 14118
rect 22574 14116 22630 14118
rect 22994 15802 23050 15804
rect 23074 15802 23130 15804
rect 23154 15802 23210 15804
rect 23234 15802 23290 15804
rect 22994 15750 23040 15802
rect 23040 15750 23050 15802
rect 23074 15750 23104 15802
rect 23104 15750 23116 15802
rect 23116 15750 23130 15802
rect 23154 15750 23168 15802
rect 23168 15750 23180 15802
rect 23180 15750 23210 15802
rect 23234 15750 23244 15802
rect 23244 15750 23290 15802
rect 22994 15748 23050 15750
rect 23074 15748 23130 15750
rect 23154 15748 23210 15750
rect 23234 15748 23290 15750
rect 22994 14714 23050 14716
rect 23074 14714 23130 14716
rect 23154 14714 23210 14716
rect 23234 14714 23290 14716
rect 22994 14662 23040 14714
rect 23040 14662 23050 14714
rect 23074 14662 23104 14714
rect 23104 14662 23116 14714
rect 23116 14662 23130 14714
rect 23154 14662 23168 14714
rect 23168 14662 23180 14714
rect 23180 14662 23210 14714
rect 23234 14662 23244 14714
rect 23244 14662 23290 14714
rect 22994 14660 23050 14662
rect 23074 14660 23130 14662
rect 23154 14660 23210 14662
rect 23234 14660 23290 14662
rect 23938 14456 23994 14512
rect 23386 13932 23442 13968
rect 23386 13912 23388 13932
rect 23388 13912 23440 13932
rect 23440 13912 23442 13932
rect 22994 13626 23050 13628
rect 23074 13626 23130 13628
rect 23154 13626 23210 13628
rect 23234 13626 23290 13628
rect 22994 13574 23040 13626
rect 23040 13574 23050 13626
rect 23074 13574 23104 13626
rect 23104 13574 23116 13626
rect 23116 13574 23130 13626
rect 23154 13574 23168 13626
rect 23168 13574 23180 13626
rect 23180 13574 23210 13626
rect 23234 13574 23244 13626
rect 23244 13574 23290 13626
rect 22994 13572 23050 13574
rect 23074 13572 23130 13574
rect 23154 13572 23210 13574
rect 23234 13572 23290 13574
rect 22334 13082 22390 13084
rect 22414 13082 22470 13084
rect 22494 13082 22550 13084
rect 22574 13082 22630 13084
rect 22334 13030 22380 13082
rect 22380 13030 22390 13082
rect 22414 13030 22444 13082
rect 22444 13030 22456 13082
rect 22456 13030 22470 13082
rect 22494 13030 22508 13082
rect 22508 13030 22520 13082
rect 22520 13030 22550 13082
rect 22574 13030 22584 13082
rect 22584 13030 22630 13082
rect 22334 13028 22390 13030
rect 22414 13028 22470 13030
rect 22494 13028 22550 13030
rect 22574 13028 22630 13030
rect 22334 11994 22390 11996
rect 22414 11994 22470 11996
rect 22494 11994 22550 11996
rect 22574 11994 22630 11996
rect 22334 11942 22380 11994
rect 22380 11942 22390 11994
rect 22414 11942 22444 11994
rect 22444 11942 22456 11994
rect 22456 11942 22470 11994
rect 22494 11942 22508 11994
rect 22508 11942 22520 11994
rect 22520 11942 22550 11994
rect 22574 11942 22584 11994
rect 22584 11942 22630 11994
rect 22334 11940 22390 11942
rect 22414 11940 22470 11942
rect 22494 11940 22550 11942
rect 22574 11940 22630 11942
rect 22994 12538 23050 12540
rect 23074 12538 23130 12540
rect 23154 12538 23210 12540
rect 23234 12538 23290 12540
rect 22994 12486 23040 12538
rect 23040 12486 23050 12538
rect 23074 12486 23104 12538
rect 23104 12486 23116 12538
rect 23116 12486 23130 12538
rect 23154 12486 23168 12538
rect 23168 12486 23180 12538
rect 23180 12486 23210 12538
rect 23234 12486 23244 12538
rect 23244 12486 23290 12538
rect 22994 12484 23050 12486
rect 23074 12484 23130 12486
rect 23154 12484 23210 12486
rect 23234 12484 23290 12486
rect 23570 12300 23626 12336
rect 23570 12280 23572 12300
rect 23572 12280 23624 12300
rect 23624 12280 23626 12300
rect 22006 11600 22062 11656
rect 22190 11600 22246 11656
rect 22334 10906 22390 10908
rect 22414 10906 22470 10908
rect 22494 10906 22550 10908
rect 22574 10906 22630 10908
rect 22334 10854 22380 10906
rect 22380 10854 22390 10906
rect 22414 10854 22444 10906
rect 22444 10854 22456 10906
rect 22456 10854 22470 10906
rect 22494 10854 22508 10906
rect 22508 10854 22520 10906
rect 22520 10854 22550 10906
rect 22574 10854 22584 10906
rect 22584 10854 22630 10906
rect 22334 10852 22390 10854
rect 22414 10852 22470 10854
rect 22494 10852 22550 10854
rect 22574 10852 22630 10854
rect 22994 11450 23050 11452
rect 23074 11450 23130 11452
rect 23154 11450 23210 11452
rect 23234 11450 23290 11452
rect 22994 11398 23040 11450
rect 23040 11398 23050 11450
rect 23074 11398 23104 11450
rect 23104 11398 23116 11450
rect 23116 11398 23130 11450
rect 23154 11398 23168 11450
rect 23168 11398 23180 11450
rect 23180 11398 23210 11450
rect 23234 11398 23244 11450
rect 23244 11398 23290 11450
rect 22994 11396 23050 11398
rect 23074 11396 23130 11398
rect 23154 11396 23210 11398
rect 23234 11396 23290 11398
rect 22334 9818 22390 9820
rect 22414 9818 22470 9820
rect 22494 9818 22550 9820
rect 22574 9818 22630 9820
rect 22334 9766 22380 9818
rect 22380 9766 22390 9818
rect 22414 9766 22444 9818
rect 22444 9766 22456 9818
rect 22456 9766 22470 9818
rect 22494 9766 22508 9818
rect 22508 9766 22520 9818
rect 22520 9766 22550 9818
rect 22574 9766 22584 9818
rect 22584 9766 22630 9818
rect 22334 9764 22390 9766
rect 22414 9764 22470 9766
rect 22494 9764 22550 9766
rect 22574 9764 22630 9766
rect 22098 8880 22154 8936
rect 22334 8730 22390 8732
rect 22414 8730 22470 8732
rect 22494 8730 22550 8732
rect 22574 8730 22630 8732
rect 22334 8678 22380 8730
rect 22380 8678 22390 8730
rect 22414 8678 22444 8730
rect 22444 8678 22456 8730
rect 22456 8678 22470 8730
rect 22494 8678 22508 8730
rect 22508 8678 22520 8730
rect 22520 8678 22550 8730
rect 22574 8678 22584 8730
rect 22584 8678 22630 8730
rect 22334 8676 22390 8678
rect 22414 8676 22470 8678
rect 22494 8676 22550 8678
rect 22574 8676 22630 8678
rect 22994 10362 23050 10364
rect 23074 10362 23130 10364
rect 23154 10362 23210 10364
rect 23234 10362 23290 10364
rect 22994 10310 23040 10362
rect 23040 10310 23050 10362
rect 23074 10310 23104 10362
rect 23104 10310 23116 10362
rect 23116 10310 23130 10362
rect 23154 10310 23168 10362
rect 23168 10310 23180 10362
rect 23180 10310 23210 10362
rect 23234 10310 23244 10362
rect 23244 10310 23290 10362
rect 22994 10308 23050 10310
rect 23074 10308 23130 10310
rect 23154 10308 23210 10310
rect 23234 10308 23290 10310
rect 22994 9274 23050 9276
rect 23074 9274 23130 9276
rect 23154 9274 23210 9276
rect 23234 9274 23290 9276
rect 22994 9222 23040 9274
rect 23040 9222 23050 9274
rect 23074 9222 23104 9274
rect 23104 9222 23116 9274
rect 23116 9222 23130 9274
rect 23154 9222 23168 9274
rect 23168 9222 23180 9274
rect 23180 9222 23210 9274
rect 23234 9222 23244 9274
rect 23244 9222 23290 9274
rect 22994 9220 23050 9222
rect 23074 9220 23130 9222
rect 23154 9220 23210 9222
rect 23234 9220 23290 9222
rect 21914 8472 21970 8528
rect 23110 8492 23166 8528
rect 23110 8472 23112 8492
rect 23112 8472 23164 8492
rect 23164 8472 23166 8492
rect 23386 8336 23442 8392
rect 22994 8186 23050 8188
rect 23074 8186 23130 8188
rect 23154 8186 23210 8188
rect 23234 8186 23290 8188
rect 22994 8134 23040 8186
rect 23040 8134 23050 8186
rect 23074 8134 23104 8186
rect 23104 8134 23116 8186
rect 23116 8134 23130 8186
rect 23154 8134 23168 8186
rect 23168 8134 23180 8186
rect 23180 8134 23210 8186
rect 23234 8134 23244 8186
rect 23244 8134 23290 8186
rect 22994 8132 23050 8134
rect 23074 8132 23130 8134
rect 23154 8132 23210 8134
rect 23234 8132 23290 8134
rect 22334 7642 22390 7644
rect 22414 7642 22470 7644
rect 22494 7642 22550 7644
rect 22574 7642 22630 7644
rect 22334 7590 22380 7642
rect 22380 7590 22390 7642
rect 22414 7590 22444 7642
rect 22444 7590 22456 7642
rect 22456 7590 22470 7642
rect 22494 7590 22508 7642
rect 22508 7590 22520 7642
rect 22520 7590 22550 7642
rect 22574 7590 22584 7642
rect 22584 7590 22630 7642
rect 22334 7588 22390 7590
rect 22414 7588 22470 7590
rect 22494 7588 22550 7590
rect 22574 7588 22630 7590
rect 22334 6554 22390 6556
rect 22414 6554 22470 6556
rect 22494 6554 22550 6556
rect 22574 6554 22630 6556
rect 22334 6502 22380 6554
rect 22380 6502 22390 6554
rect 22414 6502 22444 6554
rect 22444 6502 22456 6554
rect 22456 6502 22470 6554
rect 22494 6502 22508 6554
rect 22508 6502 22520 6554
rect 22520 6502 22550 6554
rect 22574 6502 22584 6554
rect 22584 6502 22630 6554
rect 22334 6500 22390 6502
rect 22414 6500 22470 6502
rect 22494 6500 22550 6502
rect 22574 6500 22630 6502
rect 22994 7098 23050 7100
rect 23074 7098 23130 7100
rect 23154 7098 23210 7100
rect 23234 7098 23290 7100
rect 22994 7046 23040 7098
rect 23040 7046 23050 7098
rect 23074 7046 23104 7098
rect 23104 7046 23116 7098
rect 23116 7046 23130 7098
rect 23154 7046 23168 7098
rect 23168 7046 23180 7098
rect 23180 7046 23210 7098
rect 23234 7046 23244 7098
rect 23244 7046 23290 7098
rect 22994 7044 23050 7046
rect 23074 7044 23130 7046
rect 23154 7044 23210 7046
rect 23234 7044 23290 7046
rect 22334 5466 22390 5468
rect 22414 5466 22470 5468
rect 22494 5466 22550 5468
rect 22574 5466 22630 5468
rect 22334 5414 22380 5466
rect 22380 5414 22390 5466
rect 22414 5414 22444 5466
rect 22444 5414 22456 5466
rect 22456 5414 22470 5466
rect 22494 5414 22508 5466
rect 22508 5414 22520 5466
rect 22520 5414 22550 5466
rect 22574 5414 22584 5466
rect 22584 5414 22630 5466
rect 22334 5412 22390 5414
rect 22414 5412 22470 5414
rect 22494 5412 22550 5414
rect 22574 5412 22630 5414
rect 24122 6860 24178 6896
rect 24122 6840 24124 6860
rect 24124 6840 24176 6860
rect 24176 6840 24178 6860
rect 22994 6010 23050 6012
rect 23074 6010 23130 6012
rect 23154 6010 23210 6012
rect 23234 6010 23290 6012
rect 22994 5958 23040 6010
rect 23040 5958 23050 6010
rect 23074 5958 23104 6010
rect 23104 5958 23116 6010
rect 23116 5958 23130 6010
rect 23154 5958 23168 6010
rect 23168 5958 23180 6010
rect 23180 5958 23210 6010
rect 23234 5958 23244 6010
rect 23244 5958 23290 6010
rect 22994 5956 23050 5958
rect 23074 5956 23130 5958
rect 23154 5956 23210 5958
rect 23234 5956 23290 5958
rect 22994 4922 23050 4924
rect 23074 4922 23130 4924
rect 23154 4922 23210 4924
rect 23234 4922 23290 4924
rect 22994 4870 23040 4922
rect 23040 4870 23050 4922
rect 23074 4870 23104 4922
rect 23104 4870 23116 4922
rect 23116 4870 23130 4922
rect 23154 4870 23168 4922
rect 23168 4870 23180 4922
rect 23180 4870 23210 4922
rect 23234 4870 23244 4922
rect 23244 4870 23290 4922
rect 22994 4868 23050 4870
rect 23074 4868 23130 4870
rect 23154 4868 23210 4870
rect 23234 4868 23290 4870
rect 22334 4378 22390 4380
rect 22414 4378 22470 4380
rect 22494 4378 22550 4380
rect 22574 4378 22630 4380
rect 22334 4326 22380 4378
rect 22380 4326 22390 4378
rect 22414 4326 22444 4378
rect 22444 4326 22456 4378
rect 22456 4326 22470 4378
rect 22494 4326 22508 4378
rect 22508 4326 22520 4378
rect 22520 4326 22550 4378
rect 22574 4326 22584 4378
rect 22584 4326 22630 4378
rect 22334 4324 22390 4326
rect 22414 4324 22470 4326
rect 22494 4324 22550 4326
rect 22574 4324 22630 4326
rect 22994 3834 23050 3836
rect 23074 3834 23130 3836
rect 23154 3834 23210 3836
rect 23234 3834 23290 3836
rect 22994 3782 23040 3834
rect 23040 3782 23050 3834
rect 23074 3782 23104 3834
rect 23104 3782 23116 3834
rect 23116 3782 23130 3834
rect 23154 3782 23168 3834
rect 23168 3782 23180 3834
rect 23180 3782 23210 3834
rect 23234 3782 23244 3834
rect 23244 3782 23290 3834
rect 22994 3780 23050 3782
rect 23074 3780 23130 3782
rect 23154 3780 23210 3782
rect 23234 3780 23290 3782
rect 22334 3290 22390 3292
rect 22414 3290 22470 3292
rect 22494 3290 22550 3292
rect 22574 3290 22630 3292
rect 22334 3238 22380 3290
rect 22380 3238 22390 3290
rect 22414 3238 22444 3290
rect 22444 3238 22456 3290
rect 22456 3238 22470 3290
rect 22494 3238 22508 3290
rect 22508 3238 22520 3290
rect 22520 3238 22550 3290
rect 22574 3238 22584 3290
rect 22584 3238 22630 3290
rect 22334 3236 22390 3238
rect 22414 3236 22470 3238
rect 22494 3236 22550 3238
rect 22574 3236 22630 3238
rect 27986 27512 28042 27568
rect 28906 27920 28962 27976
rect 27618 22108 27620 22128
rect 27620 22108 27672 22128
rect 27672 22108 27674 22128
rect 27618 22072 27674 22108
rect 30223 33754 30279 33756
rect 30303 33754 30359 33756
rect 30383 33754 30439 33756
rect 30463 33754 30519 33756
rect 30223 33702 30269 33754
rect 30269 33702 30279 33754
rect 30303 33702 30333 33754
rect 30333 33702 30345 33754
rect 30345 33702 30359 33754
rect 30383 33702 30397 33754
rect 30397 33702 30409 33754
rect 30409 33702 30439 33754
rect 30463 33702 30473 33754
rect 30473 33702 30519 33754
rect 30223 33700 30279 33702
rect 30303 33700 30359 33702
rect 30383 33700 30439 33702
rect 30463 33700 30519 33702
rect 30883 33210 30939 33212
rect 30963 33210 31019 33212
rect 31043 33210 31099 33212
rect 31123 33210 31179 33212
rect 30883 33158 30929 33210
rect 30929 33158 30939 33210
rect 30963 33158 30993 33210
rect 30993 33158 31005 33210
rect 31005 33158 31019 33210
rect 31043 33158 31057 33210
rect 31057 33158 31069 33210
rect 31069 33158 31099 33210
rect 31123 33158 31133 33210
rect 31133 33158 31179 33210
rect 30883 33156 30939 33158
rect 30963 33156 31019 33158
rect 31043 33156 31099 33158
rect 31123 33156 31179 33158
rect 30223 32666 30279 32668
rect 30303 32666 30359 32668
rect 30383 32666 30439 32668
rect 30463 32666 30519 32668
rect 30223 32614 30269 32666
rect 30269 32614 30279 32666
rect 30303 32614 30333 32666
rect 30333 32614 30345 32666
rect 30345 32614 30359 32666
rect 30383 32614 30397 32666
rect 30397 32614 30409 32666
rect 30409 32614 30439 32666
rect 30463 32614 30473 32666
rect 30473 32614 30519 32666
rect 30223 32612 30279 32614
rect 30303 32612 30359 32614
rect 30383 32612 30439 32614
rect 30463 32612 30519 32614
rect 30883 32122 30939 32124
rect 30963 32122 31019 32124
rect 31043 32122 31099 32124
rect 31123 32122 31179 32124
rect 30883 32070 30929 32122
rect 30929 32070 30939 32122
rect 30963 32070 30993 32122
rect 30993 32070 31005 32122
rect 31005 32070 31019 32122
rect 31043 32070 31057 32122
rect 31057 32070 31069 32122
rect 31069 32070 31099 32122
rect 31123 32070 31133 32122
rect 31133 32070 31179 32122
rect 30883 32068 30939 32070
rect 30963 32068 31019 32070
rect 31043 32068 31099 32070
rect 31123 32068 31179 32070
rect 30223 31578 30279 31580
rect 30303 31578 30359 31580
rect 30383 31578 30439 31580
rect 30463 31578 30519 31580
rect 30223 31526 30269 31578
rect 30269 31526 30279 31578
rect 30303 31526 30333 31578
rect 30333 31526 30345 31578
rect 30345 31526 30359 31578
rect 30383 31526 30397 31578
rect 30397 31526 30409 31578
rect 30409 31526 30439 31578
rect 30463 31526 30473 31578
rect 30473 31526 30519 31578
rect 30223 31524 30279 31526
rect 30303 31524 30359 31526
rect 30383 31524 30439 31526
rect 30463 31524 30519 31526
rect 30223 30490 30279 30492
rect 30303 30490 30359 30492
rect 30383 30490 30439 30492
rect 30463 30490 30519 30492
rect 30223 30438 30269 30490
rect 30269 30438 30279 30490
rect 30303 30438 30333 30490
rect 30333 30438 30345 30490
rect 30345 30438 30359 30490
rect 30383 30438 30397 30490
rect 30397 30438 30409 30490
rect 30409 30438 30439 30490
rect 30463 30438 30473 30490
rect 30473 30438 30519 30490
rect 30223 30436 30279 30438
rect 30303 30436 30359 30438
rect 30383 30436 30439 30438
rect 30463 30436 30519 30438
rect 30883 31034 30939 31036
rect 30963 31034 31019 31036
rect 31043 31034 31099 31036
rect 31123 31034 31179 31036
rect 30883 30982 30929 31034
rect 30929 30982 30939 31034
rect 30963 30982 30993 31034
rect 30993 30982 31005 31034
rect 31005 30982 31019 31034
rect 31043 30982 31057 31034
rect 31057 30982 31069 31034
rect 31069 30982 31099 31034
rect 31123 30982 31133 31034
rect 31133 30982 31179 31034
rect 30883 30980 30939 30982
rect 30963 30980 31019 30982
rect 31043 30980 31099 30982
rect 31123 30980 31179 30982
rect 33046 34040 33102 34096
rect 32126 31320 32182 31376
rect 30883 29946 30939 29948
rect 30963 29946 31019 29948
rect 31043 29946 31099 29948
rect 31123 29946 31179 29948
rect 30883 29894 30929 29946
rect 30929 29894 30939 29946
rect 30963 29894 30993 29946
rect 30993 29894 31005 29946
rect 31005 29894 31019 29946
rect 31043 29894 31057 29946
rect 31057 29894 31069 29946
rect 31069 29894 31099 29946
rect 31123 29894 31133 29946
rect 31133 29894 31179 29946
rect 30883 29892 30939 29894
rect 30963 29892 31019 29894
rect 31043 29892 31099 29894
rect 31123 29892 31179 29894
rect 30223 29402 30279 29404
rect 30303 29402 30359 29404
rect 30383 29402 30439 29404
rect 30463 29402 30519 29404
rect 30223 29350 30269 29402
rect 30269 29350 30279 29402
rect 30303 29350 30333 29402
rect 30333 29350 30345 29402
rect 30345 29350 30359 29402
rect 30383 29350 30397 29402
rect 30397 29350 30409 29402
rect 30409 29350 30439 29402
rect 30463 29350 30473 29402
rect 30473 29350 30519 29402
rect 30223 29348 30279 29350
rect 30303 29348 30359 29350
rect 30383 29348 30439 29350
rect 30463 29348 30519 29350
rect 30223 28314 30279 28316
rect 30303 28314 30359 28316
rect 30383 28314 30439 28316
rect 30463 28314 30519 28316
rect 30223 28262 30269 28314
rect 30269 28262 30279 28314
rect 30303 28262 30333 28314
rect 30333 28262 30345 28314
rect 30345 28262 30359 28314
rect 30383 28262 30397 28314
rect 30397 28262 30409 28314
rect 30409 28262 30439 28314
rect 30463 28262 30473 28314
rect 30473 28262 30519 28314
rect 30223 28260 30279 28262
rect 30303 28260 30359 28262
rect 30383 28260 30439 28262
rect 30463 28260 30519 28262
rect 30883 28858 30939 28860
rect 30963 28858 31019 28860
rect 31043 28858 31099 28860
rect 31123 28858 31179 28860
rect 30883 28806 30929 28858
rect 30929 28806 30939 28858
rect 30963 28806 30993 28858
rect 30993 28806 31005 28858
rect 31005 28806 31019 28858
rect 31043 28806 31057 28858
rect 31057 28806 31069 28858
rect 31069 28806 31099 28858
rect 31123 28806 31133 28858
rect 31133 28806 31179 28858
rect 30883 28804 30939 28806
rect 30963 28804 31019 28806
rect 31043 28804 31099 28806
rect 31123 28804 31179 28806
rect 30223 27226 30279 27228
rect 30303 27226 30359 27228
rect 30383 27226 30439 27228
rect 30463 27226 30519 27228
rect 30223 27174 30269 27226
rect 30269 27174 30279 27226
rect 30303 27174 30333 27226
rect 30333 27174 30345 27226
rect 30345 27174 30359 27226
rect 30383 27174 30397 27226
rect 30397 27174 30409 27226
rect 30409 27174 30439 27226
rect 30463 27174 30473 27226
rect 30473 27174 30519 27226
rect 30223 27172 30279 27174
rect 30303 27172 30359 27174
rect 30383 27172 30439 27174
rect 30463 27172 30519 27174
rect 30883 27770 30939 27772
rect 30963 27770 31019 27772
rect 31043 27770 31099 27772
rect 31123 27770 31179 27772
rect 30883 27718 30929 27770
rect 30929 27718 30939 27770
rect 30963 27718 30993 27770
rect 30993 27718 31005 27770
rect 31005 27718 31019 27770
rect 31043 27718 31057 27770
rect 31057 27718 31069 27770
rect 31069 27718 31099 27770
rect 31123 27718 31133 27770
rect 31133 27718 31179 27770
rect 30883 27716 30939 27718
rect 30963 27716 31019 27718
rect 31043 27716 31099 27718
rect 31123 27716 31179 27718
rect 30223 26138 30279 26140
rect 30303 26138 30359 26140
rect 30383 26138 30439 26140
rect 30463 26138 30519 26140
rect 30223 26086 30269 26138
rect 30269 26086 30279 26138
rect 30303 26086 30333 26138
rect 30333 26086 30345 26138
rect 30345 26086 30359 26138
rect 30383 26086 30397 26138
rect 30397 26086 30409 26138
rect 30409 26086 30439 26138
rect 30463 26086 30473 26138
rect 30473 26086 30519 26138
rect 30223 26084 30279 26086
rect 30303 26084 30359 26086
rect 30383 26084 30439 26086
rect 30463 26084 30519 26086
rect 30883 26682 30939 26684
rect 30963 26682 31019 26684
rect 31043 26682 31099 26684
rect 31123 26682 31179 26684
rect 30883 26630 30929 26682
rect 30929 26630 30939 26682
rect 30963 26630 30993 26682
rect 30993 26630 31005 26682
rect 31005 26630 31019 26682
rect 31043 26630 31057 26682
rect 31057 26630 31069 26682
rect 31069 26630 31099 26682
rect 31123 26630 31133 26682
rect 31133 26630 31179 26682
rect 30883 26628 30939 26630
rect 30963 26628 31019 26630
rect 31043 26628 31099 26630
rect 31123 26628 31179 26630
rect 33782 35400 33838 35456
rect 34886 32680 34942 32736
rect 33782 28600 33838 28656
rect 33046 27512 33102 27568
rect 30883 25594 30939 25596
rect 30963 25594 31019 25596
rect 31043 25594 31099 25596
rect 31123 25594 31179 25596
rect 30883 25542 30929 25594
rect 30929 25542 30939 25594
rect 30963 25542 30993 25594
rect 30993 25542 31005 25594
rect 31005 25542 31019 25594
rect 31043 25542 31057 25594
rect 31057 25542 31069 25594
rect 31069 25542 31099 25594
rect 31123 25542 31133 25594
rect 31133 25542 31179 25594
rect 30883 25540 30939 25542
rect 30963 25540 31019 25542
rect 31043 25540 31099 25542
rect 31123 25540 31179 25542
rect 28722 24112 28778 24168
rect 27986 22072 28042 22128
rect 26974 17212 26976 17232
rect 26976 17212 27028 17232
rect 27028 17212 27030 17232
rect 26974 17176 27030 17212
rect 26238 13640 26294 13696
rect 27986 19352 28042 19408
rect 28078 17856 28134 17912
rect 28262 17740 28318 17776
rect 28262 17720 28264 17740
rect 28264 17720 28316 17740
rect 28316 17720 28318 17740
rect 29182 19292 29238 19348
rect 29182 19080 29238 19136
rect 29366 18944 29422 19000
rect 30223 25050 30279 25052
rect 30303 25050 30359 25052
rect 30383 25050 30439 25052
rect 30463 25050 30519 25052
rect 30223 24998 30269 25050
rect 30269 24998 30279 25050
rect 30303 24998 30333 25050
rect 30333 24998 30345 25050
rect 30345 24998 30359 25050
rect 30383 24998 30397 25050
rect 30397 24998 30409 25050
rect 30409 24998 30439 25050
rect 30463 24998 30473 25050
rect 30473 24998 30519 25050
rect 30223 24996 30279 24998
rect 30303 24996 30359 24998
rect 30383 24996 30439 24998
rect 30463 24996 30519 24998
rect 30883 24506 30939 24508
rect 30963 24506 31019 24508
rect 31043 24506 31099 24508
rect 31123 24506 31179 24508
rect 30883 24454 30929 24506
rect 30929 24454 30939 24506
rect 30963 24454 30993 24506
rect 30993 24454 31005 24506
rect 31005 24454 31019 24506
rect 31043 24454 31057 24506
rect 31057 24454 31069 24506
rect 31069 24454 31099 24506
rect 31123 24454 31133 24506
rect 31133 24454 31179 24506
rect 30883 24452 30939 24454
rect 30963 24452 31019 24454
rect 31043 24452 31099 24454
rect 31123 24452 31179 24454
rect 30223 23962 30279 23964
rect 30303 23962 30359 23964
rect 30383 23962 30439 23964
rect 30463 23962 30519 23964
rect 30223 23910 30269 23962
rect 30269 23910 30279 23962
rect 30303 23910 30333 23962
rect 30333 23910 30345 23962
rect 30345 23910 30359 23962
rect 30383 23910 30397 23962
rect 30397 23910 30409 23962
rect 30409 23910 30439 23962
rect 30463 23910 30473 23962
rect 30473 23910 30519 23962
rect 30223 23908 30279 23910
rect 30303 23908 30359 23910
rect 30383 23908 30439 23910
rect 30463 23908 30519 23910
rect 30223 22874 30279 22876
rect 30303 22874 30359 22876
rect 30383 22874 30439 22876
rect 30463 22874 30519 22876
rect 30223 22822 30269 22874
rect 30269 22822 30279 22874
rect 30303 22822 30333 22874
rect 30333 22822 30345 22874
rect 30345 22822 30359 22874
rect 30383 22822 30397 22874
rect 30397 22822 30409 22874
rect 30409 22822 30439 22874
rect 30463 22822 30473 22874
rect 30473 22822 30519 22874
rect 30223 22820 30279 22822
rect 30303 22820 30359 22822
rect 30383 22820 30439 22822
rect 30463 22820 30519 22822
rect 30883 23418 30939 23420
rect 30963 23418 31019 23420
rect 31043 23418 31099 23420
rect 31123 23418 31179 23420
rect 30883 23366 30929 23418
rect 30929 23366 30939 23418
rect 30963 23366 30993 23418
rect 30993 23366 31005 23418
rect 31005 23366 31019 23418
rect 31043 23366 31057 23418
rect 31057 23366 31069 23418
rect 31069 23366 31099 23418
rect 31123 23366 31133 23418
rect 31133 23366 31179 23418
rect 30883 23364 30939 23366
rect 30963 23364 31019 23366
rect 31043 23364 31099 23366
rect 31123 23364 31179 23366
rect 30223 21786 30279 21788
rect 30303 21786 30359 21788
rect 30383 21786 30439 21788
rect 30463 21786 30519 21788
rect 30223 21734 30269 21786
rect 30269 21734 30279 21786
rect 30303 21734 30333 21786
rect 30333 21734 30345 21786
rect 30345 21734 30359 21786
rect 30383 21734 30397 21786
rect 30397 21734 30409 21786
rect 30409 21734 30439 21786
rect 30463 21734 30473 21786
rect 30473 21734 30519 21786
rect 30223 21732 30279 21734
rect 30303 21732 30359 21734
rect 30383 21732 30439 21734
rect 30463 21732 30519 21734
rect 30883 22330 30939 22332
rect 30963 22330 31019 22332
rect 31043 22330 31099 22332
rect 31123 22330 31179 22332
rect 30883 22278 30929 22330
rect 30929 22278 30939 22330
rect 30963 22278 30993 22330
rect 30993 22278 31005 22330
rect 31005 22278 31019 22330
rect 31043 22278 31057 22330
rect 31057 22278 31069 22330
rect 31069 22278 31099 22330
rect 31123 22278 31133 22330
rect 31133 22278 31179 22330
rect 30883 22276 30939 22278
rect 30963 22276 31019 22278
rect 31043 22276 31099 22278
rect 31123 22276 31179 22278
rect 30883 21242 30939 21244
rect 30963 21242 31019 21244
rect 31043 21242 31099 21244
rect 31123 21242 31179 21244
rect 30883 21190 30929 21242
rect 30929 21190 30939 21242
rect 30963 21190 30993 21242
rect 30993 21190 31005 21242
rect 31005 21190 31019 21242
rect 31043 21190 31057 21242
rect 31057 21190 31069 21242
rect 31069 21190 31099 21242
rect 31123 21190 31133 21242
rect 31133 21190 31179 21242
rect 30883 21188 30939 21190
rect 30963 21188 31019 21190
rect 31043 21188 31099 21190
rect 31123 21188 31179 21190
rect 30223 20698 30279 20700
rect 30303 20698 30359 20700
rect 30383 20698 30439 20700
rect 30463 20698 30519 20700
rect 30223 20646 30269 20698
rect 30269 20646 30279 20698
rect 30303 20646 30333 20698
rect 30333 20646 30345 20698
rect 30345 20646 30359 20698
rect 30383 20646 30397 20698
rect 30397 20646 30409 20698
rect 30409 20646 30439 20698
rect 30463 20646 30473 20698
rect 30473 20646 30519 20698
rect 30223 20644 30279 20646
rect 30303 20644 30359 20646
rect 30383 20644 30439 20646
rect 30463 20644 30519 20646
rect 29826 19896 29882 19952
rect 28722 17856 28778 17912
rect 28814 17720 28870 17776
rect 28262 11756 28318 11792
rect 28262 11736 28264 11756
rect 28264 11736 28316 11756
rect 28316 11736 28318 11756
rect 30883 20154 30939 20156
rect 30963 20154 31019 20156
rect 31043 20154 31099 20156
rect 31123 20154 31179 20156
rect 30883 20102 30929 20154
rect 30929 20102 30939 20154
rect 30963 20102 30993 20154
rect 30993 20102 31005 20154
rect 31005 20102 31019 20154
rect 31043 20102 31057 20154
rect 31057 20102 31069 20154
rect 31069 20102 31099 20154
rect 31123 20102 31133 20154
rect 31133 20102 31179 20154
rect 30883 20100 30939 20102
rect 30963 20100 31019 20102
rect 31043 20100 31099 20102
rect 31123 20100 31179 20102
rect 30223 19610 30279 19612
rect 30303 19610 30359 19612
rect 30383 19610 30439 19612
rect 30463 19610 30519 19612
rect 30223 19558 30269 19610
rect 30269 19558 30279 19610
rect 30303 19558 30333 19610
rect 30333 19558 30345 19610
rect 30345 19558 30359 19610
rect 30383 19558 30397 19610
rect 30397 19558 30409 19610
rect 30409 19558 30439 19610
rect 30463 19558 30473 19610
rect 30473 19558 30519 19610
rect 30223 19556 30279 19558
rect 30303 19556 30359 19558
rect 30383 19556 30439 19558
rect 30463 19556 30519 19558
rect 29826 19080 29882 19136
rect 30223 18522 30279 18524
rect 30303 18522 30359 18524
rect 30383 18522 30439 18524
rect 30463 18522 30519 18524
rect 30223 18470 30269 18522
rect 30269 18470 30279 18522
rect 30303 18470 30333 18522
rect 30333 18470 30345 18522
rect 30345 18470 30359 18522
rect 30383 18470 30397 18522
rect 30397 18470 30409 18522
rect 30409 18470 30439 18522
rect 30463 18470 30473 18522
rect 30473 18470 30519 18522
rect 30223 18468 30279 18470
rect 30303 18468 30359 18470
rect 30383 18468 30439 18470
rect 30463 18468 30519 18470
rect 30883 19066 30939 19068
rect 30963 19066 31019 19068
rect 31043 19066 31099 19068
rect 31123 19066 31179 19068
rect 30883 19014 30929 19066
rect 30929 19014 30939 19066
rect 30963 19014 30993 19066
rect 30993 19014 31005 19066
rect 31005 19014 31019 19066
rect 31043 19014 31057 19066
rect 31057 19014 31069 19066
rect 31069 19014 31099 19066
rect 31123 19014 31133 19066
rect 31133 19014 31179 19066
rect 30883 19012 30939 19014
rect 30963 19012 31019 19014
rect 31043 19012 31099 19014
rect 31123 19012 31179 19014
rect 30223 17434 30279 17436
rect 30303 17434 30359 17436
rect 30383 17434 30439 17436
rect 30463 17434 30519 17436
rect 30223 17382 30269 17434
rect 30269 17382 30279 17434
rect 30303 17382 30333 17434
rect 30333 17382 30345 17434
rect 30345 17382 30359 17434
rect 30383 17382 30397 17434
rect 30397 17382 30409 17434
rect 30409 17382 30439 17434
rect 30463 17382 30473 17434
rect 30473 17382 30519 17434
rect 30223 17380 30279 17382
rect 30303 17380 30359 17382
rect 30383 17380 30439 17382
rect 30463 17380 30519 17382
rect 30883 17978 30939 17980
rect 30963 17978 31019 17980
rect 31043 17978 31099 17980
rect 31123 17978 31179 17980
rect 30883 17926 30929 17978
rect 30929 17926 30939 17978
rect 30963 17926 30993 17978
rect 30993 17926 31005 17978
rect 31005 17926 31019 17978
rect 31043 17926 31057 17978
rect 31057 17926 31069 17978
rect 31069 17926 31099 17978
rect 31123 17926 31133 17978
rect 31133 17926 31179 17978
rect 30883 17924 30939 17926
rect 30963 17924 31019 17926
rect 31043 17924 31099 17926
rect 31123 17924 31179 17926
rect 30883 16890 30939 16892
rect 30963 16890 31019 16892
rect 31043 16890 31099 16892
rect 31123 16890 31179 16892
rect 30883 16838 30929 16890
rect 30929 16838 30939 16890
rect 30963 16838 30993 16890
rect 30993 16838 31005 16890
rect 31005 16838 31019 16890
rect 31043 16838 31057 16890
rect 31057 16838 31069 16890
rect 31069 16838 31099 16890
rect 31123 16838 31133 16890
rect 31133 16838 31179 16890
rect 30883 16836 30939 16838
rect 30963 16836 31019 16838
rect 31043 16836 31099 16838
rect 31123 16836 31179 16838
rect 30223 16346 30279 16348
rect 30303 16346 30359 16348
rect 30383 16346 30439 16348
rect 30463 16346 30519 16348
rect 30223 16294 30269 16346
rect 30269 16294 30279 16346
rect 30303 16294 30333 16346
rect 30333 16294 30345 16346
rect 30345 16294 30359 16346
rect 30383 16294 30397 16346
rect 30397 16294 30409 16346
rect 30409 16294 30439 16346
rect 30463 16294 30473 16346
rect 30473 16294 30519 16346
rect 30223 16292 30279 16294
rect 30303 16292 30359 16294
rect 30383 16292 30439 16294
rect 30463 16292 30519 16294
rect 30883 15802 30939 15804
rect 30963 15802 31019 15804
rect 31043 15802 31099 15804
rect 31123 15802 31179 15804
rect 30883 15750 30929 15802
rect 30929 15750 30939 15802
rect 30963 15750 30993 15802
rect 30993 15750 31005 15802
rect 31005 15750 31019 15802
rect 31043 15750 31057 15802
rect 31057 15750 31069 15802
rect 31069 15750 31099 15802
rect 31123 15750 31133 15802
rect 31133 15750 31179 15802
rect 30883 15748 30939 15750
rect 30963 15748 31019 15750
rect 31043 15748 31099 15750
rect 31123 15748 31179 15750
rect 28998 14492 29000 14512
rect 29000 14492 29052 14512
rect 29052 14492 29054 14512
rect 28998 14456 29054 14492
rect 30223 15258 30279 15260
rect 30303 15258 30359 15260
rect 30383 15258 30439 15260
rect 30463 15258 30519 15260
rect 30223 15206 30269 15258
rect 30269 15206 30279 15258
rect 30303 15206 30333 15258
rect 30333 15206 30345 15258
rect 30345 15206 30359 15258
rect 30383 15206 30397 15258
rect 30397 15206 30409 15258
rect 30409 15206 30439 15258
rect 30463 15206 30473 15258
rect 30473 15206 30519 15258
rect 30223 15204 30279 15206
rect 30303 15204 30359 15206
rect 30383 15204 30439 15206
rect 30463 15204 30519 15206
rect 30883 14714 30939 14716
rect 30963 14714 31019 14716
rect 31043 14714 31099 14716
rect 31123 14714 31179 14716
rect 30883 14662 30929 14714
rect 30929 14662 30939 14714
rect 30963 14662 30993 14714
rect 30993 14662 31005 14714
rect 31005 14662 31019 14714
rect 31043 14662 31057 14714
rect 31057 14662 31069 14714
rect 31069 14662 31099 14714
rect 31123 14662 31133 14714
rect 31133 14662 31179 14714
rect 30883 14660 30939 14662
rect 30963 14660 31019 14662
rect 31043 14660 31099 14662
rect 31123 14660 31179 14662
rect 30223 14170 30279 14172
rect 30303 14170 30359 14172
rect 30383 14170 30439 14172
rect 30463 14170 30519 14172
rect 30223 14118 30269 14170
rect 30269 14118 30279 14170
rect 30303 14118 30333 14170
rect 30333 14118 30345 14170
rect 30345 14118 30359 14170
rect 30383 14118 30397 14170
rect 30397 14118 30409 14170
rect 30409 14118 30439 14170
rect 30463 14118 30473 14170
rect 30473 14118 30519 14170
rect 30223 14116 30279 14118
rect 30303 14116 30359 14118
rect 30383 14116 30439 14118
rect 30463 14116 30519 14118
rect 24858 9424 24914 9480
rect 24766 9152 24822 9208
rect 24858 6160 24914 6216
rect 25410 5752 25466 5808
rect 22994 2746 23050 2748
rect 23074 2746 23130 2748
rect 23154 2746 23210 2748
rect 23234 2746 23290 2748
rect 22994 2694 23040 2746
rect 23040 2694 23050 2746
rect 23074 2694 23104 2746
rect 23104 2694 23116 2746
rect 23116 2694 23130 2746
rect 23154 2694 23168 2746
rect 23168 2694 23180 2746
rect 23180 2694 23210 2746
rect 23234 2694 23244 2746
rect 23244 2694 23290 2746
rect 22994 2692 23050 2694
rect 23074 2692 23130 2694
rect 23154 2692 23210 2694
rect 23234 2692 23290 2694
rect 26238 8880 26294 8936
rect 26330 8628 26386 8664
rect 26330 8608 26332 8628
rect 26332 8608 26384 8628
rect 26384 8608 26386 8628
rect 26974 6296 27030 6352
rect 28170 9152 28226 9208
rect 28998 8372 29000 8392
rect 29000 8372 29052 8392
rect 29052 8372 29054 8392
rect 28630 6860 28686 6896
rect 28630 6840 28632 6860
rect 28632 6840 28684 6860
rect 28684 6840 28686 6860
rect 28998 8336 29054 8372
rect 30883 13626 30939 13628
rect 30963 13626 31019 13628
rect 31043 13626 31099 13628
rect 31123 13626 31179 13628
rect 30883 13574 30929 13626
rect 30929 13574 30939 13626
rect 30963 13574 30993 13626
rect 30993 13574 31005 13626
rect 31005 13574 31019 13626
rect 31043 13574 31057 13626
rect 31057 13574 31069 13626
rect 31069 13574 31099 13626
rect 31123 13574 31133 13626
rect 31133 13574 31179 13626
rect 30883 13572 30939 13574
rect 30963 13572 31019 13574
rect 31043 13572 31099 13574
rect 31123 13572 31179 13574
rect 30223 13082 30279 13084
rect 30303 13082 30359 13084
rect 30383 13082 30439 13084
rect 30463 13082 30519 13084
rect 30223 13030 30269 13082
rect 30269 13030 30279 13082
rect 30303 13030 30333 13082
rect 30333 13030 30345 13082
rect 30345 13030 30359 13082
rect 30383 13030 30397 13082
rect 30397 13030 30409 13082
rect 30409 13030 30439 13082
rect 30463 13030 30473 13082
rect 30473 13030 30519 13082
rect 30223 13028 30279 13030
rect 30303 13028 30359 13030
rect 30383 13028 30439 13030
rect 30463 13028 30519 13030
rect 30883 12538 30939 12540
rect 30963 12538 31019 12540
rect 31043 12538 31099 12540
rect 31123 12538 31179 12540
rect 30883 12486 30929 12538
rect 30929 12486 30939 12538
rect 30963 12486 30993 12538
rect 30993 12486 31005 12538
rect 31005 12486 31019 12538
rect 31043 12486 31057 12538
rect 31057 12486 31069 12538
rect 31069 12486 31099 12538
rect 31123 12486 31133 12538
rect 31133 12486 31179 12538
rect 30883 12484 30939 12486
rect 30963 12484 31019 12486
rect 31043 12484 31099 12486
rect 31123 12484 31179 12486
rect 30223 11994 30279 11996
rect 30303 11994 30359 11996
rect 30383 11994 30439 11996
rect 30463 11994 30519 11996
rect 30223 11942 30269 11994
rect 30269 11942 30279 11994
rect 30303 11942 30333 11994
rect 30333 11942 30345 11994
rect 30345 11942 30359 11994
rect 30383 11942 30397 11994
rect 30397 11942 30409 11994
rect 30409 11942 30439 11994
rect 30463 11942 30473 11994
rect 30473 11942 30519 11994
rect 30223 11940 30279 11942
rect 30303 11940 30359 11942
rect 30383 11940 30439 11942
rect 30463 11940 30519 11942
rect 31942 12280 31998 12336
rect 30883 11450 30939 11452
rect 30963 11450 31019 11452
rect 31043 11450 31099 11452
rect 31123 11450 31179 11452
rect 30883 11398 30929 11450
rect 30929 11398 30939 11450
rect 30963 11398 30993 11450
rect 30993 11398 31005 11450
rect 31005 11398 31019 11450
rect 31043 11398 31057 11450
rect 31057 11398 31069 11450
rect 31069 11398 31099 11450
rect 31123 11398 31133 11450
rect 31133 11398 31179 11450
rect 30883 11396 30939 11398
rect 30963 11396 31019 11398
rect 31043 11396 31099 11398
rect 31123 11396 31179 11398
rect 30223 10906 30279 10908
rect 30303 10906 30359 10908
rect 30383 10906 30439 10908
rect 30463 10906 30519 10908
rect 30223 10854 30269 10906
rect 30269 10854 30279 10906
rect 30303 10854 30333 10906
rect 30333 10854 30345 10906
rect 30345 10854 30359 10906
rect 30383 10854 30397 10906
rect 30397 10854 30409 10906
rect 30409 10854 30439 10906
rect 30463 10854 30473 10906
rect 30473 10854 30519 10906
rect 30223 10852 30279 10854
rect 30303 10852 30359 10854
rect 30383 10852 30439 10854
rect 30463 10852 30519 10854
rect 30223 9818 30279 9820
rect 30303 9818 30359 9820
rect 30383 9818 30439 9820
rect 30463 9818 30519 9820
rect 30223 9766 30269 9818
rect 30269 9766 30279 9818
rect 30303 9766 30333 9818
rect 30333 9766 30345 9818
rect 30345 9766 30359 9818
rect 30383 9766 30397 9818
rect 30397 9766 30409 9818
rect 30409 9766 30439 9818
rect 30463 9766 30473 9818
rect 30473 9766 30519 9818
rect 30223 9764 30279 9766
rect 30303 9764 30359 9766
rect 30383 9764 30439 9766
rect 30463 9764 30519 9766
rect 30883 10362 30939 10364
rect 30963 10362 31019 10364
rect 31043 10362 31099 10364
rect 31123 10362 31179 10364
rect 30883 10310 30929 10362
rect 30929 10310 30939 10362
rect 30963 10310 30993 10362
rect 30993 10310 31005 10362
rect 31005 10310 31019 10362
rect 31043 10310 31057 10362
rect 31057 10310 31069 10362
rect 31069 10310 31099 10362
rect 31123 10310 31133 10362
rect 31133 10310 31179 10362
rect 30883 10308 30939 10310
rect 30963 10308 31019 10310
rect 31043 10308 31099 10310
rect 31123 10308 31179 10310
rect 30883 9274 30939 9276
rect 30963 9274 31019 9276
rect 31043 9274 31099 9276
rect 31123 9274 31179 9276
rect 30883 9222 30929 9274
rect 30929 9222 30939 9274
rect 30963 9222 30993 9274
rect 30993 9222 31005 9274
rect 31005 9222 31019 9274
rect 31043 9222 31057 9274
rect 31057 9222 31069 9274
rect 31069 9222 31099 9274
rect 31123 9222 31133 9274
rect 31133 9222 31179 9274
rect 30883 9220 30939 9222
rect 30963 9220 31019 9222
rect 31043 9220 31099 9222
rect 31123 9220 31179 9222
rect 30223 8730 30279 8732
rect 30303 8730 30359 8732
rect 30383 8730 30439 8732
rect 30463 8730 30519 8732
rect 30223 8678 30269 8730
rect 30269 8678 30279 8730
rect 30303 8678 30333 8730
rect 30333 8678 30345 8730
rect 30345 8678 30359 8730
rect 30383 8678 30397 8730
rect 30397 8678 30409 8730
rect 30409 8678 30439 8730
rect 30463 8678 30473 8730
rect 30473 8678 30519 8730
rect 30223 8676 30279 8678
rect 30303 8676 30359 8678
rect 30383 8676 30439 8678
rect 30463 8676 30519 8678
rect 29274 8064 29330 8120
rect 30562 8064 30618 8120
rect 30223 7642 30279 7644
rect 30303 7642 30359 7644
rect 30383 7642 30439 7644
rect 30463 7642 30519 7644
rect 30223 7590 30269 7642
rect 30269 7590 30279 7642
rect 30303 7590 30333 7642
rect 30333 7590 30345 7642
rect 30345 7590 30359 7642
rect 30383 7590 30397 7642
rect 30397 7590 30409 7642
rect 30409 7590 30439 7642
rect 30463 7590 30473 7642
rect 30473 7590 30519 7642
rect 30223 7588 30279 7590
rect 30303 7588 30359 7590
rect 30383 7588 30439 7590
rect 30463 7588 30519 7590
rect 30883 8186 30939 8188
rect 30963 8186 31019 8188
rect 31043 8186 31099 8188
rect 31123 8186 31179 8188
rect 30883 8134 30929 8186
rect 30929 8134 30939 8186
rect 30963 8134 30993 8186
rect 30993 8134 31005 8186
rect 31005 8134 31019 8186
rect 31043 8134 31057 8186
rect 31057 8134 31069 8186
rect 31069 8134 31099 8186
rect 31123 8134 31133 8186
rect 31133 8134 31179 8186
rect 30883 8132 30939 8134
rect 30963 8132 31019 8134
rect 31043 8132 31099 8134
rect 31123 8132 31179 8134
rect 28170 5652 28172 5672
rect 28172 5652 28224 5672
rect 28224 5652 28226 5672
rect 28170 5616 28226 5652
rect 30883 7098 30939 7100
rect 30963 7098 31019 7100
rect 31043 7098 31099 7100
rect 31123 7098 31179 7100
rect 30883 7046 30929 7098
rect 30929 7046 30939 7098
rect 30963 7046 30993 7098
rect 30993 7046 31005 7098
rect 31005 7046 31019 7098
rect 31043 7046 31057 7098
rect 31057 7046 31069 7098
rect 31069 7046 31099 7098
rect 31123 7046 31133 7098
rect 31133 7046 31179 7098
rect 30883 7044 30939 7046
rect 30963 7044 31019 7046
rect 31043 7044 31099 7046
rect 31123 7044 31179 7046
rect 30223 6554 30279 6556
rect 30303 6554 30359 6556
rect 30383 6554 30439 6556
rect 30463 6554 30519 6556
rect 30223 6502 30269 6554
rect 30269 6502 30279 6554
rect 30303 6502 30333 6554
rect 30333 6502 30345 6554
rect 30345 6502 30359 6554
rect 30383 6502 30397 6554
rect 30397 6502 30409 6554
rect 30409 6502 30439 6554
rect 30463 6502 30473 6554
rect 30473 6502 30519 6554
rect 30223 6500 30279 6502
rect 30303 6500 30359 6502
rect 30383 6500 30439 6502
rect 30463 6500 30519 6502
rect 30883 6010 30939 6012
rect 30963 6010 31019 6012
rect 31043 6010 31099 6012
rect 31123 6010 31179 6012
rect 30883 5958 30929 6010
rect 30929 5958 30939 6010
rect 30963 5958 30993 6010
rect 30993 5958 31005 6010
rect 31005 5958 31019 6010
rect 31043 5958 31057 6010
rect 31057 5958 31069 6010
rect 31069 5958 31099 6010
rect 31123 5958 31133 6010
rect 31133 5958 31179 6010
rect 30883 5956 30939 5958
rect 30963 5956 31019 5958
rect 31043 5956 31099 5958
rect 31123 5956 31179 5958
rect 30223 5466 30279 5468
rect 30303 5466 30359 5468
rect 30383 5466 30439 5468
rect 30463 5466 30519 5468
rect 30223 5414 30269 5466
rect 30269 5414 30279 5466
rect 30303 5414 30333 5466
rect 30333 5414 30345 5466
rect 30345 5414 30359 5466
rect 30383 5414 30397 5466
rect 30397 5414 30409 5466
rect 30409 5414 30439 5466
rect 30463 5414 30473 5466
rect 30473 5414 30519 5466
rect 30223 5412 30279 5414
rect 30303 5412 30359 5414
rect 30383 5412 30439 5414
rect 30463 5412 30519 5414
rect 30883 4922 30939 4924
rect 30963 4922 31019 4924
rect 31043 4922 31099 4924
rect 31123 4922 31179 4924
rect 30883 4870 30929 4922
rect 30929 4870 30939 4922
rect 30963 4870 30993 4922
rect 30993 4870 31005 4922
rect 31005 4870 31019 4922
rect 31043 4870 31057 4922
rect 31057 4870 31069 4922
rect 31069 4870 31099 4922
rect 31123 4870 31133 4922
rect 31133 4870 31179 4922
rect 30883 4868 30939 4870
rect 30963 4868 31019 4870
rect 31043 4868 31099 4870
rect 31123 4868 31179 4870
rect 30223 4378 30279 4380
rect 30303 4378 30359 4380
rect 30383 4378 30439 4380
rect 30463 4378 30519 4380
rect 30223 4326 30269 4378
rect 30269 4326 30279 4378
rect 30303 4326 30333 4378
rect 30333 4326 30345 4378
rect 30345 4326 30359 4378
rect 30383 4326 30397 4378
rect 30397 4326 30409 4378
rect 30409 4326 30439 4378
rect 30463 4326 30473 4378
rect 30473 4326 30519 4378
rect 30223 4324 30279 4326
rect 30303 4324 30359 4326
rect 30383 4324 30439 4326
rect 30463 4324 30519 4326
rect 30883 3834 30939 3836
rect 30963 3834 31019 3836
rect 31043 3834 31099 3836
rect 31123 3834 31179 3836
rect 30883 3782 30929 3834
rect 30929 3782 30939 3834
rect 30963 3782 30993 3834
rect 30993 3782 31005 3834
rect 31005 3782 31019 3834
rect 31043 3782 31057 3834
rect 31057 3782 31069 3834
rect 31069 3782 31099 3834
rect 31123 3782 31133 3834
rect 31133 3782 31179 3834
rect 30883 3780 30939 3782
rect 30963 3780 31019 3782
rect 31043 3780 31099 3782
rect 31123 3780 31179 3782
rect 30223 3290 30279 3292
rect 30303 3290 30359 3292
rect 30383 3290 30439 3292
rect 30463 3290 30519 3292
rect 30223 3238 30269 3290
rect 30269 3238 30279 3290
rect 30303 3238 30333 3290
rect 30333 3238 30345 3290
rect 30345 3238 30359 3290
rect 30383 3238 30397 3290
rect 30397 3238 30409 3290
rect 30409 3238 30439 3290
rect 30463 3238 30473 3290
rect 30473 3238 30519 3290
rect 30223 3236 30279 3238
rect 30303 3236 30359 3238
rect 30383 3236 30439 3238
rect 30463 3236 30519 3238
rect 32402 19896 32458 19952
rect 33046 25880 33102 25936
rect 33782 19760 33838 19816
rect 33046 17040 33102 17096
rect 32678 12280 32734 12336
rect 33782 9016 33838 9072
rect 33782 8508 33784 8528
rect 33784 8508 33836 8528
rect 33836 8508 33838 8528
rect 33782 8472 33838 8508
rect 32218 5616 32274 5672
rect 35162 29960 35218 30016
rect 35162 27240 35218 27296
rect 34702 23840 34758 23896
rect 35162 22516 35164 22536
rect 35164 22516 35216 22536
rect 35216 22516 35218 22536
rect 35162 22480 35218 22516
rect 34886 21120 34942 21176
rect 34518 18400 34574 18456
rect 34886 15680 34942 15736
rect 35162 13640 35218 13696
rect 34426 12280 34482 12336
rect 34886 10920 34942 10976
rect 34426 9560 34482 9616
rect 34426 8200 34482 8256
rect 34702 6860 34758 6896
rect 34702 6840 34704 6860
rect 34704 6840 34756 6860
rect 34756 6840 34758 6860
rect 34058 5752 34114 5808
rect 34886 5480 34942 5536
rect 34702 4120 34758 4176
rect 30883 2746 30939 2748
rect 30963 2746 31019 2748
rect 31043 2746 31099 2748
rect 31123 2746 31179 2748
rect 30883 2694 30929 2746
rect 30929 2694 30939 2746
rect 30963 2694 30993 2746
rect 30993 2694 31005 2746
rect 31005 2694 31019 2746
rect 31043 2694 31057 2746
rect 31057 2694 31069 2746
rect 31069 2694 31099 2746
rect 31123 2694 31133 2746
rect 31133 2694 31179 2746
rect 30883 2692 30939 2694
rect 30963 2692 31019 2694
rect 31043 2692 31099 2694
rect 31123 2692 31179 2694
rect 33046 856 33102 912
rect 34426 2080 34482 2136
<< metal3 >>
rect 0 36138 800 36168
rect 3785 36138 3851 36141
rect 0 36136 3851 36138
rect 0 36080 3790 36136
rect 3846 36080 3851 36136
rect 0 36078 3851 36080
rect 0 36048 800 36078
rect 3785 36075 3851 36078
rect 33777 35458 33843 35461
rect 36302 35458 37102 35488
rect 33777 35456 37102 35458
rect 33777 35400 33782 35456
rect 33838 35400 37102 35456
rect 33777 35398 37102 35400
rect 33777 35395 33843 35398
rect 36302 35368 37102 35398
rect 0 34778 800 34808
rect 3049 34778 3115 34781
rect 0 34776 3115 34778
rect 0 34720 3054 34776
rect 3110 34720 3115 34776
rect 0 34718 3115 34720
rect 0 34688 800 34718
rect 3049 34715 3115 34718
rect 7206 34304 7522 34305
rect 7206 34240 7212 34304
rect 7276 34240 7292 34304
rect 7356 34240 7372 34304
rect 7436 34240 7452 34304
rect 7516 34240 7522 34304
rect 7206 34239 7522 34240
rect 15095 34304 15411 34305
rect 15095 34240 15101 34304
rect 15165 34240 15181 34304
rect 15245 34240 15261 34304
rect 15325 34240 15341 34304
rect 15405 34240 15411 34304
rect 15095 34239 15411 34240
rect 22984 34304 23300 34305
rect 22984 34240 22990 34304
rect 23054 34240 23070 34304
rect 23134 34240 23150 34304
rect 23214 34240 23230 34304
rect 23294 34240 23300 34304
rect 22984 34239 23300 34240
rect 30873 34304 31189 34305
rect 30873 34240 30879 34304
rect 30943 34240 30959 34304
rect 31023 34240 31039 34304
rect 31103 34240 31119 34304
rect 31183 34240 31189 34304
rect 30873 34239 31189 34240
rect 33041 34098 33107 34101
rect 36302 34098 37102 34128
rect 33041 34096 37102 34098
rect 33041 34040 33046 34096
rect 33102 34040 37102 34096
rect 33041 34038 37102 34040
rect 33041 34035 33107 34038
rect 36302 34008 37102 34038
rect 6546 33760 6862 33761
rect 6546 33696 6552 33760
rect 6616 33696 6632 33760
rect 6696 33696 6712 33760
rect 6776 33696 6792 33760
rect 6856 33696 6862 33760
rect 6546 33695 6862 33696
rect 14435 33760 14751 33761
rect 14435 33696 14441 33760
rect 14505 33696 14521 33760
rect 14585 33696 14601 33760
rect 14665 33696 14681 33760
rect 14745 33696 14751 33760
rect 14435 33695 14751 33696
rect 22324 33760 22640 33761
rect 22324 33696 22330 33760
rect 22394 33696 22410 33760
rect 22474 33696 22490 33760
rect 22554 33696 22570 33760
rect 22634 33696 22640 33760
rect 22324 33695 22640 33696
rect 30213 33760 30529 33761
rect 30213 33696 30219 33760
rect 30283 33696 30299 33760
rect 30363 33696 30379 33760
rect 30443 33696 30459 33760
rect 30523 33696 30529 33760
rect 30213 33695 30529 33696
rect 0 33418 800 33448
rect 3233 33418 3299 33421
rect 0 33416 3299 33418
rect 0 33360 3238 33416
rect 3294 33360 3299 33416
rect 0 33358 3299 33360
rect 0 33328 800 33358
rect 3233 33355 3299 33358
rect 10869 33284 10935 33285
rect 10869 33280 10916 33284
rect 10980 33282 10986 33284
rect 11421 33282 11487 33285
rect 13077 33282 13143 33285
rect 10869 33224 10874 33280
rect 10869 33220 10916 33224
rect 10980 33222 11026 33282
rect 11421 33280 13143 33282
rect 11421 33224 11426 33280
rect 11482 33224 13082 33280
rect 13138 33224 13143 33280
rect 11421 33222 13143 33224
rect 10980 33220 10986 33222
rect 10869 33219 10935 33220
rect 11421 33219 11487 33222
rect 13077 33219 13143 33222
rect 19057 33282 19123 33285
rect 21541 33284 21607 33285
rect 19190 33282 19196 33284
rect 19057 33280 19196 33282
rect 19057 33224 19062 33280
rect 19118 33224 19196 33280
rect 19057 33222 19196 33224
rect 19057 33219 19123 33222
rect 19190 33220 19196 33222
rect 19260 33220 19266 33284
rect 21541 33280 21588 33284
rect 21652 33282 21658 33284
rect 21541 33224 21546 33280
rect 21541 33220 21588 33224
rect 21652 33222 21698 33282
rect 21652 33220 21658 33222
rect 21541 33219 21607 33220
rect 7206 33216 7522 33217
rect 7206 33152 7212 33216
rect 7276 33152 7292 33216
rect 7356 33152 7372 33216
rect 7436 33152 7452 33216
rect 7516 33152 7522 33216
rect 7206 33151 7522 33152
rect 15095 33216 15411 33217
rect 15095 33152 15101 33216
rect 15165 33152 15181 33216
rect 15245 33152 15261 33216
rect 15325 33152 15341 33216
rect 15405 33152 15411 33216
rect 15095 33151 15411 33152
rect 22984 33216 23300 33217
rect 22984 33152 22990 33216
rect 23054 33152 23070 33216
rect 23134 33152 23150 33216
rect 23214 33152 23230 33216
rect 23294 33152 23300 33216
rect 22984 33151 23300 33152
rect 30873 33216 31189 33217
rect 30873 33152 30879 33216
rect 30943 33152 30959 33216
rect 31023 33152 31039 33216
rect 31103 33152 31119 33216
rect 31183 33152 31189 33216
rect 30873 33151 31189 33152
rect 11605 33146 11671 33149
rect 12198 33146 12204 33148
rect 11605 33144 12204 33146
rect 11605 33088 11610 33144
rect 11666 33088 12204 33144
rect 11605 33086 12204 33088
rect 11605 33083 11671 33086
rect 12198 33084 12204 33086
rect 12268 33084 12274 33148
rect 12065 33010 12131 33013
rect 13997 33010 14063 33013
rect 12065 33008 14063 33010
rect 12065 32952 12070 33008
rect 12126 32952 14002 33008
rect 14058 32952 14063 33008
rect 12065 32950 14063 32952
rect 12065 32947 12131 32950
rect 13997 32947 14063 32950
rect 11053 32874 11119 32877
rect 12065 32874 12131 32877
rect 15561 32874 15627 32877
rect 11053 32872 15627 32874
rect 11053 32816 11058 32872
rect 11114 32816 12070 32872
rect 12126 32816 15566 32872
rect 15622 32816 15627 32872
rect 11053 32814 15627 32816
rect 11053 32811 11119 32814
rect 12065 32811 12131 32814
rect 15561 32811 15627 32814
rect 34881 32738 34947 32741
rect 36302 32738 37102 32768
rect 34881 32736 37102 32738
rect 34881 32680 34886 32736
rect 34942 32680 37102 32736
rect 34881 32678 37102 32680
rect 34881 32675 34947 32678
rect 6546 32672 6862 32673
rect 6546 32608 6552 32672
rect 6616 32608 6632 32672
rect 6696 32608 6712 32672
rect 6776 32608 6792 32672
rect 6856 32608 6862 32672
rect 6546 32607 6862 32608
rect 14435 32672 14751 32673
rect 14435 32608 14441 32672
rect 14505 32608 14521 32672
rect 14585 32608 14601 32672
rect 14665 32608 14681 32672
rect 14745 32608 14751 32672
rect 14435 32607 14751 32608
rect 22324 32672 22640 32673
rect 22324 32608 22330 32672
rect 22394 32608 22410 32672
rect 22474 32608 22490 32672
rect 22554 32608 22570 32672
rect 22634 32608 22640 32672
rect 22324 32607 22640 32608
rect 30213 32672 30529 32673
rect 30213 32608 30219 32672
rect 30283 32608 30299 32672
rect 30363 32608 30379 32672
rect 30443 32608 30459 32672
rect 30523 32608 30529 32672
rect 36302 32648 37102 32678
rect 30213 32607 30529 32608
rect 13261 32466 13327 32469
rect 15009 32466 15075 32469
rect 13261 32464 15075 32466
rect 13261 32408 13266 32464
rect 13322 32408 15014 32464
rect 15070 32408 15075 32464
rect 13261 32406 15075 32408
rect 13261 32403 13327 32406
rect 15009 32403 15075 32406
rect 4429 32330 4495 32333
rect 18781 32330 18847 32333
rect 4429 32328 18847 32330
rect 4429 32272 4434 32328
rect 4490 32272 18786 32328
rect 18842 32272 18847 32328
rect 4429 32270 18847 32272
rect 4429 32267 4495 32270
rect 18781 32267 18847 32270
rect 7206 32128 7522 32129
rect 7206 32064 7212 32128
rect 7276 32064 7292 32128
rect 7356 32064 7372 32128
rect 7436 32064 7452 32128
rect 7516 32064 7522 32128
rect 7206 32063 7522 32064
rect 15095 32128 15411 32129
rect 15095 32064 15101 32128
rect 15165 32064 15181 32128
rect 15245 32064 15261 32128
rect 15325 32064 15341 32128
rect 15405 32064 15411 32128
rect 15095 32063 15411 32064
rect 22984 32128 23300 32129
rect 22984 32064 22990 32128
rect 23054 32064 23070 32128
rect 23134 32064 23150 32128
rect 23214 32064 23230 32128
rect 23294 32064 23300 32128
rect 22984 32063 23300 32064
rect 30873 32128 31189 32129
rect 30873 32064 30879 32128
rect 30943 32064 30959 32128
rect 31023 32064 31039 32128
rect 31103 32064 31119 32128
rect 31183 32064 31189 32128
rect 30873 32063 31189 32064
rect 6546 31584 6862 31585
rect 6546 31520 6552 31584
rect 6616 31520 6632 31584
rect 6696 31520 6712 31584
rect 6776 31520 6792 31584
rect 6856 31520 6862 31584
rect 6546 31519 6862 31520
rect 14435 31584 14751 31585
rect 14435 31520 14441 31584
rect 14505 31520 14521 31584
rect 14585 31520 14601 31584
rect 14665 31520 14681 31584
rect 14745 31520 14751 31584
rect 14435 31519 14751 31520
rect 22324 31584 22640 31585
rect 22324 31520 22330 31584
rect 22394 31520 22410 31584
rect 22474 31520 22490 31584
rect 22554 31520 22570 31584
rect 22634 31520 22640 31584
rect 22324 31519 22640 31520
rect 30213 31584 30529 31585
rect 30213 31520 30219 31584
rect 30283 31520 30299 31584
rect 30363 31520 30379 31584
rect 30443 31520 30459 31584
rect 30523 31520 30529 31584
rect 30213 31519 30529 31520
rect 0 31378 800 31408
rect 3233 31378 3299 31381
rect 0 31376 3299 31378
rect 0 31320 3238 31376
rect 3294 31320 3299 31376
rect 0 31318 3299 31320
rect 0 31288 800 31318
rect 3233 31315 3299 31318
rect 32121 31378 32187 31381
rect 36302 31378 37102 31408
rect 32121 31376 37102 31378
rect 32121 31320 32126 31376
rect 32182 31320 37102 31376
rect 32121 31318 37102 31320
rect 32121 31315 32187 31318
rect 36302 31288 37102 31318
rect 7206 31040 7522 31041
rect 7206 30976 7212 31040
rect 7276 30976 7292 31040
rect 7356 30976 7372 31040
rect 7436 30976 7452 31040
rect 7516 30976 7522 31040
rect 7206 30975 7522 30976
rect 15095 31040 15411 31041
rect 15095 30976 15101 31040
rect 15165 30976 15181 31040
rect 15245 30976 15261 31040
rect 15325 30976 15341 31040
rect 15405 30976 15411 31040
rect 15095 30975 15411 30976
rect 22984 31040 23300 31041
rect 22984 30976 22990 31040
rect 23054 30976 23070 31040
rect 23134 30976 23150 31040
rect 23214 30976 23230 31040
rect 23294 30976 23300 31040
rect 22984 30975 23300 30976
rect 30873 31040 31189 31041
rect 30873 30976 30879 31040
rect 30943 30976 30959 31040
rect 31023 30976 31039 31040
rect 31103 30976 31119 31040
rect 31183 30976 31189 31040
rect 30873 30975 31189 30976
rect 6546 30496 6862 30497
rect 6546 30432 6552 30496
rect 6616 30432 6632 30496
rect 6696 30432 6712 30496
rect 6776 30432 6792 30496
rect 6856 30432 6862 30496
rect 6546 30431 6862 30432
rect 14435 30496 14751 30497
rect 14435 30432 14441 30496
rect 14505 30432 14521 30496
rect 14585 30432 14601 30496
rect 14665 30432 14681 30496
rect 14745 30432 14751 30496
rect 14435 30431 14751 30432
rect 22324 30496 22640 30497
rect 22324 30432 22330 30496
rect 22394 30432 22410 30496
rect 22474 30432 22490 30496
rect 22554 30432 22570 30496
rect 22634 30432 22640 30496
rect 22324 30431 22640 30432
rect 30213 30496 30529 30497
rect 30213 30432 30219 30496
rect 30283 30432 30299 30496
rect 30363 30432 30379 30496
rect 30443 30432 30459 30496
rect 30523 30432 30529 30496
rect 30213 30431 30529 30432
rect 0 30018 800 30048
rect 1301 30018 1367 30021
rect 0 30016 1367 30018
rect 0 29960 1306 30016
rect 1362 29960 1367 30016
rect 0 29958 1367 29960
rect 0 29928 800 29958
rect 1301 29955 1367 29958
rect 35157 30018 35223 30021
rect 36302 30018 37102 30048
rect 35157 30016 37102 30018
rect 35157 29960 35162 30016
rect 35218 29960 37102 30016
rect 35157 29958 37102 29960
rect 35157 29955 35223 29958
rect 7206 29952 7522 29953
rect 7206 29888 7212 29952
rect 7276 29888 7292 29952
rect 7356 29888 7372 29952
rect 7436 29888 7452 29952
rect 7516 29888 7522 29952
rect 7206 29887 7522 29888
rect 15095 29952 15411 29953
rect 15095 29888 15101 29952
rect 15165 29888 15181 29952
rect 15245 29888 15261 29952
rect 15325 29888 15341 29952
rect 15405 29888 15411 29952
rect 15095 29887 15411 29888
rect 22984 29952 23300 29953
rect 22984 29888 22990 29952
rect 23054 29888 23070 29952
rect 23134 29888 23150 29952
rect 23214 29888 23230 29952
rect 23294 29888 23300 29952
rect 22984 29887 23300 29888
rect 30873 29952 31189 29953
rect 30873 29888 30879 29952
rect 30943 29888 30959 29952
rect 31023 29888 31039 29952
rect 31103 29888 31119 29952
rect 31183 29888 31189 29952
rect 36302 29928 37102 29958
rect 30873 29887 31189 29888
rect 6546 29408 6862 29409
rect 6546 29344 6552 29408
rect 6616 29344 6632 29408
rect 6696 29344 6712 29408
rect 6776 29344 6792 29408
rect 6856 29344 6862 29408
rect 6546 29343 6862 29344
rect 14435 29408 14751 29409
rect 14435 29344 14441 29408
rect 14505 29344 14521 29408
rect 14585 29344 14601 29408
rect 14665 29344 14681 29408
rect 14745 29344 14751 29408
rect 14435 29343 14751 29344
rect 22324 29408 22640 29409
rect 22324 29344 22330 29408
rect 22394 29344 22410 29408
rect 22474 29344 22490 29408
rect 22554 29344 22570 29408
rect 22634 29344 22640 29408
rect 22324 29343 22640 29344
rect 30213 29408 30529 29409
rect 30213 29344 30219 29408
rect 30283 29344 30299 29408
rect 30363 29344 30379 29408
rect 30443 29344 30459 29408
rect 30523 29344 30529 29408
rect 30213 29343 30529 29344
rect 13077 29202 13143 29205
rect 16481 29202 16547 29205
rect 13077 29200 16547 29202
rect 13077 29144 13082 29200
rect 13138 29144 16486 29200
rect 16542 29144 16547 29200
rect 13077 29142 16547 29144
rect 13077 29139 13143 29142
rect 16481 29139 16547 29142
rect 27705 29066 27771 29069
rect 27838 29066 27844 29068
rect 27705 29064 27844 29066
rect 27705 29008 27710 29064
rect 27766 29008 27844 29064
rect 27705 29006 27844 29008
rect 27705 29003 27771 29006
rect 27838 29004 27844 29006
rect 27908 29004 27914 29068
rect 7206 28864 7522 28865
rect 7206 28800 7212 28864
rect 7276 28800 7292 28864
rect 7356 28800 7372 28864
rect 7436 28800 7452 28864
rect 7516 28800 7522 28864
rect 7206 28799 7522 28800
rect 15095 28864 15411 28865
rect 15095 28800 15101 28864
rect 15165 28800 15181 28864
rect 15245 28800 15261 28864
rect 15325 28800 15341 28864
rect 15405 28800 15411 28864
rect 15095 28799 15411 28800
rect 22984 28864 23300 28865
rect 22984 28800 22990 28864
rect 23054 28800 23070 28864
rect 23134 28800 23150 28864
rect 23214 28800 23230 28864
rect 23294 28800 23300 28864
rect 22984 28799 23300 28800
rect 30873 28864 31189 28865
rect 30873 28800 30879 28864
rect 30943 28800 30959 28864
rect 31023 28800 31039 28864
rect 31103 28800 31119 28864
rect 31183 28800 31189 28864
rect 30873 28799 31189 28800
rect 0 28658 800 28688
rect 1301 28658 1367 28661
rect 0 28656 1367 28658
rect 0 28600 1306 28656
rect 1362 28600 1367 28656
rect 0 28598 1367 28600
rect 0 28568 800 28598
rect 1301 28595 1367 28598
rect 33777 28658 33843 28661
rect 36302 28658 37102 28688
rect 33777 28656 37102 28658
rect 33777 28600 33782 28656
rect 33838 28600 37102 28656
rect 33777 28598 37102 28600
rect 33777 28595 33843 28598
rect 36302 28568 37102 28598
rect 6546 28320 6862 28321
rect 6546 28256 6552 28320
rect 6616 28256 6632 28320
rect 6696 28256 6712 28320
rect 6776 28256 6792 28320
rect 6856 28256 6862 28320
rect 6546 28255 6862 28256
rect 14435 28320 14751 28321
rect 14435 28256 14441 28320
rect 14505 28256 14521 28320
rect 14585 28256 14601 28320
rect 14665 28256 14681 28320
rect 14745 28256 14751 28320
rect 14435 28255 14751 28256
rect 22324 28320 22640 28321
rect 22324 28256 22330 28320
rect 22394 28256 22410 28320
rect 22474 28256 22490 28320
rect 22554 28256 22570 28320
rect 22634 28256 22640 28320
rect 22324 28255 22640 28256
rect 30213 28320 30529 28321
rect 30213 28256 30219 28320
rect 30283 28256 30299 28320
rect 30363 28256 30379 28320
rect 30443 28256 30459 28320
rect 30523 28256 30529 28320
rect 30213 28255 30529 28256
rect 19609 28114 19675 28117
rect 25037 28114 25103 28117
rect 19609 28112 25103 28114
rect 19609 28056 19614 28112
rect 19670 28056 25042 28112
rect 25098 28056 25103 28112
rect 19609 28054 25103 28056
rect 19609 28051 19675 28054
rect 25037 28051 25103 28054
rect 20069 27978 20135 27981
rect 28901 27978 28967 27981
rect 20069 27976 28967 27978
rect 20069 27920 20074 27976
rect 20130 27920 28906 27976
rect 28962 27920 28967 27976
rect 20069 27918 28967 27920
rect 20069 27915 20135 27918
rect 28901 27915 28967 27918
rect 7206 27776 7522 27777
rect 7206 27712 7212 27776
rect 7276 27712 7292 27776
rect 7356 27712 7372 27776
rect 7436 27712 7452 27776
rect 7516 27712 7522 27776
rect 7206 27711 7522 27712
rect 15095 27776 15411 27777
rect 15095 27712 15101 27776
rect 15165 27712 15181 27776
rect 15245 27712 15261 27776
rect 15325 27712 15341 27776
rect 15405 27712 15411 27776
rect 15095 27711 15411 27712
rect 22984 27776 23300 27777
rect 22984 27712 22990 27776
rect 23054 27712 23070 27776
rect 23134 27712 23150 27776
rect 23214 27712 23230 27776
rect 23294 27712 23300 27776
rect 22984 27711 23300 27712
rect 30873 27776 31189 27777
rect 30873 27712 30879 27776
rect 30943 27712 30959 27776
rect 31023 27712 31039 27776
rect 31103 27712 31119 27776
rect 31183 27712 31189 27776
rect 30873 27711 31189 27712
rect 27981 27570 28047 27573
rect 33041 27570 33107 27573
rect 27981 27568 33107 27570
rect 27981 27512 27986 27568
rect 28042 27512 33046 27568
rect 33102 27512 33107 27568
rect 27981 27510 33107 27512
rect 27981 27507 28047 27510
rect 33041 27507 33107 27510
rect 0 27298 800 27328
rect 1301 27298 1367 27301
rect 0 27296 1367 27298
rect 0 27240 1306 27296
rect 1362 27240 1367 27296
rect 0 27238 1367 27240
rect 0 27208 800 27238
rect 1301 27235 1367 27238
rect 35157 27298 35223 27301
rect 36302 27298 37102 27328
rect 35157 27296 37102 27298
rect 35157 27240 35162 27296
rect 35218 27240 37102 27296
rect 35157 27238 37102 27240
rect 35157 27235 35223 27238
rect 6546 27232 6862 27233
rect 6546 27168 6552 27232
rect 6616 27168 6632 27232
rect 6696 27168 6712 27232
rect 6776 27168 6792 27232
rect 6856 27168 6862 27232
rect 6546 27167 6862 27168
rect 14435 27232 14751 27233
rect 14435 27168 14441 27232
rect 14505 27168 14521 27232
rect 14585 27168 14601 27232
rect 14665 27168 14681 27232
rect 14745 27168 14751 27232
rect 14435 27167 14751 27168
rect 22324 27232 22640 27233
rect 22324 27168 22330 27232
rect 22394 27168 22410 27232
rect 22474 27168 22490 27232
rect 22554 27168 22570 27232
rect 22634 27168 22640 27232
rect 22324 27167 22640 27168
rect 30213 27232 30529 27233
rect 30213 27168 30219 27232
rect 30283 27168 30299 27232
rect 30363 27168 30379 27232
rect 30443 27168 30459 27232
rect 30523 27168 30529 27232
rect 36302 27208 37102 27238
rect 30213 27167 30529 27168
rect 13997 27026 14063 27029
rect 15929 27026 15995 27029
rect 13997 27024 15995 27026
rect 13997 26968 14002 27024
rect 14058 26968 15934 27024
rect 15990 26968 15995 27024
rect 13997 26966 15995 26968
rect 13997 26963 14063 26966
rect 15929 26963 15995 26966
rect 7206 26688 7522 26689
rect 7206 26624 7212 26688
rect 7276 26624 7292 26688
rect 7356 26624 7372 26688
rect 7436 26624 7452 26688
rect 7516 26624 7522 26688
rect 7206 26623 7522 26624
rect 15095 26688 15411 26689
rect 15095 26624 15101 26688
rect 15165 26624 15181 26688
rect 15245 26624 15261 26688
rect 15325 26624 15341 26688
rect 15405 26624 15411 26688
rect 15095 26623 15411 26624
rect 22984 26688 23300 26689
rect 22984 26624 22990 26688
rect 23054 26624 23070 26688
rect 23134 26624 23150 26688
rect 23214 26624 23230 26688
rect 23294 26624 23300 26688
rect 22984 26623 23300 26624
rect 30873 26688 31189 26689
rect 30873 26624 30879 26688
rect 30943 26624 30959 26688
rect 31023 26624 31039 26688
rect 31103 26624 31119 26688
rect 31183 26624 31189 26688
rect 30873 26623 31189 26624
rect 17401 26348 17467 26349
rect 17350 26284 17356 26348
rect 17420 26346 17467 26348
rect 17420 26344 17512 26346
rect 17462 26288 17512 26344
rect 17420 26286 17512 26288
rect 17420 26284 17467 26286
rect 17401 26283 17467 26284
rect 6546 26144 6862 26145
rect 6546 26080 6552 26144
rect 6616 26080 6632 26144
rect 6696 26080 6712 26144
rect 6776 26080 6792 26144
rect 6856 26080 6862 26144
rect 6546 26079 6862 26080
rect 14435 26144 14751 26145
rect 14435 26080 14441 26144
rect 14505 26080 14521 26144
rect 14585 26080 14601 26144
rect 14665 26080 14681 26144
rect 14745 26080 14751 26144
rect 14435 26079 14751 26080
rect 22324 26144 22640 26145
rect 22324 26080 22330 26144
rect 22394 26080 22410 26144
rect 22474 26080 22490 26144
rect 22554 26080 22570 26144
rect 22634 26080 22640 26144
rect 22324 26079 22640 26080
rect 30213 26144 30529 26145
rect 30213 26080 30219 26144
rect 30283 26080 30299 26144
rect 30363 26080 30379 26144
rect 30443 26080 30459 26144
rect 30523 26080 30529 26144
rect 30213 26079 30529 26080
rect 0 25938 800 25968
rect 3233 25938 3299 25941
rect 0 25936 3299 25938
rect 0 25880 3238 25936
rect 3294 25880 3299 25936
rect 0 25878 3299 25880
rect 0 25848 800 25878
rect 3233 25875 3299 25878
rect 33041 25938 33107 25941
rect 36302 25938 37102 25968
rect 33041 25936 37102 25938
rect 33041 25880 33046 25936
rect 33102 25880 37102 25936
rect 33041 25878 37102 25880
rect 33041 25875 33107 25878
rect 36302 25848 37102 25878
rect 18965 25802 19031 25805
rect 26693 25802 26759 25805
rect 18965 25800 26759 25802
rect 18965 25744 18970 25800
rect 19026 25744 26698 25800
rect 26754 25744 26759 25800
rect 18965 25742 26759 25744
rect 18965 25739 19031 25742
rect 26693 25739 26759 25742
rect 7206 25600 7522 25601
rect 7206 25536 7212 25600
rect 7276 25536 7292 25600
rect 7356 25536 7372 25600
rect 7436 25536 7452 25600
rect 7516 25536 7522 25600
rect 7206 25535 7522 25536
rect 15095 25600 15411 25601
rect 15095 25536 15101 25600
rect 15165 25536 15181 25600
rect 15245 25536 15261 25600
rect 15325 25536 15341 25600
rect 15405 25536 15411 25600
rect 15095 25535 15411 25536
rect 22984 25600 23300 25601
rect 22984 25536 22990 25600
rect 23054 25536 23070 25600
rect 23134 25536 23150 25600
rect 23214 25536 23230 25600
rect 23294 25536 23300 25600
rect 22984 25535 23300 25536
rect 30873 25600 31189 25601
rect 30873 25536 30879 25600
rect 30943 25536 30959 25600
rect 31023 25536 31039 25600
rect 31103 25536 31119 25600
rect 31183 25536 31189 25600
rect 30873 25535 31189 25536
rect 6546 25056 6862 25057
rect 6546 24992 6552 25056
rect 6616 24992 6632 25056
rect 6696 24992 6712 25056
rect 6776 24992 6792 25056
rect 6856 24992 6862 25056
rect 6546 24991 6862 24992
rect 14435 25056 14751 25057
rect 14435 24992 14441 25056
rect 14505 24992 14521 25056
rect 14585 24992 14601 25056
rect 14665 24992 14681 25056
rect 14745 24992 14751 25056
rect 14435 24991 14751 24992
rect 22324 25056 22640 25057
rect 22324 24992 22330 25056
rect 22394 24992 22410 25056
rect 22474 24992 22490 25056
rect 22554 24992 22570 25056
rect 22634 24992 22640 25056
rect 22324 24991 22640 24992
rect 30213 25056 30529 25057
rect 30213 24992 30219 25056
rect 30283 24992 30299 25056
rect 30363 24992 30379 25056
rect 30443 24992 30459 25056
rect 30523 24992 30529 25056
rect 30213 24991 30529 24992
rect 5574 24924 5580 24988
rect 5644 24986 5650 24988
rect 5901 24986 5967 24989
rect 5644 24984 5967 24986
rect 5644 24928 5906 24984
rect 5962 24928 5967 24984
rect 5644 24926 5967 24928
rect 5644 24924 5650 24926
rect 5901 24923 5967 24926
rect 4337 24850 4403 24853
rect 11605 24850 11671 24853
rect 16665 24850 16731 24853
rect 4337 24848 11671 24850
rect 4337 24792 4342 24848
rect 4398 24792 11610 24848
rect 11666 24792 11671 24848
rect 4337 24790 11671 24792
rect 4337 24787 4403 24790
rect 11605 24787 11671 24790
rect 12390 24848 16731 24850
rect 12390 24792 16670 24848
rect 16726 24792 16731 24848
rect 12390 24790 16731 24792
rect 8109 24714 8175 24717
rect 12390 24714 12450 24790
rect 16665 24787 16731 24790
rect 8109 24712 12450 24714
rect 8109 24656 8114 24712
rect 8170 24656 12450 24712
rect 8109 24654 12450 24656
rect 8109 24651 8175 24654
rect 0 24578 800 24608
rect 1301 24578 1367 24581
rect 0 24576 1367 24578
rect 0 24520 1306 24576
rect 1362 24520 1367 24576
rect 0 24518 1367 24520
rect 0 24488 800 24518
rect 1301 24515 1367 24518
rect 7206 24512 7522 24513
rect 7206 24448 7212 24512
rect 7276 24448 7292 24512
rect 7356 24448 7372 24512
rect 7436 24448 7452 24512
rect 7516 24448 7522 24512
rect 7206 24447 7522 24448
rect 15095 24512 15411 24513
rect 15095 24448 15101 24512
rect 15165 24448 15181 24512
rect 15245 24448 15261 24512
rect 15325 24448 15341 24512
rect 15405 24448 15411 24512
rect 15095 24447 15411 24448
rect 22984 24512 23300 24513
rect 22984 24448 22990 24512
rect 23054 24448 23070 24512
rect 23134 24448 23150 24512
rect 23214 24448 23230 24512
rect 23294 24448 23300 24512
rect 22984 24447 23300 24448
rect 30873 24512 31189 24513
rect 30873 24448 30879 24512
rect 30943 24448 30959 24512
rect 31023 24448 31039 24512
rect 31103 24448 31119 24512
rect 31183 24448 31189 24512
rect 30873 24447 31189 24448
rect 23657 24170 23723 24173
rect 28717 24170 28783 24173
rect 23657 24168 28783 24170
rect 23657 24112 23662 24168
rect 23718 24112 28722 24168
rect 28778 24112 28783 24168
rect 23657 24110 28783 24112
rect 23657 24107 23723 24110
rect 28717 24107 28783 24110
rect 26601 24036 26667 24037
rect 26550 23972 26556 24036
rect 26620 24034 26667 24036
rect 26620 24032 26712 24034
rect 26662 23976 26712 24032
rect 26620 23974 26712 23976
rect 26620 23972 26667 23974
rect 26601 23971 26667 23972
rect 6546 23968 6862 23969
rect 6546 23904 6552 23968
rect 6616 23904 6632 23968
rect 6696 23904 6712 23968
rect 6776 23904 6792 23968
rect 6856 23904 6862 23968
rect 6546 23903 6862 23904
rect 14435 23968 14751 23969
rect 14435 23904 14441 23968
rect 14505 23904 14521 23968
rect 14585 23904 14601 23968
rect 14665 23904 14681 23968
rect 14745 23904 14751 23968
rect 14435 23903 14751 23904
rect 22324 23968 22640 23969
rect 22324 23904 22330 23968
rect 22394 23904 22410 23968
rect 22474 23904 22490 23968
rect 22554 23904 22570 23968
rect 22634 23904 22640 23968
rect 22324 23903 22640 23904
rect 30213 23968 30529 23969
rect 30213 23904 30219 23968
rect 30283 23904 30299 23968
rect 30363 23904 30379 23968
rect 30443 23904 30459 23968
rect 30523 23904 30529 23968
rect 30213 23903 30529 23904
rect 34697 23898 34763 23901
rect 36302 23898 37102 23928
rect 34697 23896 37102 23898
rect 34697 23840 34702 23896
rect 34758 23840 37102 23896
rect 34697 23838 37102 23840
rect 34697 23835 34763 23838
rect 36302 23808 37102 23838
rect 15561 23762 15627 23765
rect 15694 23762 15700 23764
rect 15561 23760 15700 23762
rect 15561 23704 15566 23760
rect 15622 23704 15700 23760
rect 15561 23702 15700 23704
rect 15561 23699 15627 23702
rect 15694 23700 15700 23702
rect 15764 23700 15770 23764
rect 6177 23628 6243 23629
rect 6126 23564 6132 23628
rect 6196 23626 6243 23628
rect 10041 23626 10107 23629
rect 12617 23626 12683 23629
rect 6196 23624 6288 23626
rect 6238 23568 6288 23624
rect 6196 23566 6288 23568
rect 10041 23624 12683 23626
rect 10041 23568 10046 23624
rect 10102 23568 12622 23624
rect 12678 23568 12683 23624
rect 10041 23566 12683 23568
rect 6196 23564 6243 23566
rect 6177 23563 6243 23564
rect 10041 23563 10107 23566
rect 12617 23563 12683 23566
rect 5809 23492 5875 23493
rect 5758 23428 5764 23492
rect 5828 23490 5875 23492
rect 5828 23488 5920 23490
rect 5870 23432 5920 23488
rect 5828 23430 5920 23432
rect 5828 23428 5875 23430
rect 5809 23427 5875 23428
rect 7206 23424 7522 23425
rect 7206 23360 7212 23424
rect 7276 23360 7292 23424
rect 7356 23360 7372 23424
rect 7436 23360 7452 23424
rect 7516 23360 7522 23424
rect 7206 23359 7522 23360
rect 15095 23424 15411 23425
rect 15095 23360 15101 23424
rect 15165 23360 15181 23424
rect 15245 23360 15261 23424
rect 15325 23360 15341 23424
rect 15405 23360 15411 23424
rect 15095 23359 15411 23360
rect 22984 23424 23300 23425
rect 22984 23360 22990 23424
rect 23054 23360 23070 23424
rect 23134 23360 23150 23424
rect 23214 23360 23230 23424
rect 23294 23360 23300 23424
rect 22984 23359 23300 23360
rect 30873 23424 31189 23425
rect 30873 23360 30879 23424
rect 30943 23360 30959 23424
rect 31023 23360 31039 23424
rect 31103 23360 31119 23424
rect 31183 23360 31189 23424
rect 30873 23359 31189 23360
rect 0 23218 800 23248
rect 3509 23218 3575 23221
rect 0 23216 3575 23218
rect 0 23160 3514 23216
rect 3570 23160 3575 23216
rect 0 23158 3575 23160
rect 0 23128 800 23158
rect 3509 23155 3575 23158
rect 11605 23218 11671 23221
rect 16481 23218 16547 23221
rect 11605 23216 16547 23218
rect 11605 23160 11610 23216
rect 11666 23160 16486 23216
rect 16542 23160 16547 23216
rect 11605 23158 16547 23160
rect 11605 23155 11671 23158
rect 16481 23155 16547 23158
rect 6546 22880 6862 22881
rect 6546 22816 6552 22880
rect 6616 22816 6632 22880
rect 6696 22816 6712 22880
rect 6776 22816 6792 22880
rect 6856 22816 6862 22880
rect 6546 22815 6862 22816
rect 14435 22880 14751 22881
rect 14435 22816 14441 22880
rect 14505 22816 14521 22880
rect 14585 22816 14601 22880
rect 14665 22816 14681 22880
rect 14745 22816 14751 22880
rect 14435 22815 14751 22816
rect 22324 22880 22640 22881
rect 22324 22816 22330 22880
rect 22394 22816 22410 22880
rect 22474 22816 22490 22880
rect 22554 22816 22570 22880
rect 22634 22816 22640 22880
rect 22324 22815 22640 22816
rect 30213 22880 30529 22881
rect 30213 22816 30219 22880
rect 30283 22816 30299 22880
rect 30363 22816 30379 22880
rect 30443 22816 30459 22880
rect 30523 22816 30529 22880
rect 30213 22815 30529 22816
rect 35157 22538 35223 22541
rect 36302 22538 37102 22568
rect 35157 22536 37102 22538
rect 35157 22480 35162 22536
rect 35218 22480 37102 22536
rect 35157 22478 37102 22480
rect 35157 22475 35223 22478
rect 36302 22448 37102 22478
rect 7206 22336 7522 22337
rect 7206 22272 7212 22336
rect 7276 22272 7292 22336
rect 7356 22272 7372 22336
rect 7436 22272 7452 22336
rect 7516 22272 7522 22336
rect 7206 22271 7522 22272
rect 15095 22336 15411 22337
rect 15095 22272 15101 22336
rect 15165 22272 15181 22336
rect 15245 22272 15261 22336
rect 15325 22272 15341 22336
rect 15405 22272 15411 22336
rect 15095 22271 15411 22272
rect 22984 22336 23300 22337
rect 22984 22272 22990 22336
rect 23054 22272 23070 22336
rect 23134 22272 23150 22336
rect 23214 22272 23230 22336
rect 23294 22272 23300 22336
rect 22984 22271 23300 22272
rect 30873 22336 31189 22337
rect 30873 22272 30879 22336
rect 30943 22272 30959 22336
rect 31023 22272 31039 22336
rect 31103 22272 31119 22336
rect 31183 22272 31189 22336
rect 30873 22271 31189 22272
rect 23197 22130 23263 22133
rect 26049 22130 26115 22133
rect 23197 22128 26115 22130
rect 23197 22072 23202 22128
rect 23258 22072 26054 22128
rect 26110 22072 26115 22128
rect 23197 22070 26115 22072
rect 23197 22067 23263 22070
rect 26049 22067 26115 22070
rect 27613 22130 27679 22133
rect 27981 22130 28047 22133
rect 27613 22128 28047 22130
rect 27613 22072 27618 22128
rect 27674 22072 27986 22128
rect 28042 22072 28047 22128
rect 27613 22070 28047 22072
rect 27613 22067 27679 22070
rect 27981 22067 28047 22070
rect 6546 21792 6862 21793
rect 6546 21728 6552 21792
rect 6616 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6862 21792
rect 6546 21727 6862 21728
rect 14435 21792 14751 21793
rect 14435 21728 14441 21792
rect 14505 21728 14521 21792
rect 14585 21728 14601 21792
rect 14665 21728 14681 21792
rect 14745 21728 14751 21792
rect 14435 21727 14751 21728
rect 22324 21792 22640 21793
rect 22324 21728 22330 21792
rect 22394 21728 22410 21792
rect 22474 21728 22490 21792
rect 22554 21728 22570 21792
rect 22634 21728 22640 21792
rect 22324 21727 22640 21728
rect 30213 21792 30529 21793
rect 30213 21728 30219 21792
rect 30283 21728 30299 21792
rect 30363 21728 30379 21792
rect 30443 21728 30459 21792
rect 30523 21728 30529 21792
rect 30213 21727 30529 21728
rect 11697 21722 11763 21725
rect 11830 21722 11836 21724
rect 11697 21720 11836 21722
rect 11697 21664 11702 21720
rect 11758 21664 11836 21720
rect 11697 21662 11836 21664
rect 11697 21659 11763 21662
rect 11830 21660 11836 21662
rect 11900 21660 11906 21724
rect 9857 21586 9923 21589
rect 17125 21586 17191 21589
rect 9857 21584 17191 21586
rect 9857 21528 9862 21584
rect 9918 21528 17130 21584
rect 17186 21528 17191 21584
rect 9857 21526 17191 21528
rect 9857 21523 9923 21526
rect 17125 21523 17191 21526
rect 7206 21248 7522 21249
rect 0 21178 800 21208
rect 7206 21184 7212 21248
rect 7276 21184 7292 21248
rect 7356 21184 7372 21248
rect 7436 21184 7452 21248
rect 7516 21184 7522 21248
rect 7206 21183 7522 21184
rect 15095 21248 15411 21249
rect 15095 21184 15101 21248
rect 15165 21184 15181 21248
rect 15245 21184 15261 21248
rect 15325 21184 15341 21248
rect 15405 21184 15411 21248
rect 15095 21183 15411 21184
rect 22984 21248 23300 21249
rect 22984 21184 22990 21248
rect 23054 21184 23070 21248
rect 23134 21184 23150 21248
rect 23214 21184 23230 21248
rect 23294 21184 23300 21248
rect 22984 21183 23300 21184
rect 30873 21248 31189 21249
rect 30873 21184 30879 21248
rect 30943 21184 30959 21248
rect 31023 21184 31039 21248
rect 31103 21184 31119 21248
rect 31183 21184 31189 21248
rect 30873 21183 31189 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 34881 21178 34947 21181
rect 36302 21178 37102 21208
rect 34881 21176 37102 21178
rect 34881 21120 34886 21176
rect 34942 21120 37102 21176
rect 34881 21118 37102 21120
rect 34881 21115 34947 21118
rect 36302 21088 37102 21118
rect 5533 21042 5599 21045
rect 12709 21042 12775 21045
rect 5533 21040 12775 21042
rect 5533 20984 5538 21040
rect 5594 20984 12714 21040
rect 12770 20984 12775 21040
rect 5533 20982 12775 20984
rect 5533 20979 5599 20982
rect 12709 20979 12775 20982
rect 10041 20906 10107 20909
rect 11513 20906 11579 20909
rect 10041 20904 11579 20906
rect 10041 20848 10046 20904
rect 10102 20848 11518 20904
rect 11574 20848 11579 20904
rect 10041 20846 11579 20848
rect 10041 20843 10107 20846
rect 11513 20843 11579 20846
rect 19374 20708 19380 20772
rect 19444 20770 19450 20772
rect 19701 20770 19767 20773
rect 19444 20768 19767 20770
rect 19444 20712 19706 20768
rect 19762 20712 19767 20768
rect 19444 20710 19767 20712
rect 19444 20708 19450 20710
rect 19701 20707 19767 20710
rect 6546 20704 6862 20705
rect 6546 20640 6552 20704
rect 6616 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6862 20704
rect 6546 20639 6862 20640
rect 14435 20704 14751 20705
rect 14435 20640 14441 20704
rect 14505 20640 14521 20704
rect 14585 20640 14601 20704
rect 14665 20640 14681 20704
rect 14745 20640 14751 20704
rect 14435 20639 14751 20640
rect 22324 20704 22640 20705
rect 22324 20640 22330 20704
rect 22394 20640 22410 20704
rect 22474 20640 22490 20704
rect 22554 20640 22570 20704
rect 22634 20640 22640 20704
rect 22324 20639 22640 20640
rect 30213 20704 30529 20705
rect 30213 20640 30219 20704
rect 30283 20640 30299 20704
rect 30363 20640 30379 20704
rect 30443 20640 30459 20704
rect 30523 20640 30529 20704
rect 30213 20639 30529 20640
rect 11881 20500 11947 20501
rect 11830 20436 11836 20500
rect 11900 20498 11947 20500
rect 11900 20496 11992 20498
rect 11942 20440 11992 20496
rect 11900 20438 11992 20440
rect 11900 20436 11947 20438
rect 12198 20436 12204 20500
rect 12268 20498 12274 20500
rect 17125 20498 17191 20501
rect 12268 20496 17191 20498
rect 12268 20440 17130 20496
rect 17186 20440 17191 20496
rect 12268 20438 17191 20440
rect 12268 20436 12274 20438
rect 11881 20435 11947 20436
rect 17125 20435 17191 20438
rect 10501 20362 10567 20365
rect 19057 20362 19123 20365
rect 10501 20360 19123 20362
rect 10501 20304 10506 20360
rect 10562 20304 19062 20360
rect 19118 20304 19123 20360
rect 10501 20302 19123 20304
rect 10501 20299 10567 20302
rect 19057 20299 19123 20302
rect 20529 20362 20595 20365
rect 21909 20362 21975 20365
rect 20529 20360 21975 20362
rect 20529 20304 20534 20360
rect 20590 20304 21914 20360
rect 21970 20304 21975 20360
rect 20529 20302 21975 20304
rect 20529 20299 20595 20302
rect 21909 20299 21975 20302
rect 5809 20226 5875 20229
rect 6126 20226 6132 20228
rect 5809 20224 6132 20226
rect 5809 20168 5814 20224
rect 5870 20168 6132 20224
rect 5809 20166 6132 20168
rect 5809 20163 5875 20166
rect 6126 20164 6132 20166
rect 6196 20164 6202 20228
rect 7206 20160 7522 20161
rect 7206 20096 7212 20160
rect 7276 20096 7292 20160
rect 7356 20096 7372 20160
rect 7436 20096 7452 20160
rect 7516 20096 7522 20160
rect 7206 20095 7522 20096
rect 15095 20160 15411 20161
rect 15095 20096 15101 20160
rect 15165 20096 15181 20160
rect 15245 20096 15261 20160
rect 15325 20096 15341 20160
rect 15405 20096 15411 20160
rect 15095 20095 15411 20096
rect 22984 20160 23300 20161
rect 22984 20096 22990 20160
rect 23054 20096 23070 20160
rect 23134 20096 23150 20160
rect 23214 20096 23230 20160
rect 23294 20096 23300 20160
rect 22984 20095 23300 20096
rect 30873 20160 31189 20161
rect 30873 20096 30879 20160
rect 30943 20096 30959 20160
rect 31023 20096 31039 20160
rect 31103 20096 31119 20160
rect 31183 20096 31189 20160
rect 30873 20095 31189 20096
rect 10869 20090 10935 20093
rect 13813 20090 13879 20093
rect 10869 20088 13879 20090
rect 10869 20032 10874 20088
rect 10930 20032 13818 20088
rect 13874 20032 13879 20088
rect 10869 20030 13879 20032
rect 10869 20027 10935 20030
rect 13813 20027 13879 20030
rect 11053 19954 11119 19957
rect 14181 19954 14247 19957
rect 11053 19952 14247 19954
rect 11053 19896 11058 19952
rect 11114 19896 14186 19952
rect 14242 19896 14247 19952
rect 11053 19894 14247 19896
rect 11053 19891 11119 19894
rect 14181 19891 14247 19894
rect 29821 19954 29887 19957
rect 32397 19954 32463 19957
rect 29821 19952 32463 19954
rect 29821 19896 29826 19952
rect 29882 19896 32402 19952
rect 32458 19896 32463 19952
rect 29821 19894 32463 19896
rect 29821 19891 29887 19894
rect 32397 19891 32463 19894
rect 0 19818 800 19848
rect 3233 19818 3299 19821
rect 0 19816 3299 19818
rect 0 19760 3238 19816
rect 3294 19760 3299 19816
rect 0 19758 3299 19760
rect 0 19728 800 19758
rect 3233 19755 3299 19758
rect 9029 19818 9095 19821
rect 11329 19818 11395 19821
rect 9029 19816 11395 19818
rect 9029 19760 9034 19816
rect 9090 19760 11334 19816
rect 11390 19760 11395 19816
rect 9029 19758 11395 19760
rect 9029 19755 9095 19758
rect 11329 19755 11395 19758
rect 33777 19818 33843 19821
rect 36302 19818 37102 19848
rect 33777 19816 37102 19818
rect 33777 19760 33782 19816
rect 33838 19760 37102 19816
rect 33777 19758 37102 19760
rect 33777 19755 33843 19758
rect 36302 19728 37102 19758
rect 6546 19616 6862 19617
rect 6546 19552 6552 19616
rect 6616 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6862 19616
rect 6546 19551 6862 19552
rect 14435 19616 14751 19617
rect 14435 19552 14441 19616
rect 14505 19552 14521 19616
rect 14585 19552 14601 19616
rect 14665 19552 14681 19616
rect 14745 19552 14751 19616
rect 14435 19551 14751 19552
rect 22324 19616 22640 19617
rect 22324 19552 22330 19616
rect 22394 19552 22410 19616
rect 22474 19552 22490 19616
rect 22554 19552 22570 19616
rect 22634 19552 22640 19616
rect 22324 19551 22640 19552
rect 30213 19616 30529 19617
rect 30213 19552 30219 19616
rect 30283 19552 30299 19616
rect 30363 19552 30379 19616
rect 30443 19552 30459 19616
rect 30523 19552 30529 19616
rect 30213 19551 30529 19552
rect 10685 19546 10751 19549
rect 11237 19546 11303 19549
rect 10685 19544 11303 19546
rect 10685 19488 10690 19544
rect 10746 19488 11242 19544
rect 11298 19488 11303 19544
rect 10685 19486 11303 19488
rect 10685 19483 10751 19486
rect 11237 19483 11303 19486
rect 5165 19410 5231 19413
rect 6361 19410 6427 19413
rect 5165 19408 6427 19410
rect 5165 19352 5170 19408
rect 5226 19352 6366 19408
rect 6422 19352 6427 19408
rect 5165 19350 6427 19352
rect 5165 19347 5231 19350
rect 6361 19347 6427 19350
rect 20069 19410 20135 19413
rect 27981 19410 28047 19413
rect 20069 19408 28047 19410
rect 20069 19352 20074 19408
rect 20130 19352 27986 19408
rect 28042 19352 28047 19408
rect 20069 19350 28047 19352
rect 29177 19350 29243 19353
rect 20069 19347 20135 19350
rect 27981 19347 28047 19350
rect 28996 19348 29243 19350
rect 28996 19292 29182 19348
rect 29238 19292 29243 19348
rect 28996 19290 29243 19292
rect 6729 19274 6795 19277
rect 12801 19274 12867 19277
rect 14365 19274 14431 19277
rect 6729 19272 9690 19274
rect 6729 19216 6734 19272
rect 6790 19216 9690 19272
rect 6729 19214 9690 19216
rect 6729 19211 6795 19214
rect 7206 19072 7522 19073
rect 7206 19008 7212 19072
rect 7276 19008 7292 19072
rect 7356 19008 7372 19072
rect 7436 19008 7452 19072
rect 7516 19008 7522 19072
rect 7206 19007 7522 19008
rect 9630 19002 9690 19214
rect 12801 19272 14431 19274
rect 12801 19216 12806 19272
rect 12862 19216 14370 19272
rect 14426 19216 14431 19272
rect 12801 19214 14431 19216
rect 12801 19211 12867 19214
rect 14365 19211 14431 19214
rect 15095 19072 15411 19073
rect 15095 19008 15101 19072
rect 15165 19008 15181 19072
rect 15245 19008 15261 19072
rect 15325 19008 15341 19072
rect 15405 19008 15411 19072
rect 15095 19007 15411 19008
rect 22984 19072 23300 19073
rect 22984 19008 22990 19072
rect 23054 19008 23070 19072
rect 23134 19008 23150 19072
rect 23214 19008 23230 19072
rect 23294 19008 23300 19072
rect 22984 19007 23300 19008
rect 9949 19002 10015 19005
rect 9630 19000 10015 19002
rect 9630 18944 9954 19000
rect 10010 18944 10015 19000
rect 9630 18942 10015 18944
rect 28996 19002 29056 19290
rect 29177 19287 29243 19290
rect 29177 19138 29243 19141
rect 29821 19138 29887 19141
rect 29177 19136 29887 19138
rect 29177 19080 29182 19136
rect 29238 19080 29826 19136
rect 29882 19080 29887 19136
rect 29177 19078 29887 19080
rect 29177 19075 29243 19078
rect 29821 19075 29887 19078
rect 30873 19072 31189 19073
rect 30873 19008 30879 19072
rect 30943 19008 30959 19072
rect 31023 19008 31039 19072
rect 31103 19008 31119 19072
rect 31183 19008 31189 19072
rect 30873 19007 31189 19008
rect 29361 19002 29427 19005
rect 28996 19000 29427 19002
rect 28996 18944 29366 19000
rect 29422 18944 29427 19000
rect 28996 18942 29427 18944
rect 9949 18939 10015 18942
rect 29361 18939 29427 18942
rect 19517 18866 19583 18869
rect 20345 18866 20411 18869
rect 19517 18864 20411 18866
rect 19517 18808 19522 18864
rect 19578 18808 20350 18864
rect 20406 18808 20411 18864
rect 19517 18806 20411 18808
rect 19517 18803 19583 18806
rect 20345 18803 20411 18806
rect 6546 18528 6862 18529
rect 0 18458 800 18488
rect 6546 18464 6552 18528
rect 6616 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6862 18528
rect 6546 18463 6862 18464
rect 14435 18528 14751 18529
rect 14435 18464 14441 18528
rect 14505 18464 14521 18528
rect 14585 18464 14601 18528
rect 14665 18464 14681 18528
rect 14745 18464 14751 18528
rect 14435 18463 14751 18464
rect 22324 18528 22640 18529
rect 22324 18464 22330 18528
rect 22394 18464 22410 18528
rect 22474 18464 22490 18528
rect 22554 18464 22570 18528
rect 22634 18464 22640 18528
rect 22324 18463 22640 18464
rect 30213 18528 30529 18529
rect 30213 18464 30219 18528
rect 30283 18464 30299 18528
rect 30363 18464 30379 18528
rect 30443 18464 30459 18528
rect 30523 18464 30529 18528
rect 30213 18463 30529 18464
rect 1301 18458 1367 18461
rect 0 18456 1367 18458
rect 0 18400 1306 18456
rect 1362 18400 1367 18456
rect 0 18398 1367 18400
rect 0 18368 800 18398
rect 1301 18395 1367 18398
rect 34513 18458 34579 18461
rect 36302 18458 37102 18488
rect 34513 18456 37102 18458
rect 34513 18400 34518 18456
rect 34574 18400 37102 18456
rect 34513 18398 37102 18400
rect 34513 18395 34579 18398
rect 36302 18368 37102 18398
rect 5717 18322 5783 18325
rect 8661 18322 8727 18325
rect 5717 18320 8727 18322
rect 5717 18264 5722 18320
rect 5778 18264 8666 18320
rect 8722 18264 8727 18320
rect 5717 18262 8727 18264
rect 5717 18259 5783 18262
rect 8661 18259 8727 18262
rect 14917 18322 14983 18325
rect 18781 18322 18847 18325
rect 14917 18320 18847 18322
rect 14917 18264 14922 18320
rect 14978 18264 18786 18320
rect 18842 18264 18847 18320
rect 14917 18262 18847 18264
rect 14917 18259 14983 18262
rect 18781 18259 18847 18262
rect 14273 18186 14339 18189
rect 14273 18184 15578 18186
rect 14273 18128 14278 18184
rect 14334 18128 15578 18184
rect 14273 18126 15578 18128
rect 14273 18123 14339 18126
rect 7206 17984 7522 17985
rect 7206 17920 7212 17984
rect 7276 17920 7292 17984
rect 7356 17920 7372 17984
rect 7436 17920 7452 17984
rect 7516 17920 7522 17984
rect 7206 17919 7522 17920
rect 15095 17984 15411 17985
rect 15095 17920 15101 17984
rect 15165 17920 15181 17984
rect 15245 17920 15261 17984
rect 15325 17920 15341 17984
rect 15405 17920 15411 17984
rect 15095 17919 15411 17920
rect 15518 17914 15578 18126
rect 19517 18052 19583 18053
rect 19517 18048 19564 18052
rect 19628 18050 19634 18052
rect 19517 17992 19522 18048
rect 19517 17988 19564 17992
rect 19628 17990 19674 18050
rect 19628 17988 19634 17990
rect 19517 17987 19583 17988
rect 22984 17984 23300 17985
rect 22984 17920 22990 17984
rect 23054 17920 23070 17984
rect 23134 17920 23150 17984
rect 23214 17920 23230 17984
rect 23294 17920 23300 17984
rect 22984 17919 23300 17920
rect 30873 17984 31189 17985
rect 30873 17920 30879 17984
rect 30943 17920 30959 17984
rect 31023 17920 31039 17984
rect 31103 17920 31119 17984
rect 31183 17920 31189 17984
rect 30873 17919 31189 17920
rect 16021 17914 16087 17917
rect 19701 17916 19767 17917
rect 19701 17914 19748 17916
rect 15518 17912 19748 17914
rect 19812 17914 19818 17916
rect 28073 17914 28139 17917
rect 28717 17914 28783 17917
rect 15518 17856 16026 17912
rect 16082 17856 19706 17912
rect 15518 17854 19748 17856
rect 16021 17851 16087 17854
rect 19701 17852 19748 17854
rect 19812 17854 19894 17914
rect 28073 17912 28783 17914
rect 28073 17856 28078 17912
rect 28134 17856 28722 17912
rect 28778 17856 28783 17912
rect 28073 17854 28783 17856
rect 19812 17852 19818 17854
rect 19701 17851 19767 17852
rect 28073 17851 28139 17854
rect 28717 17851 28783 17854
rect 7741 17778 7807 17781
rect 19517 17778 19583 17781
rect 7741 17776 19583 17778
rect 7741 17720 7746 17776
rect 7802 17720 19522 17776
rect 19578 17720 19583 17776
rect 7741 17718 19583 17720
rect 7741 17715 7807 17718
rect 19517 17715 19583 17718
rect 22134 17716 22140 17780
rect 22204 17778 22210 17780
rect 22645 17778 22711 17781
rect 22204 17776 22711 17778
rect 22204 17720 22650 17776
rect 22706 17720 22711 17776
rect 22204 17718 22711 17720
rect 22204 17716 22210 17718
rect 22645 17715 22711 17718
rect 28257 17778 28323 17781
rect 28809 17778 28875 17781
rect 28257 17776 28875 17778
rect 28257 17720 28262 17776
rect 28318 17720 28814 17776
rect 28870 17720 28875 17776
rect 28257 17718 28875 17720
rect 28257 17715 28323 17718
rect 28809 17715 28875 17718
rect 13629 17642 13695 17645
rect 18137 17642 18203 17645
rect 13629 17640 18203 17642
rect 13629 17584 13634 17640
rect 13690 17584 18142 17640
rect 18198 17584 18203 17640
rect 13629 17582 18203 17584
rect 13629 17579 13695 17582
rect 18137 17579 18203 17582
rect 6546 17440 6862 17441
rect 6546 17376 6552 17440
rect 6616 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6862 17440
rect 6546 17375 6862 17376
rect 14435 17440 14751 17441
rect 14435 17376 14441 17440
rect 14505 17376 14521 17440
rect 14585 17376 14601 17440
rect 14665 17376 14681 17440
rect 14745 17376 14751 17440
rect 14435 17375 14751 17376
rect 22324 17440 22640 17441
rect 22324 17376 22330 17440
rect 22394 17376 22410 17440
rect 22474 17376 22490 17440
rect 22554 17376 22570 17440
rect 22634 17376 22640 17440
rect 22324 17375 22640 17376
rect 30213 17440 30529 17441
rect 30213 17376 30219 17440
rect 30283 17376 30299 17440
rect 30363 17376 30379 17440
rect 30443 17376 30459 17440
rect 30523 17376 30529 17440
rect 30213 17375 30529 17376
rect 20529 17234 20595 17237
rect 26969 17234 27035 17237
rect 20529 17232 27035 17234
rect 20529 17176 20534 17232
rect 20590 17176 26974 17232
rect 27030 17176 27035 17232
rect 20529 17174 27035 17176
rect 20529 17171 20595 17174
rect 26969 17171 27035 17174
rect 0 17098 800 17128
rect 1301 17098 1367 17101
rect 0 17096 1367 17098
rect 0 17040 1306 17096
rect 1362 17040 1367 17096
rect 0 17038 1367 17040
rect 0 17008 800 17038
rect 1301 17035 1367 17038
rect 12801 17098 12867 17101
rect 18137 17098 18203 17101
rect 12801 17096 18203 17098
rect 12801 17040 12806 17096
rect 12862 17040 18142 17096
rect 18198 17040 18203 17096
rect 12801 17038 18203 17040
rect 12801 17035 12867 17038
rect 18137 17035 18203 17038
rect 33041 17098 33107 17101
rect 36302 17098 37102 17128
rect 33041 17096 37102 17098
rect 33041 17040 33046 17096
rect 33102 17040 37102 17096
rect 33041 17038 37102 17040
rect 33041 17035 33107 17038
rect 36302 17008 37102 17038
rect 7206 16896 7522 16897
rect 7206 16832 7212 16896
rect 7276 16832 7292 16896
rect 7356 16832 7372 16896
rect 7436 16832 7452 16896
rect 7516 16832 7522 16896
rect 7206 16831 7522 16832
rect 15095 16896 15411 16897
rect 15095 16832 15101 16896
rect 15165 16832 15181 16896
rect 15245 16832 15261 16896
rect 15325 16832 15341 16896
rect 15405 16832 15411 16896
rect 15095 16831 15411 16832
rect 22984 16896 23300 16897
rect 22984 16832 22990 16896
rect 23054 16832 23070 16896
rect 23134 16832 23150 16896
rect 23214 16832 23230 16896
rect 23294 16832 23300 16896
rect 22984 16831 23300 16832
rect 30873 16896 31189 16897
rect 30873 16832 30879 16896
rect 30943 16832 30959 16896
rect 31023 16832 31039 16896
rect 31103 16832 31119 16896
rect 31183 16832 31189 16896
rect 30873 16831 31189 16832
rect 6546 16352 6862 16353
rect 6546 16288 6552 16352
rect 6616 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6862 16352
rect 6546 16287 6862 16288
rect 14435 16352 14751 16353
rect 14435 16288 14441 16352
rect 14505 16288 14521 16352
rect 14585 16288 14601 16352
rect 14665 16288 14681 16352
rect 14745 16288 14751 16352
rect 14435 16287 14751 16288
rect 22324 16352 22640 16353
rect 22324 16288 22330 16352
rect 22394 16288 22410 16352
rect 22474 16288 22490 16352
rect 22554 16288 22570 16352
rect 22634 16288 22640 16352
rect 22324 16287 22640 16288
rect 30213 16352 30529 16353
rect 30213 16288 30219 16352
rect 30283 16288 30299 16352
rect 30363 16288 30379 16352
rect 30443 16288 30459 16352
rect 30523 16288 30529 16352
rect 30213 16287 30529 16288
rect 20161 16010 20227 16013
rect 20161 16008 20914 16010
rect 20161 15952 20166 16008
rect 20222 15952 20914 16008
rect 20161 15950 20914 15952
rect 20161 15947 20227 15950
rect 20854 15877 20914 15950
rect 20854 15872 20963 15877
rect 20854 15816 20902 15872
rect 20958 15816 20963 15872
rect 20854 15814 20963 15816
rect 20897 15811 20963 15814
rect 7206 15808 7522 15809
rect 0 15738 800 15768
rect 7206 15744 7212 15808
rect 7276 15744 7292 15808
rect 7356 15744 7372 15808
rect 7436 15744 7452 15808
rect 7516 15744 7522 15808
rect 7206 15743 7522 15744
rect 15095 15808 15411 15809
rect 15095 15744 15101 15808
rect 15165 15744 15181 15808
rect 15245 15744 15261 15808
rect 15325 15744 15341 15808
rect 15405 15744 15411 15808
rect 15095 15743 15411 15744
rect 22984 15808 23300 15809
rect 22984 15744 22990 15808
rect 23054 15744 23070 15808
rect 23134 15744 23150 15808
rect 23214 15744 23230 15808
rect 23294 15744 23300 15808
rect 22984 15743 23300 15744
rect 30873 15808 31189 15809
rect 30873 15744 30879 15808
rect 30943 15744 30959 15808
rect 31023 15744 31039 15808
rect 31103 15744 31119 15808
rect 31183 15744 31189 15808
rect 30873 15743 31189 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 34881 15738 34947 15741
rect 36302 15738 37102 15768
rect 34881 15736 37102 15738
rect 34881 15680 34886 15736
rect 34942 15680 37102 15736
rect 34881 15678 37102 15680
rect 34881 15675 34947 15678
rect 36302 15648 37102 15678
rect 18822 15268 18828 15332
rect 18892 15330 18898 15332
rect 19241 15330 19307 15333
rect 18892 15328 19307 15330
rect 18892 15272 19246 15328
rect 19302 15272 19307 15328
rect 18892 15270 19307 15272
rect 18892 15268 18898 15270
rect 19241 15267 19307 15270
rect 6546 15264 6862 15265
rect 6546 15200 6552 15264
rect 6616 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6862 15264
rect 6546 15199 6862 15200
rect 14435 15264 14751 15265
rect 14435 15200 14441 15264
rect 14505 15200 14521 15264
rect 14585 15200 14601 15264
rect 14665 15200 14681 15264
rect 14745 15200 14751 15264
rect 14435 15199 14751 15200
rect 22324 15264 22640 15265
rect 22324 15200 22330 15264
rect 22394 15200 22410 15264
rect 22474 15200 22490 15264
rect 22554 15200 22570 15264
rect 22634 15200 22640 15264
rect 22324 15199 22640 15200
rect 30213 15264 30529 15265
rect 30213 15200 30219 15264
rect 30283 15200 30299 15264
rect 30363 15200 30379 15264
rect 30443 15200 30459 15264
rect 30523 15200 30529 15264
rect 30213 15199 30529 15200
rect 5574 15132 5580 15196
rect 5644 15194 5650 15196
rect 5717 15194 5783 15197
rect 5644 15192 5783 15194
rect 5644 15136 5722 15192
rect 5778 15136 5783 15192
rect 5644 15134 5783 15136
rect 5644 15132 5650 15134
rect 5717 15131 5783 15134
rect 19742 15132 19748 15196
rect 19812 15194 19818 15196
rect 20069 15194 20135 15197
rect 19812 15192 20135 15194
rect 19812 15136 20074 15192
rect 20130 15136 20135 15192
rect 19812 15134 20135 15136
rect 19812 15132 19818 15134
rect 20069 15131 20135 15134
rect 21817 14786 21883 14789
rect 22185 14786 22251 14789
rect 21817 14784 22251 14786
rect 21817 14728 21822 14784
rect 21878 14728 22190 14784
rect 22246 14728 22251 14784
rect 21817 14726 22251 14728
rect 21817 14723 21883 14726
rect 22185 14723 22251 14726
rect 7206 14720 7522 14721
rect 7206 14656 7212 14720
rect 7276 14656 7292 14720
rect 7356 14656 7372 14720
rect 7436 14656 7452 14720
rect 7516 14656 7522 14720
rect 7206 14655 7522 14656
rect 15095 14720 15411 14721
rect 15095 14656 15101 14720
rect 15165 14656 15181 14720
rect 15245 14656 15261 14720
rect 15325 14656 15341 14720
rect 15405 14656 15411 14720
rect 15095 14655 15411 14656
rect 22984 14720 23300 14721
rect 22984 14656 22990 14720
rect 23054 14656 23070 14720
rect 23134 14656 23150 14720
rect 23214 14656 23230 14720
rect 23294 14656 23300 14720
rect 22984 14655 23300 14656
rect 30873 14720 31189 14721
rect 30873 14656 30879 14720
rect 30943 14656 30959 14720
rect 31023 14656 31039 14720
rect 31103 14656 31119 14720
rect 31183 14656 31189 14720
rect 30873 14655 31189 14656
rect 23933 14514 23999 14517
rect 28993 14514 29059 14517
rect 23933 14512 29059 14514
rect 23933 14456 23938 14512
rect 23994 14456 28998 14512
rect 29054 14456 29059 14512
rect 23933 14454 29059 14456
rect 23933 14451 23999 14454
rect 28993 14451 29059 14454
rect 0 14378 800 14408
rect 1301 14378 1367 14381
rect 0 14376 1367 14378
rect 0 14320 1306 14376
rect 1362 14320 1367 14376
rect 0 14318 1367 14320
rect 0 14288 800 14318
rect 1301 14315 1367 14318
rect 6546 14176 6862 14177
rect 6546 14112 6552 14176
rect 6616 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6862 14176
rect 6546 14111 6862 14112
rect 14435 14176 14751 14177
rect 14435 14112 14441 14176
rect 14505 14112 14521 14176
rect 14585 14112 14601 14176
rect 14665 14112 14681 14176
rect 14745 14112 14751 14176
rect 14435 14111 14751 14112
rect 22324 14176 22640 14177
rect 22324 14112 22330 14176
rect 22394 14112 22410 14176
rect 22474 14112 22490 14176
rect 22554 14112 22570 14176
rect 22634 14112 22640 14176
rect 22324 14111 22640 14112
rect 30213 14176 30529 14177
rect 30213 14112 30219 14176
rect 30283 14112 30299 14176
rect 30363 14112 30379 14176
rect 30443 14112 30459 14176
rect 30523 14112 30529 14176
rect 30213 14111 30529 14112
rect 15469 14106 15535 14109
rect 17677 14106 17743 14109
rect 15469 14104 17743 14106
rect 15469 14048 15474 14104
rect 15530 14048 17682 14104
rect 17738 14048 17743 14104
rect 15469 14046 17743 14048
rect 15469 14043 15535 14046
rect 17677 14043 17743 14046
rect 10910 13908 10916 13972
rect 10980 13970 10986 13972
rect 23381 13970 23447 13973
rect 10980 13968 23447 13970
rect 10980 13912 23386 13968
rect 23442 13912 23447 13968
rect 10980 13910 23447 13912
rect 10980 13908 10986 13910
rect 23381 13907 23447 13910
rect 14733 13834 14799 13837
rect 15561 13834 15627 13837
rect 14733 13832 15627 13834
rect 14733 13776 14738 13832
rect 14794 13776 15566 13832
rect 15622 13776 15627 13832
rect 14733 13774 15627 13776
rect 14733 13771 14799 13774
rect 15561 13771 15627 13774
rect 17350 13772 17356 13836
rect 17420 13834 17426 13836
rect 18781 13834 18847 13837
rect 17420 13832 18847 13834
rect 17420 13776 18786 13832
rect 18842 13776 18847 13832
rect 17420 13774 18847 13776
rect 17420 13772 17426 13774
rect 15561 13698 15627 13701
rect 17358 13698 17418 13772
rect 18781 13771 18847 13774
rect 15561 13696 17418 13698
rect 15561 13640 15566 13696
rect 15622 13640 17418 13696
rect 15561 13638 17418 13640
rect 17585 13698 17651 13701
rect 18965 13698 19031 13701
rect 17585 13696 19031 13698
rect 17585 13640 17590 13696
rect 17646 13640 18970 13696
rect 19026 13640 19031 13696
rect 17585 13638 19031 13640
rect 15561 13635 15627 13638
rect 17585 13635 17651 13638
rect 18965 13635 19031 13638
rect 20069 13698 20135 13701
rect 22001 13698 22067 13701
rect 26233 13698 26299 13701
rect 20069 13696 22067 13698
rect 20069 13640 20074 13696
rect 20130 13640 22006 13696
rect 22062 13640 22067 13696
rect 20069 13638 22067 13640
rect 20069 13635 20135 13638
rect 22001 13635 22067 13638
rect 24350 13696 26299 13698
rect 24350 13640 26238 13696
rect 26294 13640 26299 13696
rect 24350 13638 26299 13640
rect 7206 13632 7522 13633
rect 7206 13568 7212 13632
rect 7276 13568 7292 13632
rect 7356 13568 7372 13632
rect 7436 13568 7452 13632
rect 7516 13568 7522 13632
rect 7206 13567 7522 13568
rect 15095 13632 15411 13633
rect 15095 13568 15101 13632
rect 15165 13568 15181 13632
rect 15245 13568 15261 13632
rect 15325 13568 15341 13632
rect 15405 13568 15411 13632
rect 15095 13567 15411 13568
rect 22984 13632 23300 13633
rect 22984 13568 22990 13632
rect 23054 13568 23070 13632
rect 23134 13568 23150 13632
rect 23214 13568 23230 13632
rect 23294 13568 23300 13632
rect 22984 13567 23300 13568
rect 16297 13426 16363 13429
rect 17309 13426 17375 13429
rect 16297 13424 17375 13426
rect 16297 13368 16302 13424
rect 16358 13368 17314 13424
rect 17370 13368 17375 13424
rect 16297 13366 17375 13368
rect 16297 13363 16363 13366
rect 17309 13363 17375 13366
rect 15193 13290 15259 13293
rect 24350 13290 24410 13638
rect 26233 13635 26299 13638
rect 35157 13698 35223 13701
rect 36302 13698 37102 13728
rect 35157 13696 37102 13698
rect 35157 13640 35162 13696
rect 35218 13640 37102 13696
rect 35157 13638 37102 13640
rect 35157 13635 35223 13638
rect 30873 13632 31189 13633
rect 30873 13568 30879 13632
rect 30943 13568 30959 13632
rect 31023 13568 31039 13632
rect 31103 13568 31119 13632
rect 31183 13568 31189 13632
rect 36302 13608 37102 13638
rect 30873 13567 31189 13568
rect 15193 13288 24410 13290
rect 15193 13232 15198 13288
rect 15254 13232 24410 13288
rect 15193 13230 24410 13232
rect 15193 13227 15259 13230
rect 16573 13154 16639 13157
rect 17125 13154 17191 13157
rect 16573 13152 17191 13154
rect 16573 13096 16578 13152
rect 16634 13096 17130 13152
rect 17186 13096 17191 13152
rect 16573 13094 17191 13096
rect 16573 13091 16639 13094
rect 17125 13091 17191 13094
rect 6546 13088 6862 13089
rect 0 13018 800 13048
rect 6546 13024 6552 13088
rect 6616 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6862 13088
rect 6546 13023 6862 13024
rect 14435 13088 14751 13089
rect 14435 13024 14441 13088
rect 14505 13024 14521 13088
rect 14585 13024 14601 13088
rect 14665 13024 14681 13088
rect 14745 13024 14751 13088
rect 14435 13023 14751 13024
rect 22324 13088 22640 13089
rect 22324 13024 22330 13088
rect 22394 13024 22410 13088
rect 22474 13024 22490 13088
rect 22554 13024 22570 13088
rect 22634 13024 22640 13088
rect 22324 13023 22640 13024
rect 30213 13088 30529 13089
rect 30213 13024 30219 13088
rect 30283 13024 30299 13088
rect 30363 13024 30379 13088
rect 30443 13024 30459 13088
rect 30523 13024 30529 13088
rect 30213 13023 30529 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 16849 13018 16915 13021
rect 17953 13018 18019 13021
rect 16849 13016 18019 13018
rect 16849 12960 16854 13016
rect 16910 12960 17958 13016
rect 18014 12960 18019 13016
rect 16849 12958 18019 12960
rect 16849 12955 16915 12958
rect 17953 12955 18019 12958
rect 15469 12882 15535 12885
rect 27838 12882 27844 12884
rect 15469 12880 27844 12882
rect 15469 12824 15474 12880
rect 15530 12824 27844 12880
rect 15469 12822 27844 12824
rect 15469 12819 15535 12822
rect 27838 12820 27844 12822
rect 27908 12820 27914 12884
rect 17401 12746 17467 12749
rect 18689 12746 18755 12749
rect 17401 12744 18755 12746
rect 17401 12688 17406 12744
rect 17462 12688 18694 12744
rect 18750 12688 18755 12744
rect 17401 12686 18755 12688
rect 17401 12683 17467 12686
rect 18689 12683 18755 12686
rect 7206 12544 7522 12545
rect 7206 12480 7212 12544
rect 7276 12480 7292 12544
rect 7356 12480 7372 12544
rect 7436 12480 7452 12544
rect 7516 12480 7522 12544
rect 7206 12479 7522 12480
rect 15095 12544 15411 12545
rect 15095 12480 15101 12544
rect 15165 12480 15181 12544
rect 15245 12480 15261 12544
rect 15325 12480 15341 12544
rect 15405 12480 15411 12544
rect 15095 12479 15411 12480
rect 22984 12544 23300 12545
rect 22984 12480 22990 12544
rect 23054 12480 23070 12544
rect 23134 12480 23150 12544
rect 23214 12480 23230 12544
rect 23294 12480 23300 12544
rect 22984 12479 23300 12480
rect 30873 12544 31189 12545
rect 30873 12480 30879 12544
rect 30943 12480 30959 12544
rect 31023 12480 31039 12544
rect 31103 12480 31119 12544
rect 31183 12480 31189 12544
rect 30873 12479 31189 12480
rect 18045 12338 18111 12341
rect 18413 12338 18479 12341
rect 18045 12336 18479 12338
rect 18045 12280 18050 12336
rect 18106 12280 18418 12336
rect 18474 12280 18479 12336
rect 18045 12278 18479 12280
rect 18045 12275 18111 12278
rect 18413 12275 18479 12278
rect 19517 12338 19583 12341
rect 23565 12338 23631 12341
rect 31937 12338 32003 12341
rect 32673 12338 32739 12341
rect 19517 12336 32003 12338
rect 19517 12280 19522 12336
rect 19578 12280 23570 12336
rect 23626 12280 31942 12336
rect 31998 12280 32003 12336
rect 19517 12278 32003 12280
rect 19517 12275 19583 12278
rect 23565 12275 23631 12278
rect 31937 12275 32003 12278
rect 32078 12336 32739 12338
rect 32078 12280 32678 12336
rect 32734 12280 32739 12336
rect 32078 12278 32739 12280
rect 15469 12202 15535 12205
rect 32078 12202 32138 12278
rect 32673 12275 32739 12278
rect 34421 12338 34487 12341
rect 36302 12338 37102 12368
rect 34421 12336 37102 12338
rect 34421 12280 34426 12336
rect 34482 12280 37102 12336
rect 34421 12278 37102 12280
rect 34421 12275 34487 12278
rect 36302 12248 37102 12278
rect 15469 12200 32138 12202
rect 15469 12144 15474 12200
rect 15530 12144 32138 12200
rect 15469 12142 32138 12144
rect 15469 12139 15535 12142
rect 6546 12000 6862 12001
rect 6546 11936 6552 12000
rect 6616 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6862 12000
rect 6546 11935 6862 11936
rect 14435 12000 14751 12001
rect 14435 11936 14441 12000
rect 14505 11936 14521 12000
rect 14585 11936 14601 12000
rect 14665 11936 14681 12000
rect 14745 11936 14751 12000
rect 14435 11935 14751 11936
rect 22324 12000 22640 12001
rect 22324 11936 22330 12000
rect 22394 11936 22410 12000
rect 22474 11936 22490 12000
rect 22554 11936 22570 12000
rect 22634 11936 22640 12000
rect 22324 11935 22640 11936
rect 30213 12000 30529 12001
rect 30213 11936 30219 12000
rect 30283 11936 30299 12000
rect 30363 11936 30379 12000
rect 30443 11936 30459 12000
rect 30523 11936 30529 12000
rect 30213 11935 30529 11936
rect 17401 11930 17467 11933
rect 19241 11930 19307 11933
rect 17401 11928 19307 11930
rect 17401 11872 17406 11928
rect 17462 11872 19246 11928
rect 19302 11872 19307 11928
rect 17401 11870 19307 11872
rect 17401 11867 17467 11870
rect 19241 11867 19307 11870
rect 13905 11794 13971 11797
rect 18045 11794 18111 11797
rect 13905 11792 18111 11794
rect 13905 11736 13910 11792
rect 13966 11736 18050 11792
rect 18106 11736 18111 11792
rect 13905 11734 18111 11736
rect 13905 11731 13971 11734
rect 18045 11731 18111 11734
rect 21265 11794 21331 11797
rect 28257 11794 28323 11797
rect 21265 11792 28323 11794
rect 21265 11736 21270 11792
rect 21326 11736 28262 11792
rect 28318 11736 28323 11792
rect 21265 11734 28323 11736
rect 21265 11731 21331 11734
rect 28257 11731 28323 11734
rect 0 11658 800 11688
rect 1301 11658 1367 11661
rect 0 11656 1367 11658
rect 0 11600 1306 11656
rect 1362 11600 1367 11656
rect 0 11598 1367 11600
rect 0 11568 800 11598
rect 1301 11595 1367 11598
rect 19333 11658 19399 11661
rect 22001 11658 22067 11661
rect 22185 11660 22251 11661
rect 19333 11656 22067 11658
rect 19333 11600 19338 11656
rect 19394 11600 22006 11656
rect 22062 11600 22067 11656
rect 19333 11598 22067 11600
rect 19333 11595 19399 11598
rect 22001 11595 22067 11598
rect 22134 11596 22140 11660
rect 22204 11658 22251 11660
rect 22204 11656 22296 11658
rect 22246 11600 22296 11656
rect 22204 11598 22296 11600
rect 22204 11596 22251 11598
rect 22185 11595 22251 11596
rect 7206 11456 7522 11457
rect 7206 11392 7212 11456
rect 7276 11392 7292 11456
rect 7356 11392 7372 11456
rect 7436 11392 7452 11456
rect 7516 11392 7522 11456
rect 7206 11391 7522 11392
rect 15095 11456 15411 11457
rect 15095 11392 15101 11456
rect 15165 11392 15181 11456
rect 15245 11392 15261 11456
rect 15325 11392 15341 11456
rect 15405 11392 15411 11456
rect 15095 11391 15411 11392
rect 22984 11456 23300 11457
rect 22984 11392 22990 11456
rect 23054 11392 23070 11456
rect 23134 11392 23150 11456
rect 23214 11392 23230 11456
rect 23294 11392 23300 11456
rect 22984 11391 23300 11392
rect 30873 11456 31189 11457
rect 30873 11392 30879 11456
rect 30943 11392 30959 11456
rect 31023 11392 31039 11456
rect 31103 11392 31119 11456
rect 31183 11392 31189 11456
rect 30873 11391 31189 11392
rect 15929 11250 15995 11253
rect 17585 11250 17651 11253
rect 15929 11248 17651 11250
rect 15929 11192 15934 11248
rect 15990 11192 17590 11248
rect 17646 11192 17651 11248
rect 15929 11190 17651 11192
rect 15929 11187 15995 11190
rect 17585 11187 17651 11190
rect 12157 11114 12223 11117
rect 14733 11114 14799 11117
rect 12157 11112 14799 11114
rect 12157 11056 12162 11112
rect 12218 11056 14738 11112
rect 14794 11056 14799 11112
rect 12157 11054 14799 11056
rect 12157 11051 12223 11054
rect 14733 11051 14799 11054
rect 16941 10978 17007 10981
rect 19558 10978 19564 10980
rect 16941 10976 19564 10978
rect 16941 10920 16946 10976
rect 17002 10920 19564 10976
rect 16941 10918 19564 10920
rect 16941 10915 17007 10918
rect 19558 10916 19564 10918
rect 19628 10916 19634 10980
rect 34881 10978 34947 10981
rect 36302 10978 37102 11008
rect 34881 10976 37102 10978
rect 34881 10920 34886 10976
rect 34942 10920 37102 10976
rect 34881 10918 37102 10920
rect 34881 10915 34947 10918
rect 6546 10912 6862 10913
rect 6546 10848 6552 10912
rect 6616 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6862 10912
rect 6546 10847 6862 10848
rect 14435 10912 14751 10913
rect 14435 10848 14441 10912
rect 14505 10848 14521 10912
rect 14585 10848 14601 10912
rect 14665 10848 14681 10912
rect 14745 10848 14751 10912
rect 14435 10847 14751 10848
rect 22324 10912 22640 10913
rect 22324 10848 22330 10912
rect 22394 10848 22410 10912
rect 22474 10848 22490 10912
rect 22554 10848 22570 10912
rect 22634 10848 22640 10912
rect 22324 10847 22640 10848
rect 30213 10912 30529 10913
rect 30213 10848 30219 10912
rect 30283 10848 30299 10912
rect 30363 10848 30379 10912
rect 30443 10848 30459 10912
rect 30523 10848 30529 10912
rect 36302 10888 37102 10918
rect 30213 10847 30529 10848
rect 7206 10368 7522 10369
rect 7206 10304 7212 10368
rect 7276 10304 7292 10368
rect 7356 10304 7372 10368
rect 7436 10304 7452 10368
rect 7516 10304 7522 10368
rect 7206 10303 7522 10304
rect 15095 10368 15411 10369
rect 15095 10304 15101 10368
rect 15165 10304 15181 10368
rect 15245 10304 15261 10368
rect 15325 10304 15341 10368
rect 15405 10304 15411 10368
rect 15095 10303 15411 10304
rect 22984 10368 23300 10369
rect 22984 10304 22990 10368
rect 23054 10304 23070 10368
rect 23134 10304 23150 10368
rect 23214 10304 23230 10368
rect 23294 10304 23300 10368
rect 22984 10303 23300 10304
rect 30873 10368 31189 10369
rect 30873 10304 30879 10368
rect 30943 10304 30959 10368
rect 31023 10304 31039 10368
rect 31103 10304 31119 10368
rect 31183 10304 31189 10368
rect 30873 10303 31189 10304
rect 6546 9824 6862 9825
rect 6546 9760 6552 9824
rect 6616 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6862 9824
rect 6546 9759 6862 9760
rect 14435 9824 14751 9825
rect 14435 9760 14441 9824
rect 14505 9760 14521 9824
rect 14585 9760 14601 9824
rect 14665 9760 14681 9824
rect 14745 9760 14751 9824
rect 14435 9759 14751 9760
rect 22324 9824 22640 9825
rect 22324 9760 22330 9824
rect 22394 9760 22410 9824
rect 22474 9760 22490 9824
rect 22554 9760 22570 9824
rect 22634 9760 22640 9824
rect 22324 9759 22640 9760
rect 30213 9824 30529 9825
rect 30213 9760 30219 9824
rect 30283 9760 30299 9824
rect 30363 9760 30379 9824
rect 30443 9760 30459 9824
rect 30523 9760 30529 9824
rect 30213 9759 30529 9760
rect 0 9618 800 9648
rect 1301 9618 1367 9621
rect 5717 9620 5783 9621
rect 5717 9618 5764 9620
rect 0 9616 1367 9618
rect 0 9560 1306 9616
rect 1362 9560 1367 9616
rect 0 9558 1367 9560
rect 5672 9616 5764 9618
rect 5672 9560 5722 9616
rect 5672 9558 5764 9560
rect 0 9528 800 9558
rect 1301 9555 1367 9558
rect 5717 9556 5764 9558
rect 5828 9556 5834 9620
rect 19190 9556 19196 9620
rect 19260 9618 19266 9620
rect 19609 9618 19675 9621
rect 19260 9616 19675 9618
rect 19260 9560 19614 9616
rect 19670 9560 19675 9616
rect 19260 9558 19675 9560
rect 19260 9556 19266 9558
rect 5717 9555 5783 9556
rect 19609 9555 19675 9558
rect 34421 9618 34487 9621
rect 36302 9618 37102 9648
rect 34421 9616 37102 9618
rect 34421 9560 34426 9616
rect 34482 9560 37102 9616
rect 34421 9558 37102 9560
rect 34421 9555 34487 9558
rect 36302 9528 37102 9558
rect 17493 9482 17559 9485
rect 17861 9482 17927 9485
rect 17493 9480 17927 9482
rect 17493 9424 17498 9480
rect 17554 9424 17866 9480
rect 17922 9424 17927 9480
rect 17493 9422 17927 9424
rect 17493 9419 17559 9422
rect 17861 9419 17927 9422
rect 21582 9420 21588 9484
rect 21652 9482 21658 9484
rect 24853 9482 24919 9485
rect 21652 9480 24919 9482
rect 21652 9424 24858 9480
rect 24914 9424 24919 9480
rect 21652 9422 24919 9424
rect 21652 9420 21658 9422
rect 24853 9419 24919 9422
rect 7206 9280 7522 9281
rect 7206 9216 7212 9280
rect 7276 9216 7292 9280
rect 7356 9216 7372 9280
rect 7436 9216 7452 9280
rect 7516 9216 7522 9280
rect 7206 9215 7522 9216
rect 15095 9280 15411 9281
rect 15095 9216 15101 9280
rect 15165 9216 15181 9280
rect 15245 9216 15261 9280
rect 15325 9216 15341 9280
rect 15405 9216 15411 9280
rect 15095 9215 15411 9216
rect 22984 9280 23300 9281
rect 22984 9216 22990 9280
rect 23054 9216 23070 9280
rect 23134 9216 23150 9280
rect 23214 9216 23230 9280
rect 23294 9216 23300 9280
rect 22984 9215 23300 9216
rect 30873 9280 31189 9281
rect 30873 9216 30879 9280
rect 30943 9216 30959 9280
rect 31023 9216 31039 9280
rect 31103 9216 31119 9280
rect 31183 9216 31189 9280
rect 30873 9215 31189 9216
rect 24761 9210 24827 9213
rect 28165 9210 28231 9213
rect 24761 9208 28231 9210
rect 24761 9152 24766 9208
rect 24822 9152 28170 9208
rect 28226 9152 28231 9208
rect 24761 9150 28231 9152
rect 24761 9147 24827 9150
rect 28165 9147 28231 9150
rect 14549 9074 14615 9077
rect 18045 9074 18111 9077
rect 14549 9072 18111 9074
rect 14549 9016 14554 9072
rect 14610 9016 18050 9072
rect 18106 9016 18111 9072
rect 14549 9014 18111 9016
rect 14549 9011 14615 9014
rect 18045 9011 18111 9014
rect 18781 9074 18847 9077
rect 33777 9074 33843 9077
rect 18781 9072 33843 9074
rect 18781 9016 18786 9072
rect 18842 9016 33782 9072
rect 33838 9016 33843 9072
rect 18781 9014 33843 9016
rect 18781 9011 18847 9014
rect 33777 9011 33843 9014
rect 22093 8938 22159 8941
rect 26233 8938 26299 8941
rect 22093 8936 26299 8938
rect 22093 8880 22098 8936
rect 22154 8880 26238 8936
rect 26294 8880 26299 8936
rect 22093 8878 26299 8880
rect 22093 8875 22159 8878
rect 26233 8875 26299 8878
rect 6546 8736 6862 8737
rect 6546 8672 6552 8736
rect 6616 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6862 8736
rect 6546 8671 6862 8672
rect 14435 8736 14751 8737
rect 14435 8672 14441 8736
rect 14505 8672 14521 8736
rect 14585 8672 14601 8736
rect 14665 8672 14681 8736
rect 14745 8672 14751 8736
rect 14435 8671 14751 8672
rect 22324 8736 22640 8737
rect 22324 8672 22330 8736
rect 22394 8672 22410 8736
rect 22474 8672 22490 8736
rect 22554 8672 22570 8736
rect 22634 8672 22640 8736
rect 22324 8671 22640 8672
rect 30213 8736 30529 8737
rect 30213 8672 30219 8736
rect 30283 8672 30299 8736
rect 30363 8672 30379 8736
rect 30443 8672 30459 8736
rect 30523 8672 30529 8736
rect 30213 8671 30529 8672
rect 26325 8666 26391 8669
rect 22878 8664 26391 8666
rect 22878 8608 26330 8664
rect 26386 8608 26391 8664
rect 22878 8606 26391 8608
rect 21909 8530 21975 8533
rect 22878 8530 22938 8606
rect 26325 8603 26391 8606
rect 21909 8528 22938 8530
rect 21909 8472 21914 8528
rect 21970 8472 22938 8528
rect 21909 8470 22938 8472
rect 23105 8530 23171 8533
rect 33777 8530 33843 8533
rect 23105 8528 33843 8530
rect 23105 8472 23110 8528
rect 23166 8472 33782 8528
rect 33838 8472 33843 8528
rect 23105 8470 33843 8472
rect 21909 8467 21975 8470
rect 23105 8467 23171 8470
rect 33777 8467 33843 8470
rect 23381 8394 23447 8397
rect 28993 8394 29059 8397
rect 23381 8392 29059 8394
rect 23381 8336 23386 8392
rect 23442 8336 28998 8392
rect 29054 8336 29059 8392
rect 23381 8334 29059 8336
rect 23381 8331 23447 8334
rect 28993 8331 29059 8334
rect 0 8258 800 8288
rect 1301 8258 1367 8261
rect 18781 8260 18847 8261
rect 18781 8258 18828 8260
rect 0 8256 1367 8258
rect 0 8200 1306 8256
rect 1362 8200 1367 8256
rect 0 8198 1367 8200
rect 18736 8256 18828 8258
rect 18736 8200 18786 8256
rect 18736 8198 18828 8200
rect 0 8168 800 8198
rect 1301 8195 1367 8198
rect 18781 8196 18828 8198
rect 18892 8196 18898 8260
rect 34421 8258 34487 8261
rect 36302 8258 37102 8288
rect 34421 8256 37102 8258
rect 34421 8200 34426 8256
rect 34482 8200 37102 8256
rect 34421 8198 37102 8200
rect 18781 8195 18847 8196
rect 34421 8195 34487 8198
rect 7206 8192 7522 8193
rect 7206 8128 7212 8192
rect 7276 8128 7292 8192
rect 7356 8128 7372 8192
rect 7436 8128 7452 8192
rect 7516 8128 7522 8192
rect 7206 8127 7522 8128
rect 15095 8192 15411 8193
rect 15095 8128 15101 8192
rect 15165 8128 15181 8192
rect 15245 8128 15261 8192
rect 15325 8128 15341 8192
rect 15405 8128 15411 8192
rect 15095 8127 15411 8128
rect 22984 8192 23300 8193
rect 22984 8128 22990 8192
rect 23054 8128 23070 8192
rect 23134 8128 23150 8192
rect 23214 8128 23230 8192
rect 23294 8128 23300 8192
rect 22984 8127 23300 8128
rect 30873 8192 31189 8193
rect 30873 8128 30879 8192
rect 30943 8128 30959 8192
rect 31023 8128 31039 8192
rect 31103 8128 31119 8192
rect 31183 8128 31189 8192
rect 36302 8168 37102 8198
rect 30873 8127 31189 8128
rect 18597 8122 18663 8125
rect 19374 8122 19380 8124
rect 18597 8120 19380 8122
rect 18597 8064 18602 8120
rect 18658 8064 19380 8120
rect 18597 8062 19380 8064
rect 18597 8059 18663 8062
rect 19374 8060 19380 8062
rect 19444 8060 19450 8124
rect 29269 8122 29335 8125
rect 30557 8122 30623 8125
rect 29269 8120 30623 8122
rect 29269 8064 29274 8120
rect 29330 8064 30562 8120
rect 30618 8064 30623 8120
rect 29269 8062 30623 8064
rect 29269 8059 29335 8062
rect 30557 8059 30623 8062
rect 9213 7986 9279 7989
rect 26550 7986 26556 7988
rect 9213 7984 26556 7986
rect 9213 7928 9218 7984
rect 9274 7928 26556 7984
rect 9213 7926 26556 7928
rect 9213 7923 9279 7926
rect 26550 7924 26556 7926
rect 26620 7924 26626 7988
rect 4061 7850 4127 7853
rect 8661 7850 8727 7853
rect 4061 7848 8727 7850
rect 4061 7792 4066 7848
rect 4122 7792 8666 7848
rect 8722 7792 8727 7848
rect 4061 7790 8727 7792
rect 4061 7787 4127 7790
rect 8661 7787 8727 7790
rect 6546 7648 6862 7649
rect 6546 7584 6552 7648
rect 6616 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6862 7648
rect 6546 7583 6862 7584
rect 14435 7648 14751 7649
rect 14435 7584 14441 7648
rect 14505 7584 14521 7648
rect 14585 7584 14601 7648
rect 14665 7584 14681 7648
rect 14745 7584 14751 7648
rect 14435 7583 14751 7584
rect 22324 7648 22640 7649
rect 22324 7584 22330 7648
rect 22394 7584 22410 7648
rect 22474 7584 22490 7648
rect 22554 7584 22570 7648
rect 22634 7584 22640 7648
rect 22324 7583 22640 7584
rect 30213 7648 30529 7649
rect 30213 7584 30219 7648
rect 30283 7584 30299 7648
rect 30363 7584 30379 7648
rect 30443 7584 30459 7648
rect 30523 7584 30529 7648
rect 30213 7583 30529 7584
rect 7206 7104 7522 7105
rect 7206 7040 7212 7104
rect 7276 7040 7292 7104
rect 7356 7040 7372 7104
rect 7436 7040 7452 7104
rect 7516 7040 7522 7104
rect 7206 7039 7522 7040
rect 15095 7104 15411 7105
rect 15095 7040 15101 7104
rect 15165 7040 15181 7104
rect 15245 7040 15261 7104
rect 15325 7040 15341 7104
rect 15405 7040 15411 7104
rect 15095 7039 15411 7040
rect 22984 7104 23300 7105
rect 22984 7040 22990 7104
rect 23054 7040 23070 7104
rect 23134 7040 23150 7104
rect 23214 7040 23230 7104
rect 23294 7040 23300 7104
rect 22984 7039 23300 7040
rect 30873 7104 31189 7105
rect 30873 7040 30879 7104
rect 30943 7040 30959 7104
rect 31023 7040 31039 7104
rect 31103 7040 31119 7104
rect 31183 7040 31189 7104
rect 30873 7039 31189 7040
rect 0 6898 800 6928
rect 3509 6898 3575 6901
rect 0 6896 3575 6898
rect 0 6840 3514 6896
rect 3570 6840 3575 6896
rect 0 6838 3575 6840
rect 0 6808 800 6838
rect 3509 6835 3575 6838
rect 24117 6898 24183 6901
rect 28625 6898 28691 6901
rect 24117 6896 28691 6898
rect 24117 6840 24122 6896
rect 24178 6840 28630 6896
rect 28686 6840 28691 6896
rect 24117 6838 28691 6840
rect 24117 6835 24183 6838
rect 28625 6835 28691 6838
rect 34697 6898 34763 6901
rect 36302 6898 37102 6928
rect 34697 6896 37102 6898
rect 34697 6840 34702 6896
rect 34758 6840 37102 6896
rect 34697 6838 37102 6840
rect 34697 6835 34763 6838
rect 36302 6808 37102 6838
rect 6546 6560 6862 6561
rect 6546 6496 6552 6560
rect 6616 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6862 6560
rect 6546 6495 6862 6496
rect 14435 6560 14751 6561
rect 14435 6496 14441 6560
rect 14505 6496 14521 6560
rect 14585 6496 14601 6560
rect 14665 6496 14681 6560
rect 14745 6496 14751 6560
rect 14435 6495 14751 6496
rect 22324 6560 22640 6561
rect 22324 6496 22330 6560
rect 22394 6496 22410 6560
rect 22474 6496 22490 6560
rect 22554 6496 22570 6560
rect 22634 6496 22640 6560
rect 22324 6495 22640 6496
rect 30213 6560 30529 6561
rect 30213 6496 30219 6560
rect 30283 6496 30299 6560
rect 30363 6496 30379 6560
rect 30443 6496 30459 6560
rect 30523 6496 30529 6560
rect 30213 6495 30529 6496
rect 19333 6354 19399 6357
rect 26969 6354 27035 6357
rect 19333 6352 27035 6354
rect 19333 6296 19338 6352
rect 19394 6296 26974 6352
rect 27030 6296 27035 6352
rect 19333 6294 27035 6296
rect 19333 6291 19399 6294
rect 26969 6291 27035 6294
rect 4061 6218 4127 6221
rect 24853 6218 24919 6221
rect 4061 6216 24919 6218
rect 4061 6160 4066 6216
rect 4122 6160 24858 6216
rect 24914 6160 24919 6216
rect 4061 6158 24919 6160
rect 4061 6155 4127 6158
rect 24853 6155 24919 6158
rect 7206 6016 7522 6017
rect 7206 5952 7212 6016
rect 7276 5952 7292 6016
rect 7356 5952 7372 6016
rect 7436 5952 7452 6016
rect 7516 5952 7522 6016
rect 7206 5951 7522 5952
rect 15095 6016 15411 6017
rect 15095 5952 15101 6016
rect 15165 5952 15181 6016
rect 15245 5952 15261 6016
rect 15325 5952 15341 6016
rect 15405 5952 15411 6016
rect 15095 5951 15411 5952
rect 22984 6016 23300 6017
rect 22984 5952 22990 6016
rect 23054 5952 23070 6016
rect 23134 5952 23150 6016
rect 23214 5952 23230 6016
rect 23294 5952 23300 6016
rect 22984 5951 23300 5952
rect 30873 6016 31189 6017
rect 30873 5952 30879 6016
rect 30943 5952 30959 6016
rect 31023 5952 31039 6016
rect 31103 5952 31119 6016
rect 31183 5952 31189 6016
rect 30873 5951 31189 5952
rect 25405 5810 25471 5813
rect 34053 5810 34119 5813
rect 25405 5808 34119 5810
rect 25405 5752 25410 5808
rect 25466 5752 34058 5808
rect 34114 5752 34119 5808
rect 25405 5750 34119 5752
rect 25405 5747 25471 5750
rect 34053 5747 34119 5750
rect 12157 5674 12223 5677
rect 16665 5674 16731 5677
rect 12157 5672 16731 5674
rect 12157 5616 12162 5672
rect 12218 5616 16670 5672
rect 16726 5616 16731 5672
rect 12157 5614 16731 5616
rect 12157 5611 12223 5614
rect 16665 5611 16731 5614
rect 28165 5674 28231 5677
rect 32213 5674 32279 5677
rect 28165 5672 32279 5674
rect 28165 5616 28170 5672
rect 28226 5616 32218 5672
rect 32274 5616 32279 5672
rect 28165 5614 32279 5616
rect 28165 5611 28231 5614
rect 32213 5611 32279 5614
rect 0 5538 800 5568
rect 3049 5538 3115 5541
rect 0 5536 3115 5538
rect 0 5480 3054 5536
rect 3110 5480 3115 5536
rect 0 5478 3115 5480
rect 0 5448 800 5478
rect 3049 5475 3115 5478
rect 34881 5538 34947 5541
rect 36302 5538 37102 5568
rect 34881 5536 37102 5538
rect 34881 5480 34886 5536
rect 34942 5480 37102 5536
rect 34881 5478 37102 5480
rect 34881 5475 34947 5478
rect 6546 5472 6862 5473
rect 6546 5408 6552 5472
rect 6616 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6862 5472
rect 6546 5407 6862 5408
rect 14435 5472 14751 5473
rect 14435 5408 14441 5472
rect 14505 5408 14521 5472
rect 14585 5408 14601 5472
rect 14665 5408 14681 5472
rect 14745 5408 14751 5472
rect 14435 5407 14751 5408
rect 22324 5472 22640 5473
rect 22324 5408 22330 5472
rect 22394 5408 22410 5472
rect 22474 5408 22490 5472
rect 22554 5408 22570 5472
rect 22634 5408 22640 5472
rect 22324 5407 22640 5408
rect 30213 5472 30529 5473
rect 30213 5408 30219 5472
rect 30283 5408 30299 5472
rect 30363 5408 30379 5472
rect 30443 5408 30459 5472
rect 30523 5408 30529 5472
rect 36302 5448 37102 5478
rect 30213 5407 30529 5408
rect 7206 4928 7522 4929
rect 7206 4864 7212 4928
rect 7276 4864 7292 4928
rect 7356 4864 7372 4928
rect 7436 4864 7452 4928
rect 7516 4864 7522 4928
rect 7206 4863 7522 4864
rect 15095 4928 15411 4929
rect 15095 4864 15101 4928
rect 15165 4864 15181 4928
rect 15245 4864 15261 4928
rect 15325 4864 15341 4928
rect 15405 4864 15411 4928
rect 15095 4863 15411 4864
rect 22984 4928 23300 4929
rect 22984 4864 22990 4928
rect 23054 4864 23070 4928
rect 23134 4864 23150 4928
rect 23214 4864 23230 4928
rect 23294 4864 23300 4928
rect 22984 4863 23300 4864
rect 30873 4928 31189 4929
rect 30873 4864 30879 4928
rect 30943 4864 30959 4928
rect 31023 4864 31039 4928
rect 31103 4864 31119 4928
rect 31183 4864 31189 4928
rect 30873 4863 31189 4864
rect 6546 4384 6862 4385
rect 6546 4320 6552 4384
rect 6616 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6862 4384
rect 6546 4319 6862 4320
rect 14435 4384 14751 4385
rect 14435 4320 14441 4384
rect 14505 4320 14521 4384
rect 14585 4320 14601 4384
rect 14665 4320 14681 4384
rect 14745 4320 14751 4384
rect 14435 4319 14751 4320
rect 22324 4384 22640 4385
rect 22324 4320 22330 4384
rect 22394 4320 22410 4384
rect 22474 4320 22490 4384
rect 22554 4320 22570 4384
rect 22634 4320 22640 4384
rect 22324 4319 22640 4320
rect 30213 4384 30529 4385
rect 30213 4320 30219 4384
rect 30283 4320 30299 4384
rect 30363 4320 30379 4384
rect 30443 4320 30459 4384
rect 30523 4320 30529 4384
rect 30213 4319 30529 4320
rect 0 4178 800 4208
rect 1301 4178 1367 4181
rect 0 4176 1367 4178
rect 0 4120 1306 4176
rect 1362 4120 1367 4176
rect 0 4118 1367 4120
rect 0 4088 800 4118
rect 1301 4115 1367 4118
rect 34697 4178 34763 4181
rect 36302 4178 37102 4208
rect 34697 4176 37102 4178
rect 34697 4120 34702 4176
rect 34758 4120 37102 4176
rect 34697 4118 37102 4120
rect 34697 4115 34763 4118
rect 36302 4088 37102 4118
rect 7206 3840 7522 3841
rect 7206 3776 7212 3840
rect 7276 3776 7292 3840
rect 7356 3776 7372 3840
rect 7436 3776 7452 3840
rect 7516 3776 7522 3840
rect 7206 3775 7522 3776
rect 15095 3840 15411 3841
rect 15095 3776 15101 3840
rect 15165 3776 15181 3840
rect 15245 3776 15261 3840
rect 15325 3776 15341 3840
rect 15405 3776 15411 3840
rect 15095 3775 15411 3776
rect 22984 3840 23300 3841
rect 22984 3776 22990 3840
rect 23054 3776 23070 3840
rect 23134 3776 23150 3840
rect 23214 3776 23230 3840
rect 23294 3776 23300 3840
rect 22984 3775 23300 3776
rect 30873 3840 31189 3841
rect 30873 3776 30879 3840
rect 30943 3776 30959 3840
rect 31023 3776 31039 3840
rect 31103 3776 31119 3840
rect 31183 3776 31189 3840
rect 30873 3775 31189 3776
rect 6546 3296 6862 3297
rect 6546 3232 6552 3296
rect 6616 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6862 3296
rect 6546 3231 6862 3232
rect 14435 3296 14751 3297
rect 14435 3232 14441 3296
rect 14505 3232 14521 3296
rect 14585 3232 14601 3296
rect 14665 3232 14681 3296
rect 14745 3232 14751 3296
rect 14435 3231 14751 3232
rect 22324 3296 22640 3297
rect 22324 3232 22330 3296
rect 22394 3232 22410 3296
rect 22474 3232 22490 3296
rect 22554 3232 22570 3296
rect 22634 3232 22640 3296
rect 22324 3231 22640 3232
rect 30213 3296 30529 3297
rect 30213 3232 30219 3296
rect 30283 3232 30299 3296
rect 30363 3232 30379 3296
rect 30443 3232 30459 3296
rect 30523 3232 30529 3296
rect 30213 3231 30529 3232
rect 5717 3090 5783 3093
rect 15694 3090 15700 3092
rect 5717 3088 15700 3090
rect 5717 3032 5722 3088
rect 5778 3032 15700 3088
rect 5717 3030 15700 3032
rect 5717 3027 5783 3030
rect 15694 3028 15700 3030
rect 15764 3028 15770 3092
rect 0 2818 800 2848
rect 1301 2818 1367 2821
rect 0 2816 1367 2818
rect 0 2760 1306 2816
rect 1362 2760 1367 2816
rect 0 2758 1367 2760
rect 0 2728 800 2758
rect 1301 2755 1367 2758
rect 7206 2752 7522 2753
rect 7206 2688 7212 2752
rect 7276 2688 7292 2752
rect 7356 2688 7372 2752
rect 7436 2688 7452 2752
rect 7516 2688 7522 2752
rect 7206 2687 7522 2688
rect 15095 2752 15411 2753
rect 15095 2688 15101 2752
rect 15165 2688 15181 2752
rect 15245 2688 15261 2752
rect 15325 2688 15341 2752
rect 15405 2688 15411 2752
rect 15095 2687 15411 2688
rect 22984 2752 23300 2753
rect 22984 2688 22990 2752
rect 23054 2688 23070 2752
rect 23134 2688 23150 2752
rect 23214 2688 23230 2752
rect 23294 2688 23300 2752
rect 22984 2687 23300 2688
rect 30873 2752 31189 2753
rect 30873 2688 30879 2752
rect 30943 2688 30959 2752
rect 31023 2688 31039 2752
rect 31103 2688 31119 2752
rect 31183 2688 31189 2752
rect 30873 2687 31189 2688
rect 34421 2138 34487 2141
rect 36302 2138 37102 2168
rect 34421 2136 37102 2138
rect 34421 2080 34426 2136
rect 34482 2080 37102 2136
rect 34421 2078 37102 2080
rect 34421 2075 34487 2078
rect 36302 2048 37102 2078
rect 0 1458 800 1488
rect 3049 1458 3115 1461
rect 0 1456 3115 1458
rect 0 1400 3054 1456
rect 3110 1400 3115 1456
rect 0 1398 3115 1400
rect 0 1368 800 1398
rect 3049 1395 3115 1398
rect 33041 914 33107 917
rect 33041 912 33610 914
rect 33041 856 33046 912
rect 33102 856 33610 912
rect 33041 854 33610 856
rect 33041 851 33107 854
rect 33550 778 33610 854
rect 36302 778 37102 808
rect 33550 718 37102 778
rect 36302 688 37102 718
<< via3 >>
rect 7212 34300 7276 34304
rect 7212 34244 7216 34300
rect 7216 34244 7272 34300
rect 7272 34244 7276 34300
rect 7212 34240 7276 34244
rect 7292 34300 7356 34304
rect 7292 34244 7296 34300
rect 7296 34244 7352 34300
rect 7352 34244 7356 34300
rect 7292 34240 7356 34244
rect 7372 34300 7436 34304
rect 7372 34244 7376 34300
rect 7376 34244 7432 34300
rect 7432 34244 7436 34300
rect 7372 34240 7436 34244
rect 7452 34300 7516 34304
rect 7452 34244 7456 34300
rect 7456 34244 7512 34300
rect 7512 34244 7516 34300
rect 7452 34240 7516 34244
rect 15101 34300 15165 34304
rect 15101 34244 15105 34300
rect 15105 34244 15161 34300
rect 15161 34244 15165 34300
rect 15101 34240 15165 34244
rect 15181 34300 15245 34304
rect 15181 34244 15185 34300
rect 15185 34244 15241 34300
rect 15241 34244 15245 34300
rect 15181 34240 15245 34244
rect 15261 34300 15325 34304
rect 15261 34244 15265 34300
rect 15265 34244 15321 34300
rect 15321 34244 15325 34300
rect 15261 34240 15325 34244
rect 15341 34300 15405 34304
rect 15341 34244 15345 34300
rect 15345 34244 15401 34300
rect 15401 34244 15405 34300
rect 15341 34240 15405 34244
rect 22990 34300 23054 34304
rect 22990 34244 22994 34300
rect 22994 34244 23050 34300
rect 23050 34244 23054 34300
rect 22990 34240 23054 34244
rect 23070 34300 23134 34304
rect 23070 34244 23074 34300
rect 23074 34244 23130 34300
rect 23130 34244 23134 34300
rect 23070 34240 23134 34244
rect 23150 34300 23214 34304
rect 23150 34244 23154 34300
rect 23154 34244 23210 34300
rect 23210 34244 23214 34300
rect 23150 34240 23214 34244
rect 23230 34300 23294 34304
rect 23230 34244 23234 34300
rect 23234 34244 23290 34300
rect 23290 34244 23294 34300
rect 23230 34240 23294 34244
rect 30879 34300 30943 34304
rect 30879 34244 30883 34300
rect 30883 34244 30939 34300
rect 30939 34244 30943 34300
rect 30879 34240 30943 34244
rect 30959 34300 31023 34304
rect 30959 34244 30963 34300
rect 30963 34244 31019 34300
rect 31019 34244 31023 34300
rect 30959 34240 31023 34244
rect 31039 34300 31103 34304
rect 31039 34244 31043 34300
rect 31043 34244 31099 34300
rect 31099 34244 31103 34300
rect 31039 34240 31103 34244
rect 31119 34300 31183 34304
rect 31119 34244 31123 34300
rect 31123 34244 31179 34300
rect 31179 34244 31183 34300
rect 31119 34240 31183 34244
rect 6552 33756 6616 33760
rect 6552 33700 6556 33756
rect 6556 33700 6612 33756
rect 6612 33700 6616 33756
rect 6552 33696 6616 33700
rect 6632 33756 6696 33760
rect 6632 33700 6636 33756
rect 6636 33700 6692 33756
rect 6692 33700 6696 33756
rect 6632 33696 6696 33700
rect 6712 33756 6776 33760
rect 6712 33700 6716 33756
rect 6716 33700 6772 33756
rect 6772 33700 6776 33756
rect 6712 33696 6776 33700
rect 6792 33756 6856 33760
rect 6792 33700 6796 33756
rect 6796 33700 6852 33756
rect 6852 33700 6856 33756
rect 6792 33696 6856 33700
rect 14441 33756 14505 33760
rect 14441 33700 14445 33756
rect 14445 33700 14501 33756
rect 14501 33700 14505 33756
rect 14441 33696 14505 33700
rect 14521 33756 14585 33760
rect 14521 33700 14525 33756
rect 14525 33700 14581 33756
rect 14581 33700 14585 33756
rect 14521 33696 14585 33700
rect 14601 33756 14665 33760
rect 14601 33700 14605 33756
rect 14605 33700 14661 33756
rect 14661 33700 14665 33756
rect 14601 33696 14665 33700
rect 14681 33756 14745 33760
rect 14681 33700 14685 33756
rect 14685 33700 14741 33756
rect 14741 33700 14745 33756
rect 14681 33696 14745 33700
rect 22330 33756 22394 33760
rect 22330 33700 22334 33756
rect 22334 33700 22390 33756
rect 22390 33700 22394 33756
rect 22330 33696 22394 33700
rect 22410 33756 22474 33760
rect 22410 33700 22414 33756
rect 22414 33700 22470 33756
rect 22470 33700 22474 33756
rect 22410 33696 22474 33700
rect 22490 33756 22554 33760
rect 22490 33700 22494 33756
rect 22494 33700 22550 33756
rect 22550 33700 22554 33756
rect 22490 33696 22554 33700
rect 22570 33756 22634 33760
rect 22570 33700 22574 33756
rect 22574 33700 22630 33756
rect 22630 33700 22634 33756
rect 22570 33696 22634 33700
rect 30219 33756 30283 33760
rect 30219 33700 30223 33756
rect 30223 33700 30279 33756
rect 30279 33700 30283 33756
rect 30219 33696 30283 33700
rect 30299 33756 30363 33760
rect 30299 33700 30303 33756
rect 30303 33700 30359 33756
rect 30359 33700 30363 33756
rect 30299 33696 30363 33700
rect 30379 33756 30443 33760
rect 30379 33700 30383 33756
rect 30383 33700 30439 33756
rect 30439 33700 30443 33756
rect 30379 33696 30443 33700
rect 30459 33756 30523 33760
rect 30459 33700 30463 33756
rect 30463 33700 30519 33756
rect 30519 33700 30523 33756
rect 30459 33696 30523 33700
rect 10916 33280 10980 33284
rect 10916 33224 10930 33280
rect 10930 33224 10980 33280
rect 10916 33220 10980 33224
rect 19196 33220 19260 33284
rect 21588 33280 21652 33284
rect 21588 33224 21602 33280
rect 21602 33224 21652 33280
rect 21588 33220 21652 33224
rect 7212 33212 7276 33216
rect 7212 33156 7216 33212
rect 7216 33156 7272 33212
rect 7272 33156 7276 33212
rect 7212 33152 7276 33156
rect 7292 33212 7356 33216
rect 7292 33156 7296 33212
rect 7296 33156 7352 33212
rect 7352 33156 7356 33212
rect 7292 33152 7356 33156
rect 7372 33212 7436 33216
rect 7372 33156 7376 33212
rect 7376 33156 7432 33212
rect 7432 33156 7436 33212
rect 7372 33152 7436 33156
rect 7452 33212 7516 33216
rect 7452 33156 7456 33212
rect 7456 33156 7512 33212
rect 7512 33156 7516 33212
rect 7452 33152 7516 33156
rect 15101 33212 15165 33216
rect 15101 33156 15105 33212
rect 15105 33156 15161 33212
rect 15161 33156 15165 33212
rect 15101 33152 15165 33156
rect 15181 33212 15245 33216
rect 15181 33156 15185 33212
rect 15185 33156 15241 33212
rect 15241 33156 15245 33212
rect 15181 33152 15245 33156
rect 15261 33212 15325 33216
rect 15261 33156 15265 33212
rect 15265 33156 15321 33212
rect 15321 33156 15325 33212
rect 15261 33152 15325 33156
rect 15341 33212 15405 33216
rect 15341 33156 15345 33212
rect 15345 33156 15401 33212
rect 15401 33156 15405 33212
rect 15341 33152 15405 33156
rect 22990 33212 23054 33216
rect 22990 33156 22994 33212
rect 22994 33156 23050 33212
rect 23050 33156 23054 33212
rect 22990 33152 23054 33156
rect 23070 33212 23134 33216
rect 23070 33156 23074 33212
rect 23074 33156 23130 33212
rect 23130 33156 23134 33212
rect 23070 33152 23134 33156
rect 23150 33212 23214 33216
rect 23150 33156 23154 33212
rect 23154 33156 23210 33212
rect 23210 33156 23214 33212
rect 23150 33152 23214 33156
rect 23230 33212 23294 33216
rect 23230 33156 23234 33212
rect 23234 33156 23290 33212
rect 23290 33156 23294 33212
rect 23230 33152 23294 33156
rect 30879 33212 30943 33216
rect 30879 33156 30883 33212
rect 30883 33156 30939 33212
rect 30939 33156 30943 33212
rect 30879 33152 30943 33156
rect 30959 33212 31023 33216
rect 30959 33156 30963 33212
rect 30963 33156 31019 33212
rect 31019 33156 31023 33212
rect 30959 33152 31023 33156
rect 31039 33212 31103 33216
rect 31039 33156 31043 33212
rect 31043 33156 31099 33212
rect 31099 33156 31103 33212
rect 31039 33152 31103 33156
rect 31119 33212 31183 33216
rect 31119 33156 31123 33212
rect 31123 33156 31179 33212
rect 31179 33156 31183 33212
rect 31119 33152 31183 33156
rect 12204 33084 12268 33148
rect 6552 32668 6616 32672
rect 6552 32612 6556 32668
rect 6556 32612 6612 32668
rect 6612 32612 6616 32668
rect 6552 32608 6616 32612
rect 6632 32668 6696 32672
rect 6632 32612 6636 32668
rect 6636 32612 6692 32668
rect 6692 32612 6696 32668
rect 6632 32608 6696 32612
rect 6712 32668 6776 32672
rect 6712 32612 6716 32668
rect 6716 32612 6772 32668
rect 6772 32612 6776 32668
rect 6712 32608 6776 32612
rect 6792 32668 6856 32672
rect 6792 32612 6796 32668
rect 6796 32612 6852 32668
rect 6852 32612 6856 32668
rect 6792 32608 6856 32612
rect 14441 32668 14505 32672
rect 14441 32612 14445 32668
rect 14445 32612 14501 32668
rect 14501 32612 14505 32668
rect 14441 32608 14505 32612
rect 14521 32668 14585 32672
rect 14521 32612 14525 32668
rect 14525 32612 14581 32668
rect 14581 32612 14585 32668
rect 14521 32608 14585 32612
rect 14601 32668 14665 32672
rect 14601 32612 14605 32668
rect 14605 32612 14661 32668
rect 14661 32612 14665 32668
rect 14601 32608 14665 32612
rect 14681 32668 14745 32672
rect 14681 32612 14685 32668
rect 14685 32612 14741 32668
rect 14741 32612 14745 32668
rect 14681 32608 14745 32612
rect 22330 32668 22394 32672
rect 22330 32612 22334 32668
rect 22334 32612 22390 32668
rect 22390 32612 22394 32668
rect 22330 32608 22394 32612
rect 22410 32668 22474 32672
rect 22410 32612 22414 32668
rect 22414 32612 22470 32668
rect 22470 32612 22474 32668
rect 22410 32608 22474 32612
rect 22490 32668 22554 32672
rect 22490 32612 22494 32668
rect 22494 32612 22550 32668
rect 22550 32612 22554 32668
rect 22490 32608 22554 32612
rect 22570 32668 22634 32672
rect 22570 32612 22574 32668
rect 22574 32612 22630 32668
rect 22630 32612 22634 32668
rect 22570 32608 22634 32612
rect 30219 32668 30283 32672
rect 30219 32612 30223 32668
rect 30223 32612 30279 32668
rect 30279 32612 30283 32668
rect 30219 32608 30283 32612
rect 30299 32668 30363 32672
rect 30299 32612 30303 32668
rect 30303 32612 30359 32668
rect 30359 32612 30363 32668
rect 30299 32608 30363 32612
rect 30379 32668 30443 32672
rect 30379 32612 30383 32668
rect 30383 32612 30439 32668
rect 30439 32612 30443 32668
rect 30379 32608 30443 32612
rect 30459 32668 30523 32672
rect 30459 32612 30463 32668
rect 30463 32612 30519 32668
rect 30519 32612 30523 32668
rect 30459 32608 30523 32612
rect 7212 32124 7276 32128
rect 7212 32068 7216 32124
rect 7216 32068 7272 32124
rect 7272 32068 7276 32124
rect 7212 32064 7276 32068
rect 7292 32124 7356 32128
rect 7292 32068 7296 32124
rect 7296 32068 7352 32124
rect 7352 32068 7356 32124
rect 7292 32064 7356 32068
rect 7372 32124 7436 32128
rect 7372 32068 7376 32124
rect 7376 32068 7432 32124
rect 7432 32068 7436 32124
rect 7372 32064 7436 32068
rect 7452 32124 7516 32128
rect 7452 32068 7456 32124
rect 7456 32068 7512 32124
rect 7512 32068 7516 32124
rect 7452 32064 7516 32068
rect 15101 32124 15165 32128
rect 15101 32068 15105 32124
rect 15105 32068 15161 32124
rect 15161 32068 15165 32124
rect 15101 32064 15165 32068
rect 15181 32124 15245 32128
rect 15181 32068 15185 32124
rect 15185 32068 15241 32124
rect 15241 32068 15245 32124
rect 15181 32064 15245 32068
rect 15261 32124 15325 32128
rect 15261 32068 15265 32124
rect 15265 32068 15321 32124
rect 15321 32068 15325 32124
rect 15261 32064 15325 32068
rect 15341 32124 15405 32128
rect 15341 32068 15345 32124
rect 15345 32068 15401 32124
rect 15401 32068 15405 32124
rect 15341 32064 15405 32068
rect 22990 32124 23054 32128
rect 22990 32068 22994 32124
rect 22994 32068 23050 32124
rect 23050 32068 23054 32124
rect 22990 32064 23054 32068
rect 23070 32124 23134 32128
rect 23070 32068 23074 32124
rect 23074 32068 23130 32124
rect 23130 32068 23134 32124
rect 23070 32064 23134 32068
rect 23150 32124 23214 32128
rect 23150 32068 23154 32124
rect 23154 32068 23210 32124
rect 23210 32068 23214 32124
rect 23150 32064 23214 32068
rect 23230 32124 23294 32128
rect 23230 32068 23234 32124
rect 23234 32068 23290 32124
rect 23290 32068 23294 32124
rect 23230 32064 23294 32068
rect 30879 32124 30943 32128
rect 30879 32068 30883 32124
rect 30883 32068 30939 32124
rect 30939 32068 30943 32124
rect 30879 32064 30943 32068
rect 30959 32124 31023 32128
rect 30959 32068 30963 32124
rect 30963 32068 31019 32124
rect 31019 32068 31023 32124
rect 30959 32064 31023 32068
rect 31039 32124 31103 32128
rect 31039 32068 31043 32124
rect 31043 32068 31099 32124
rect 31099 32068 31103 32124
rect 31039 32064 31103 32068
rect 31119 32124 31183 32128
rect 31119 32068 31123 32124
rect 31123 32068 31179 32124
rect 31179 32068 31183 32124
rect 31119 32064 31183 32068
rect 6552 31580 6616 31584
rect 6552 31524 6556 31580
rect 6556 31524 6612 31580
rect 6612 31524 6616 31580
rect 6552 31520 6616 31524
rect 6632 31580 6696 31584
rect 6632 31524 6636 31580
rect 6636 31524 6692 31580
rect 6692 31524 6696 31580
rect 6632 31520 6696 31524
rect 6712 31580 6776 31584
rect 6712 31524 6716 31580
rect 6716 31524 6772 31580
rect 6772 31524 6776 31580
rect 6712 31520 6776 31524
rect 6792 31580 6856 31584
rect 6792 31524 6796 31580
rect 6796 31524 6852 31580
rect 6852 31524 6856 31580
rect 6792 31520 6856 31524
rect 14441 31580 14505 31584
rect 14441 31524 14445 31580
rect 14445 31524 14501 31580
rect 14501 31524 14505 31580
rect 14441 31520 14505 31524
rect 14521 31580 14585 31584
rect 14521 31524 14525 31580
rect 14525 31524 14581 31580
rect 14581 31524 14585 31580
rect 14521 31520 14585 31524
rect 14601 31580 14665 31584
rect 14601 31524 14605 31580
rect 14605 31524 14661 31580
rect 14661 31524 14665 31580
rect 14601 31520 14665 31524
rect 14681 31580 14745 31584
rect 14681 31524 14685 31580
rect 14685 31524 14741 31580
rect 14741 31524 14745 31580
rect 14681 31520 14745 31524
rect 22330 31580 22394 31584
rect 22330 31524 22334 31580
rect 22334 31524 22390 31580
rect 22390 31524 22394 31580
rect 22330 31520 22394 31524
rect 22410 31580 22474 31584
rect 22410 31524 22414 31580
rect 22414 31524 22470 31580
rect 22470 31524 22474 31580
rect 22410 31520 22474 31524
rect 22490 31580 22554 31584
rect 22490 31524 22494 31580
rect 22494 31524 22550 31580
rect 22550 31524 22554 31580
rect 22490 31520 22554 31524
rect 22570 31580 22634 31584
rect 22570 31524 22574 31580
rect 22574 31524 22630 31580
rect 22630 31524 22634 31580
rect 22570 31520 22634 31524
rect 30219 31580 30283 31584
rect 30219 31524 30223 31580
rect 30223 31524 30279 31580
rect 30279 31524 30283 31580
rect 30219 31520 30283 31524
rect 30299 31580 30363 31584
rect 30299 31524 30303 31580
rect 30303 31524 30359 31580
rect 30359 31524 30363 31580
rect 30299 31520 30363 31524
rect 30379 31580 30443 31584
rect 30379 31524 30383 31580
rect 30383 31524 30439 31580
rect 30439 31524 30443 31580
rect 30379 31520 30443 31524
rect 30459 31580 30523 31584
rect 30459 31524 30463 31580
rect 30463 31524 30519 31580
rect 30519 31524 30523 31580
rect 30459 31520 30523 31524
rect 7212 31036 7276 31040
rect 7212 30980 7216 31036
rect 7216 30980 7272 31036
rect 7272 30980 7276 31036
rect 7212 30976 7276 30980
rect 7292 31036 7356 31040
rect 7292 30980 7296 31036
rect 7296 30980 7352 31036
rect 7352 30980 7356 31036
rect 7292 30976 7356 30980
rect 7372 31036 7436 31040
rect 7372 30980 7376 31036
rect 7376 30980 7432 31036
rect 7432 30980 7436 31036
rect 7372 30976 7436 30980
rect 7452 31036 7516 31040
rect 7452 30980 7456 31036
rect 7456 30980 7512 31036
rect 7512 30980 7516 31036
rect 7452 30976 7516 30980
rect 15101 31036 15165 31040
rect 15101 30980 15105 31036
rect 15105 30980 15161 31036
rect 15161 30980 15165 31036
rect 15101 30976 15165 30980
rect 15181 31036 15245 31040
rect 15181 30980 15185 31036
rect 15185 30980 15241 31036
rect 15241 30980 15245 31036
rect 15181 30976 15245 30980
rect 15261 31036 15325 31040
rect 15261 30980 15265 31036
rect 15265 30980 15321 31036
rect 15321 30980 15325 31036
rect 15261 30976 15325 30980
rect 15341 31036 15405 31040
rect 15341 30980 15345 31036
rect 15345 30980 15401 31036
rect 15401 30980 15405 31036
rect 15341 30976 15405 30980
rect 22990 31036 23054 31040
rect 22990 30980 22994 31036
rect 22994 30980 23050 31036
rect 23050 30980 23054 31036
rect 22990 30976 23054 30980
rect 23070 31036 23134 31040
rect 23070 30980 23074 31036
rect 23074 30980 23130 31036
rect 23130 30980 23134 31036
rect 23070 30976 23134 30980
rect 23150 31036 23214 31040
rect 23150 30980 23154 31036
rect 23154 30980 23210 31036
rect 23210 30980 23214 31036
rect 23150 30976 23214 30980
rect 23230 31036 23294 31040
rect 23230 30980 23234 31036
rect 23234 30980 23290 31036
rect 23290 30980 23294 31036
rect 23230 30976 23294 30980
rect 30879 31036 30943 31040
rect 30879 30980 30883 31036
rect 30883 30980 30939 31036
rect 30939 30980 30943 31036
rect 30879 30976 30943 30980
rect 30959 31036 31023 31040
rect 30959 30980 30963 31036
rect 30963 30980 31019 31036
rect 31019 30980 31023 31036
rect 30959 30976 31023 30980
rect 31039 31036 31103 31040
rect 31039 30980 31043 31036
rect 31043 30980 31099 31036
rect 31099 30980 31103 31036
rect 31039 30976 31103 30980
rect 31119 31036 31183 31040
rect 31119 30980 31123 31036
rect 31123 30980 31179 31036
rect 31179 30980 31183 31036
rect 31119 30976 31183 30980
rect 6552 30492 6616 30496
rect 6552 30436 6556 30492
rect 6556 30436 6612 30492
rect 6612 30436 6616 30492
rect 6552 30432 6616 30436
rect 6632 30492 6696 30496
rect 6632 30436 6636 30492
rect 6636 30436 6692 30492
rect 6692 30436 6696 30492
rect 6632 30432 6696 30436
rect 6712 30492 6776 30496
rect 6712 30436 6716 30492
rect 6716 30436 6772 30492
rect 6772 30436 6776 30492
rect 6712 30432 6776 30436
rect 6792 30492 6856 30496
rect 6792 30436 6796 30492
rect 6796 30436 6852 30492
rect 6852 30436 6856 30492
rect 6792 30432 6856 30436
rect 14441 30492 14505 30496
rect 14441 30436 14445 30492
rect 14445 30436 14501 30492
rect 14501 30436 14505 30492
rect 14441 30432 14505 30436
rect 14521 30492 14585 30496
rect 14521 30436 14525 30492
rect 14525 30436 14581 30492
rect 14581 30436 14585 30492
rect 14521 30432 14585 30436
rect 14601 30492 14665 30496
rect 14601 30436 14605 30492
rect 14605 30436 14661 30492
rect 14661 30436 14665 30492
rect 14601 30432 14665 30436
rect 14681 30492 14745 30496
rect 14681 30436 14685 30492
rect 14685 30436 14741 30492
rect 14741 30436 14745 30492
rect 14681 30432 14745 30436
rect 22330 30492 22394 30496
rect 22330 30436 22334 30492
rect 22334 30436 22390 30492
rect 22390 30436 22394 30492
rect 22330 30432 22394 30436
rect 22410 30492 22474 30496
rect 22410 30436 22414 30492
rect 22414 30436 22470 30492
rect 22470 30436 22474 30492
rect 22410 30432 22474 30436
rect 22490 30492 22554 30496
rect 22490 30436 22494 30492
rect 22494 30436 22550 30492
rect 22550 30436 22554 30492
rect 22490 30432 22554 30436
rect 22570 30492 22634 30496
rect 22570 30436 22574 30492
rect 22574 30436 22630 30492
rect 22630 30436 22634 30492
rect 22570 30432 22634 30436
rect 30219 30492 30283 30496
rect 30219 30436 30223 30492
rect 30223 30436 30279 30492
rect 30279 30436 30283 30492
rect 30219 30432 30283 30436
rect 30299 30492 30363 30496
rect 30299 30436 30303 30492
rect 30303 30436 30359 30492
rect 30359 30436 30363 30492
rect 30299 30432 30363 30436
rect 30379 30492 30443 30496
rect 30379 30436 30383 30492
rect 30383 30436 30439 30492
rect 30439 30436 30443 30492
rect 30379 30432 30443 30436
rect 30459 30492 30523 30496
rect 30459 30436 30463 30492
rect 30463 30436 30519 30492
rect 30519 30436 30523 30492
rect 30459 30432 30523 30436
rect 7212 29948 7276 29952
rect 7212 29892 7216 29948
rect 7216 29892 7272 29948
rect 7272 29892 7276 29948
rect 7212 29888 7276 29892
rect 7292 29948 7356 29952
rect 7292 29892 7296 29948
rect 7296 29892 7352 29948
rect 7352 29892 7356 29948
rect 7292 29888 7356 29892
rect 7372 29948 7436 29952
rect 7372 29892 7376 29948
rect 7376 29892 7432 29948
rect 7432 29892 7436 29948
rect 7372 29888 7436 29892
rect 7452 29948 7516 29952
rect 7452 29892 7456 29948
rect 7456 29892 7512 29948
rect 7512 29892 7516 29948
rect 7452 29888 7516 29892
rect 15101 29948 15165 29952
rect 15101 29892 15105 29948
rect 15105 29892 15161 29948
rect 15161 29892 15165 29948
rect 15101 29888 15165 29892
rect 15181 29948 15245 29952
rect 15181 29892 15185 29948
rect 15185 29892 15241 29948
rect 15241 29892 15245 29948
rect 15181 29888 15245 29892
rect 15261 29948 15325 29952
rect 15261 29892 15265 29948
rect 15265 29892 15321 29948
rect 15321 29892 15325 29948
rect 15261 29888 15325 29892
rect 15341 29948 15405 29952
rect 15341 29892 15345 29948
rect 15345 29892 15401 29948
rect 15401 29892 15405 29948
rect 15341 29888 15405 29892
rect 22990 29948 23054 29952
rect 22990 29892 22994 29948
rect 22994 29892 23050 29948
rect 23050 29892 23054 29948
rect 22990 29888 23054 29892
rect 23070 29948 23134 29952
rect 23070 29892 23074 29948
rect 23074 29892 23130 29948
rect 23130 29892 23134 29948
rect 23070 29888 23134 29892
rect 23150 29948 23214 29952
rect 23150 29892 23154 29948
rect 23154 29892 23210 29948
rect 23210 29892 23214 29948
rect 23150 29888 23214 29892
rect 23230 29948 23294 29952
rect 23230 29892 23234 29948
rect 23234 29892 23290 29948
rect 23290 29892 23294 29948
rect 23230 29888 23294 29892
rect 30879 29948 30943 29952
rect 30879 29892 30883 29948
rect 30883 29892 30939 29948
rect 30939 29892 30943 29948
rect 30879 29888 30943 29892
rect 30959 29948 31023 29952
rect 30959 29892 30963 29948
rect 30963 29892 31019 29948
rect 31019 29892 31023 29948
rect 30959 29888 31023 29892
rect 31039 29948 31103 29952
rect 31039 29892 31043 29948
rect 31043 29892 31099 29948
rect 31099 29892 31103 29948
rect 31039 29888 31103 29892
rect 31119 29948 31183 29952
rect 31119 29892 31123 29948
rect 31123 29892 31179 29948
rect 31179 29892 31183 29948
rect 31119 29888 31183 29892
rect 6552 29404 6616 29408
rect 6552 29348 6556 29404
rect 6556 29348 6612 29404
rect 6612 29348 6616 29404
rect 6552 29344 6616 29348
rect 6632 29404 6696 29408
rect 6632 29348 6636 29404
rect 6636 29348 6692 29404
rect 6692 29348 6696 29404
rect 6632 29344 6696 29348
rect 6712 29404 6776 29408
rect 6712 29348 6716 29404
rect 6716 29348 6772 29404
rect 6772 29348 6776 29404
rect 6712 29344 6776 29348
rect 6792 29404 6856 29408
rect 6792 29348 6796 29404
rect 6796 29348 6852 29404
rect 6852 29348 6856 29404
rect 6792 29344 6856 29348
rect 14441 29404 14505 29408
rect 14441 29348 14445 29404
rect 14445 29348 14501 29404
rect 14501 29348 14505 29404
rect 14441 29344 14505 29348
rect 14521 29404 14585 29408
rect 14521 29348 14525 29404
rect 14525 29348 14581 29404
rect 14581 29348 14585 29404
rect 14521 29344 14585 29348
rect 14601 29404 14665 29408
rect 14601 29348 14605 29404
rect 14605 29348 14661 29404
rect 14661 29348 14665 29404
rect 14601 29344 14665 29348
rect 14681 29404 14745 29408
rect 14681 29348 14685 29404
rect 14685 29348 14741 29404
rect 14741 29348 14745 29404
rect 14681 29344 14745 29348
rect 22330 29404 22394 29408
rect 22330 29348 22334 29404
rect 22334 29348 22390 29404
rect 22390 29348 22394 29404
rect 22330 29344 22394 29348
rect 22410 29404 22474 29408
rect 22410 29348 22414 29404
rect 22414 29348 22470 29404
rect 22470 29348 22474 29404
rect 22410 29344 22474 29348
rect 22490 29404 22554 29408
rect 22490 29348 22494 29404
rect 22494 29348 22550 29404
rect 22550 29348 22554 29404
rect 22490 29344 22554 29348
rect 22570 29404 22634 29408
rect 22570 29348 22574 29404
rect 22574 29348 22630 29404
rect 22630 29348 22634 29404
rect 22570 29344 22634 29348
rect 30219 29404 30283 29408
rect 30219 29348 30223 29404
rect 30223 29348 30279 29404
rect 30279 29348 30283 29404
rect 30219 29344 30283 29348
rect 30299 29404 30363 29408
rect 30299 29348 30303 29404
rect 30303 29348 30359 29404
rect 30359 29348 30363 29404
rect 30299 29344 30363 29348
rect 30379 29404 30443 29408
rect 30379 29348 30383 29404
rect 30383 29348 30439 29404
rect 30439 29348 30443 29404
rect 30379 29344 30443 29348
rect 30459 29404 30523 29408
rect 30459 29348 30463 29404
rect 30463 29348 30519 29404
rect 30519 29348 30523 29404
rect 30459 29344 30523 29348
rect 27844 29004 27908 29068
rect 7212 28860 7276 28864
rect 7212 28804 7216 28860
rect 7216 28804 7272 28860
rect 7272 28804 7276 28860
rect 7212 28800 7276 28804
rect 7292 28860 7356 28864
rect 7292 28804 7296 28860
rect 7296 28804 7352 28860
rect 7352 28804 7356 28860
rect 7292 28800 7356 28804
rect 7372 28860 7436 28864
rect 7372 28804 7376 28860
rect 7376 28804 7432 28860
rect 7432 28804 7436 28860
rect 7372 28800 7436 28804
rect 7452 28860 7516 28864
rect 7452 28804 7456 28860
rect 7456 28804 7512 28860
rect 7512 28804 7516 28860
rect 7452 28800 7516 28804
rect 15101 28860 15165 28864
rect 15101 28804 15105 28860
rect 15105 28804 15161 28860
rect 15161 28804 15165 28860
rect 15101 28800 15165 28804
rect 15181 28860 15245 28864
rect 15181 28804 15185 28860
rect 15185 28804 15241 28860
rect 15241 28804 15245 28860
rect 15181 28800 15245 28804
rect 15261 28860 15325 28864
rect 15261 28804 15265 28860
rect 15265 28804 15321 28860
rect 15321 28804 15325 28860
rect 15261 28800 15325 28804
rect 15341 28860 15405 28864
rect 15341 28804 15345 28860
rect 15345 28804 15401 28860
rect 15401 28804 15405 28860
rect 15341 28800 15405 28804
rect 22990 28860 23054 28864
rect 22990 28804 22994 28860
rect 22994 28804 23050 28860
rect 23050 28804 23054 28860
rect 22990 28800 23054 28804
rect 23070 28860 23134 28864
rect 23070 28804 23074 28860
rect 23074 28804 23130 28860
rect 23130 28804 23134 28860
rect 23070 28800 23134 28804
rect 23150 28860 23214 28864
rect 23150 28804 23154 28860
rect 23154 28804 23210 28860
rect 23210 28804 23214 28860
rect 23150 28800 23214 28804
rect 23230 28860 23294 28864
rect 23230 28804 23234 28860
rect 23234 28804 23290 28860
rect 23290 28804 23294 28860
rect 23230 28800 23294 28804
rect 30879 28860 30943 28864
rect 30879 28804 30883 28860
rect 30883 28804 30939 28860
rect 30939 28804 30943 28860
rect 30879 28800 30943 28804
rect 30959 28860 31023 28864
rect 30959 28804 30963 28860
rect 30963 28804 31019 28860
rect 31019 28804 31023 28860
rect 30959 28800 31023 28804
rect 31039 28860 31103 28864
rect 31039 28804 31043 28860
rect 31043 28804 31099 28860
rect 31099 28804 31103 28860
rect 31039 28800 31103 28804
rect 31119 28860 31183 28864
rect 31119 28804 31123 28860
rect 31123 28804 31179 28860
rect 31179 28804 31183 28860
rect 31119 28800 31183 28804
rect 6552 28316 6616 28320
rect 6552 28260 6556 28316
rect 6556 28260 6612 28316
rect 6612 28260 6616 28316
rect 6552 28256 6616 28260
rect 6632 28316 6696 28320
rect 6632 28260 6636 28316
rect 6636 28260 6692 28316
rect 6692 28260 6696 28316
rect 6632 28256 6696 28260
rect 6712 28316 6776 28320
rect 6712 28260 6716 28316
rect 6716 28260 6772 28316
rect 6772 28260 6776 28316
rect 6712 28256 6776 28260
rect 6792 28316 6856 28320
rect 6792 28260 6796 28316
rect 6796 28260 6852 28316
rect 6852 28260 6856 28316
rect 6792 28256 6856 28260
rect 14441 28316 14505 28320
rect 14441 28260 14445 28316
rect 14445 28260 14501 28316
rect 14501 28260 14505 28316
rect 14441 28256 14505 28260
rect 14521 28316 14585 28320
rect 14521 28260 14525 28316
rect 14525 28260 14581 28316
rect 14581 28260 14585 28316
rect 14521 28256 14585 28260
rect 14601 28316 14665 28320
rect 14601 28260 14605 28316
rect 14605 28260 14661 28316
rect 14661 28260 14665 28316
rect 14601 28256 14665 28260
rect 14681 28316 14745 28320
rect 14681 28260 14685 28316
rect 14685 28260 14741 28316
rect 14741 28260 14745 28316
rect 14681 28256 14745 28260
rect 22330 28316 22394 28320
rect 22330 28260 22334 28316
rect 22334 28260 22390 28316
rect 22390 28260 22394 28316
rect 22330 28256 22394 28260
rect 22410 28316 22474 28320
rect 22410 28260 22414 28316
rect 22414 28260 22470 28316
rect 22470 28260 22474 28316
rect 22410 28256 22474 28260
rect 22490 28316 22554 28320
rect 22490 28260 22494 28316
rect 22494 28260 22550 28316
rect 22550 28260 22554 28316
rect 22490 28256 22554 28260
rect 22570 28316 22634 28320
rect 22570 28260 22574 28316
rect 22574 28260 22630 28316
rect 22630 28260 22634 28316
rect 22570 28256 22634 28260
rect 30219 28316 30283 28320
rect 30219 28260 30223 28316
rect 30223 28260 30279 28316
rect 30279 28260 30283 28316
rect 30219 28256 30283 28260
rect 30299 28316 30363 28320
rect 30299 28260 30303 28316
rect 30303 28260 30359 28316
rect 30359 28260 30363 28316
rect 30299 28256 30363 28260
rect 30379 28316 30443 28320
rect 30379 28260 30383 28316
rect 30383 28260 30439 28316
rect 30439 28260 30443 28316
rect 30379 28256 30443 28260
rect 30459 28316 30523 28320
rect 30459 28260 30463 28316
rect 30463 28260 30519 28316
rect 30519 28260 30523 28316
rect 30459 28256 30523 28260
rect 7212 27772 7276 27776
rect 7212 27716 7216 27772
rect 7216 27716 7272 27772
rect 7272 27716 7276 27772
rect 7212 27712 7276 27716
rect 7292 27772 7356 27776
rect 7292 27716 7296 27772
rect 7296 27716 7352 27772
rect 7352 27716 7356 27772
rect 7292 27712 7356 27716
rect 7372 27772 7436 27776
rect 7372 27716 7376 27772
rect 7376 27716 7432 27772
rect 7432 27716 7436 27772
rect 7372 27712 7436 27716
rect 7452 27772 7516 27776
rect 7452 27716 7456 27772
rect 7456 27716 7512 27772
rect 7512 27716 7516 27772
rect 7452 27712 7516 27716
rect 15101 27772 15165 27776
rect 15101 27716 15105 27772
rect 15105 27716 15161 27772
rect 15161 27716 15165 27772
rect 15101 27712 15165 27716
rect 15181 27772 15245 27776
rect 15181 27716 15185 27772
rect 15185 27716 15241 27772
rect 15241 27716 15245 27772
rect 15181 27712 15245 27716
rect 15261 27772 15325 27776
rect 15261 27716 15265 27772
rect 15265 27716 15321 27772
rect 15321 27716 15325 27772
rect 15261 27712 15325 27716
rect 15341 27772 15405 27776
rect 15341 27716 15345 27772
rect 15345 27716 15401 27772
rect 15401 27716 15405 27772
rect 15341 27712 15405 27716
rect 22990 27772 23054 27776
rect 22990 27716 22994 27772
rect 22994 27716 23050 27772
rect 23050 27716 23054 27772
rect 22990 27712 23054 27716
rect 23070 27772 23134 27776
rect 23070 27716 23074 27772
rect 23074 27716 23130 27772
rect 23130 27716 23134 27772
rect 23070 27712 23134 27716
rect 23150 27772 23214 27776
rect 23150 27716 23154 27772
rect 23154 27716 23210 27772
rect 23210 27716 23214 27772
rect 23150 27712 23214 27716
rect 23230 27772 23294 27776
rect 23230 27716 23234 27772
rect 23234 27716 23290 27772
rect 23290 27716 23294 27772
rect 23230 27712 23294 27716
rect 30879 27772 30943 27776
rect 30879 27716 30883 27772
rect 30883 27716 30939 27772
rect 30939 27716 30943 27772
rect 30879 27712 30943 27716
rect 30959 27772 31023 27776
rect 30959 27716 30963 27772
rect 30963 27716 31019 27772
rect 31019 27716 31023 27772
rect 30959 27712 31023 27716
rect 31039 27772 31103 27776
rect 31039 27716 31043 27772
rect 31043 27716 31099 27772
rect 31099 27716 31103 27772
rect 31039 27712 31103 27716
rect 31119 27772 31183 27776
rect 31119 27716 31123 27772
rect 31123 27716 31179 27772
rect 31179 27716 31183 27772
rect 31119 27712 31183 27716
rect 6552 27228 6616 27232
rect 6552 27172 6556 27228
rect 6556 27172 6612 27228
rect 6612 27172 6616 27228
rect 6552 27168 6616 27172
rect 6632 27228 6696 27232
rect 6632 27172 6636 27228
rect 6636 27172 6692 27228
rect 6692 27172 6696 27228
rect 6632 27168 6696 27172
rect 6712 27228 6776 27232
rect 6712 27172 6716 27228
rect 6716 27172 6772 27228
rect 6772 27172 6776 27228
rect 6712 27168 6776 27172
rect 6792 27228 6856 27232
rect 6792 27172 6796 27228
rect 6796 27172 6852 27228
rect 6852 27172 6856 27228
rect 6792 27168 6856 27172
rect 14441 27228 14505 27232
rect 14441 27172 14445 27228
rect 14445 27172 14501 27228
rect 14501 27172 14505 27228
rect 14441 27168 14505 27172
rect 14521 27228 14585 27232
rect 14521 27172 14525 27228
rect 14525 27172 14581 27228
rect 14581 27172 14585 27228
rect 14521 27168 14585 27172
rect 14601 27228 14665 27232
rect 14601 27172 14605 27228
rect 14605 27172 14661 27228
rect 14661 27172 14665 27228
rect 14601 27168 14665 27172
rect 14681 27228 14745 27232
rect 14681 27172 14685 27228
rect 14685 27172 14741 27228
rect 14741 27172 14745 27228
rect 14681 27168 14745 27172
rect 22330 27228 22394 27232
rect 22330 27172 22334 27228
rect 22334 27172 22390 27228
rect 22390 27172 22394 27228
rect 22330 27168 22394 27172
rect 22410 27228 22474 27232
rect 22410 27172 22414 27228
rect 22414 27172 22470 27228
rect 22470 27172 22474 27228
rect 22410 27168 22474 27172
rect 22490 27228 22554 27232
rect 22490 27172 22494 27228
rect 22494 27172 22550 27228
rect 22550 27172 22554 27228
rect 22490 27168 22554 27172
rect 22570 27228 22634 27232
rect 22570 27172 22574 27228
rect 22574 27172 22630 27228
rect 22630 27172 22634 27228
rect 22570 27168 22634 27172
rect 30219 27228 30283 27232
rect 30219 27172 30223 27228
rect 30223 27172 30279 27228
rect 30279 27172 30283 27228
rect 30219 27168 30283 27172
rect 30299 27228 30363 27232
rect 30299 27172 30303 27228
rect 30303 27172 30359 27228
rect 30359 27172 30363 27228
rect 30299 27168 30363 27172
rect 30379 27228 30443 27232
rect 30379 27172 30383 27228
rect 30383 27172 30439 27228
rect 30439 27172 30443 27228
rect 30379 27168 30443 27172
rect 30459 27228 30523 27232
rect 30459 27172 30463 27228
rect 30463 27172 30519 27228
rect 30519 27172 30523 27228
rect 30459 27168 30523 27172
rect 7212 26684 7276 26688
rect 7212 26628 7216 26684
rect 7216 26628 7272 26684
rect 7272 26628 7276 26684
rect 7212 26624 7276 26628
rect 7292 26684 7356 26688
rect 7292 26628 7296 26684
rect 7296 26628 7352 26684
rect 7352 26628 7356 26684
rect 7292 26624 7356 26628
rect 7372 26684 7436 26688
rect 7372 26628 7376 26684
rect 7376 26628 7432 26684
rect 7432 26628 7436 26684
rect 7372 26624 7436 26628
rect 7452 26684 7516 26688
rect 7452 26628 7456 26684
rect 7456 26628 7512 26684
rect 7512 26628 7516 26684
rect 7452 26624 7516 26628
rect 15101 26684 15165 26688
rect 15101 26628 15105 26684
rect 15105 26628 15161 26684
rect 15161 26628 15165 26684
rect 15101 26624 15165 26628
rect 15181 26684 15245 26688
rect 15181 26628 15185 26684
rect 15185 26628 15241 26684
rect 15241 26628 15245 26684
rect 15181 26624 15245 26628
rect 15261 26684 15325 26688
rect 15261 26628 15265 26684
rect 15265 26628 15321 26684
rect 15321 26628 15325 26684
rect 15261 26624 15325 26628
rect 15341 26684 15405 26688
rect 15341 26628 15345 26684
rect 15345 26628 15401 26684
rect 15401 26628 15405 26684
rect 15341 26624 15405 26628
rect 22990 26684 23054 26688
rect 22990 26628 22994 26684
rect 22994 26628 23050 26684
rect 23050 26628 23054 26684
rect 22990 26624 23054 26628
rect 23070 26684 23134 26688
rect 23070 26628 23074 26684
rect 23074 26628 23130 26684
rect 23130 26628 23134 26684
rect 23070 26624 23134 26628
rect 23150 26684 23214 26688
rect 23150 26628 23154 26684
rect 23154 26628 23210 26684
rect 23210 26628 23214 26684
rect 23150 26624 23214 26628
rect 23230 26684 23294 26688
rect 23230 26628 23234 26684
rect 23234 26628 23290 26684
rect 23290 26628 23294 26684
rect 23230 26624 23294 26628
rect 30879 26684 30943 26688
rect 30879 26628 30883 26684
rect 30883 26628 30939 26684
rect 30939 26628 30943 26684
rect 30879 26624 30943 26628
rect 30959 26684 31023 26688
rect 30959 26628 30963 26684
rect 30963 26628 31019 26684
rect 31019 26628 31023 26684
rect 30959 26624 31023 26628
rect 31039 26684 31103 26688
rect 31039 26628 31043 26684
rect 31043 26628 31099 26684
rect 31099 26628 31103 26684
rect 31039 26624 31103 26628
rect 31119 26684 31183 26688
rect 31119 26628 31123 26684
rect 31123 26628 31179 26684
rect 31179 26628 31183 26684
rect 31119 26624 31183 26628
rect 17356 26344 17420 26348
rect 17356 26288 17406 26344
rect 17406 26288 17420 26344
rect 17356 26284 17420 26288
rect 6552 26140 6616 26144
rect 6552 26084 6556 26140
rect 6556 26084 6612 26140
rect 6612 26084 6616 26140
rect 6552 26080 6616 26084
rect 6632 26140 6696 26144
rect 6632 26084 6636 26140
rect 6636 26084 6692 26140
rect 6692 26084 6696 26140
rect 6632 26080 6696 26084
rect 6712 26140 6776 26144
rect 6712 26084 6716 26140
rect 6716 26084 6772 26140
rect 6772 26084 6776 26140
rect 6712 26080 6776 26084
rect 6792 26140 6856 26144
rect 6792 26084 6796 26140
rect 6796 26084 6852 26140
rect 6852 26084 6856 26140
rect 6792 26080 6856 26084
rect 14441 26140 14505 26144
rect 14441 26084 14445 26140
rect 14445 26084 14501 26140
rect 14501 26084 14505 26140
rect 14441 26080 14505 26084
rect 14521 26140 14585 26144
rect 14521 26084 14525 26140
rect 14525 26084 14581 26140
rect 14581 26084 14585 26140
rect 14521 26080 14585 26084
rect 14601 26140 14665 26144
rect 14601 26084 14605 26140
rect 14605 26084 14661 26140
rect 14661 26084 14665 26140
rect 14601 26080 14665 26084
rect 14681 26140 14745 26144
rect 14681 26084 14685 26140
rect 14685 26084 14741 26140
rect 14741 26084 14745 26140
rect 14681 26080 14745 26084
rect 22330 26140 22394 26144
rect 22330 26084 22334 26140
rect 22334 26084 22390 26140
rect 22390 26084 22394 26140
rect 22330 26080 22394 26084
rect 22410 26140 22474 26144
rect 22410 26084 22414 26140
rect 22414 26084 22470 26140
rect 22470 26084 22474 26140
rect 22410 26080 22474 26084
rect 22490 26140 22554 26144
rect 22490 26084 22494 26140
rect 22494 26084 22550 26140
rect 22550 26084 22554 26140
rect 22490 26080 22554 26084
rect 22570 26140 22634 26144
rect 22570 26084 22574 26140
rect 22574 26084 22630 26140
rect 22630 26084 22634 26140
rect 22570 26080 22634 26084
rect 30219 26140 30283 26144
rect 30219 26084 30223 26140
rect 30223 26084 30279 26140
rect 30279 26084 30283 26140
rect 30219 26080 30283 26084
rect 30299 26140 30363 26144
rect 30299 26084 30303 26140
rect 30303 26084 30359 26140
rect 30359 26084 30363 26140
rect 30299 26080 30363 26084
rect 30379 26140 30443 26144
rect 30379 26084 30383 26140
rect 30383 26084 30439 26140
rect 30439 26084 30443 26140
rect 30379 26080 30443 26084
rect 30459 26140 30523 26144
rect 30459 26084 30463 26140
rect 30463 26084 30519 26140
rect 30519 26084 30523 26140
rect 30459 26080 30523 26084
rect 7212 25596 7276 25600
rect 7212 25540 7216 25596
rect 7216 25540 7272 25596
rect 7272 25540 7276 25596
rect 7212 25536 7276 25540
rect 7292 25596 7356 25600
rect 7292 25540 7296 25596
rect 7296 25540 7352 25596
rect 7352 25540 7356 25596
rect 7292 25536 7356 25540
rect 7372 25596 7436 25600
rect 7372 25540 7376 25596
rect 7376 25540 7432 25596
rect 7432 25540 7436 25596
rect 7372 25536 7436 25540
rect 7452 25596 7516 25600
rect 7452 25540 7456 25596
rect 7456 25540 7512 25596
rect 7512 25540 7516 25596
rect 7452 25536 7516 25540
rect 15101 25596 15165 25600
rect 15101 25540 15105 25596
rect 15105 25540 15161 25596
rect 15161 25540 15165 25596
rect 15101 25536 15165 25540
rect 15181 25596 15245 25600
rect 15181 25540 15185 25596
rect 15185 25540 15241 25596
rect 15241 25540 15245 25596
rect 15181 25536 15245 25540
rect 15261 25596 15325 25600
rect 15261 25540 15265 25596
rect 15265 25540 15321 25596
rect 15321 25540 15325 25596
rect 15261 25536 15325 25540
rect 15341 25596 15405 25600
rect 15341 25540 15345 25596
rect 15345 25540 15401 25596
rect 15401 25540 15405 25596
rect 15341 25536 15405 25540
rect 22990 25596 23054 25600
rect 22990 25540 22994 25596
rect 22994 25540 23050 25596
rect 23050 25540 23054 25596
rect 22990 25536 23054 25540
rect 23070 25596 23134 25600
rect 23070 25540 23074 25596
rect 23074 25540 23130 25596
rect 23130 25540 23134 25596
rect 23070 25536 23134 25540
rect 23150 25596 23214 25600
rect 23150 25540 23154 25596
rect 23154 25540 23210 25596
rect 23210 25540 23214 25596
rect 23150 25536 23214 25540
rect 23230 25596 23294 25600
rect 23230 25540 23234 25596
rect 23234 25540 23290 25596
rect 23290 25540 23294 25596
rect 23230 25536 23294 25540
rect 30879 25596 30943 25600
rect 30879 25540 30883 25596
rect 30883 25540 30939 25596
rect 30939 25540 30943 25596
rect 30879 25536 30943 25540
rect 30959 25596 31023 25600
rect 30959 25540 30963 25596
rect 30963 25540 31019 25596
rect 31019 25540 31023 25596
rect 30959 25536 31023 25540
rect 31039 25596 31103 25600
rect 31039 25540 31043 25596
rect 31043 25540 31099 25596
rect 31099 25540 31103 25596
rect 31039 25536 31103 25540
rect 31119 25596 31183 25600
rect 31119 25540 31123 25596
rect 31123 25540 31179 25596
rect 31179 25540 31183 25596
rect 31119 25536 31183 25540
rect 6552 25052 6616 25056
rect 6552 24996 6556 25052
rect 6556 24996 6612 25052
rect 6612 24996 6616 25052
rect 6552 24992 6616 24996
rect 6632 25052 6696 25056
rect 6632 24996 6636 25052
rect 6636 24996 6692 25052
rect 6692 24996 6696 25052
rect 6632 24992 6696 24996
rect 6712 25052 6776 25056
rect 6712 24996 6716 25052
rect 6716 24996 6772 25052
rect 6772 24996 6776 25052
rect 6712 24992 6776 24996
rect 6792 25052 6856 25056
rect 6792 24996 6796 25052
rect 6796 24996 6852 25052
rect 6852 24996 6856 25052
rect 6792 24992 6856 24996
rect 14441 25052 14505 25056
rect 14441 24996 14445 25052
rect 14445 24996 14501 25052
rect 14501 24996 14505 25052
rect 14441 24992 14505 24996
rect 14521 25052 14585 25056
rect 14521 24996 14525 25052
rect 14525 24996 14581 25052
rect 14581 24996 14585 25052
rect 14521 24992 14585 24996
rect 14601 25052 14665 25056
rect 14601 24996 14605 25052
rect 14605 24996 14661 25052
rect 14661 24996 14665 25052
rect 14601 24992 14665 24996
rect 14681 25052 14745 25056
rect 14681 24996 14685 25052
rect 14685 24996 14741 25052
rect 14741 24996 14745 25052
rect 14681 24992 14745 24996
rect 22330 25052 22394 25056
rect 22330 24996 22334 25052
rect 22334 24996 22390 25052
rect 22390 24996 22394 25052
rect 22330 24992 22394 24996
rect 22410 25052 22474 25056
rect 22410 24996 22414 25052
rect 22414 24996 22470 25052
rect 22470 24996 22474 25052
rect 22410 24992 22474 24996
rect 22490 25052 22554 25056
rect 22490 24996 22494 25052
rect 22494 24996 22550 25052
rect 22550 24996 22554 25052
rect 22490 24992 22554 24996
rect 22570 25052 22634 25056
rect 22570 24996 22574 25052
rect 22574 24996 22630 25052
rect 22630 24996 22634 25052
rect 22570 24992 22634 24996
rect 30219 25052 30283 25056
rect 30219 24996 30223 25052
rect 30223 24996 30279 25052
rect 30279 24996 30283 25052
rect 30219 24992 30283 24996
rect 30299 25052 30363 25056
rect 30299 24996 30303 25052
rect 30303 24996 30359 25052
rect 30359 24996 30363 25052
rect 30299 24992 30363 24996
rect 30379 25052 30443 25056
rect 30379 24996 30383 25052
rect 30383 24996 30439 25052
rect 30439 24996 30443 25052
rect 30379 24992 30443 24996
rect 30459 25052 30523 25056
rect 30459 24996 30463 25052
rect 30463 24996 30519 25052
rect 30519 24996 30523 25052
rect 30459 24992 30523 24996
rect 5580 24924 5644 24988
rect 7212 24508 7276 24512
rect 7212 24452 7216 24508
rect 7216 24452 7272 24508
rect 7272 24452 7276 24508
rect 7212 24448 7276 24452
rect 7292 24508 7356 24512
rect 7292 24452 7296 24508
rect 7296 24452 7352 24508
rect 7352 24452 7356 24508
rect 7292 24448 7356 24452
rect 7372 24508 7436 24512
rect 7372 24452 7376 24508
rect 7376 24452 7432 24508
rect 7432 24452 7436 24508
rect 7372 24448 7436 24452
rect 7452 24508 7516 24512
rect 7452 24452 7456 24508
rect 7456 24452 7512 24508
rect 7512 24452 7516 24508
rect 7452 24448 7516 24452
rect 15101 24508 15165 24512
rect 15101 24452 15105 24508
rect 15105 24452 15161 24508
rect 15161 24452 15165 24508
rect 15101 24448 15165 24452
rect 15181 24508 15245 24512
rect 15181 24452 15185 24508
rect 15185 24452 15241 24508
rect 15241 24452 15245 24508
rect 15181 24448 15245 24452
rect 15261 24508 15325 24512
rect 15261 24452 15265 24508
rect 15265 24452 15321 24508
rect 15321 24452 15325 24508
rect 15261 24448 15325 24452
rect 15341 24508 15405 24512
rect 15341 24452 15345 24508
rect 15345 24452 15401 24508
rect 15401 24452 15405 24508
rect 15341 24448 15405 24452
rect 22990 24508 23054 24512
rect 22990 24452 22994 24508
rect 22994 24452 23050 24508
rect 23050 24452 23054 24508
rect 22990 24448 23054 24452
rect 23070 24508 23134 24512
rect 23070 24452 23074 24508
rect 23074 24452 23130 24508
rect 23130 24452 23134 24508
rect 23070 24448 23134 24452
rect 23150 24508 23214 24512
rect 23150 24452 23154 24508
rect 23154 24452 23210 24508
rect 23210 24452 23214 24508
rect 23150 24448 23214 24452
rect 23230 24508 23294 24512
rect 23230 24452 23234 24508
rect 23234 24452 23290 24508
rect 23290 24452 23294 24508
rect 23230 24448 23294 24452
rect 30879 24508 30943 24512
rect 30879 24452 30883 24508
rect 30883 24452 30939 24508
rect 30939 24452 30943 24508
rect 30879 24448 30943 24452
rect 30959 24508 31023 24512
rect 30959 24452 30963 24508
rect 30963 24452 31019 24508
rect 31019 24452 31023 24508
rect 30959 24448 31023 24452
rect 31039 24508 31103 24512
rect 31039 24452 31043 24508
rect 31043 24452 31099 24508
rect 31099 24452 31103 24508
rect 31039 24448 31103 24452
rect 31119 24508 31183 24512
rect 31119 24452 31123 24508
rect 31123 24452 31179 24508
rect 31179 24452 31183 24508
rect 31119 24448 31183 24452
rect 26556 24032 26620 24036
rect 26556 23976 26606 24032
rect 26606 23976 26620 24032
rect 26556 23972 26620 23976
rect 6552 23964 6616 23968
rect 6552 23908 6556 23964
rect 6556 23908 6612 23964
rect 6612 23908 6616 23964
rect 6552 23904 6616 23908
rect 6632 23964 6696 23968
rect 6632 23908 6636 23964
rect 6636 23908 6692 23964
rect 6692 23908 6696 23964
rect 6632 23904 6696 23908
rect 6712 23964 6776 23968
rect 6712 23908 6716 23964
rect 6716 23908 6772 23964
rect 6772 23908 6776 23964
rect 6712 23904 6776 23908
rect 6792 23964 6856 23968
rect 6792 23908 6796 23964
rect 6796 23908 6852 23964
rect 6852 23908 6856 23964
rect 6792 23904 6856 23908
rect 14441 23964 14505 23968
rect 14441 23908 14445 23964
rect 14445 23908 14501 23964
rect 14501 23908 14505 23964
rect 14441 23904 14505 23908
rect 14521 23964 14585 23968
rect 14521 23908 14525 23964
rect 14525 23908 14581 23964
rect 14581 23908 14585 23964
rect 14521 23904 14585 23908
rect 14601 23964 14665 23968
rect 14601 23908 14605 23964
rect 14605 23908 14661 23964
rect 14661 23908 14665 23964
rect 14601 23904 14665 23908
rect 14681 23964 14745 23968
rect 14681 23908 14685 23964
rect 14685 23908 14741 23964
rect 14741 23908 14745 23964
rect 14681 23904 14745 23908
rect 22330 23964 22394 23968
rect 22330 23908 22334 23964
rect 22334 23908 22390 23964
rect 22390 23908 22394 23964
rect 22330 23904 22394 23908
rect 22410 23964 22474 23968
rect 22410 23908 22414 23964
rect 22414 23908 22470 23964
rect 22470 23908 22474 23964
rect 22410 23904 22474 23908
rect 22490 23964 22554 23968
rect 22490 23908 22494 23964
rect 22494 23908 22550 23964
rect 22550 23908 22554 23964
rect 22490 23904 22554 23908
rect 22570 23964 22634 23968
rect 22570 23908 22574 23964
rect 22574 23908 22630 23964
rect 22630 23908 22634 23964
rect 22570 23904 22634 23908
rect 30219 23964 30283 23968
rect 30219 23908 30223 23964
rect 30223 23908 30279 23964
rect 30279 23908 30283 23964
rect 30219 23904 30283 23908
rect 30299 23964 30363 23968
rect 30299 23908 30303 23964
rect 30303 23908 30359 23964
rect 30359 23908 30363 23964
rect 30299 23904 30363 23908
rect 30379 23964 30443 23968
rect 30379 23908 30383 23964
rect 30383 23908 30439 23964
rect 30439 23908 30443 23964
rect 30379 23904 30443 23908
rect 30459 23964 30523 23968
rect 30459 23908 30463 23964
rect 30463 23908 30519 23964
rect 30519 23908 30523 23964
rect 30459 23904 30523 23908
rect 15700 23700 15764 23764
rect 6132 23624 6196 23628
rect 6132 23568 6182 23624
rect 6182 23568 6196 23624
rect 6132 23564 6196 23568
rect 5764 23488 5828 23492
rect 5764 23432 5814 23488
rect 5814 23432 5828 23488
rect 5764 23428 5828 23432
rect 7212 23420 7276 23424
rect 7212 23364 7216 23420
rect 7216 23364 7272 23420
rect 7272 23364 7276 23420
rect 7212 23360 7276 23364
rect 7292 23420 7356 23424
rect 7292 23364 7296 23420
rect 7296 23364 7352 23420
rect 7352 23364 7356 23420
rect 7292 23360 7356 23364
rect 7372 23420 7436 23424
rect 7372 23364 7376 23420
rect 7376 23364 7432 23420
rect 7432 23364 7436 23420
rect 7372 23360 7436 23364
rect 7452 23420 7516 23424
rect 7452 23364 7456 23420
rect 7456 23364 7512 23420
rect 7512 23364 7516 23420
rect 7452 23360 7516 23364
rect 15101 23420 15165 23424
rect 15101 23364 15105 23420
rect 15105 23364 15161 23420
rect 15161 23364 15165 23420
rect 15101 23360 15165 23364
rect 15181 23420 15245 23424
rect 15181 23364 15185 23420
rect 15185 23364 15241 23420
rect 15241 23364 15245 23420
rect 15181 23360 15245 23364
rect 15261 23420 15325 23424
rect 15261 23364 15265 23420
rect 15265 23364 15321 23420
rect 15321 23364 15325 23420
rect 15261 23360 15325 23364
rect 15341 23420 15405 23424
rect 15341 23364 15345 23420
rect 15345 23364 15401 23420
rect 15401 23364 15405 23420
rect 15341 23360 15405 23364
rect 22990 23420 23054 23424
rect 22990 23364 22994 23420
rect 22994 23364 23050 23420
rect 23050 23364 23054 23420
rect 22990 23360 23054 23364
rect 23070 23420 23134 23424
rect 23070 23364 23074 23420
rect 23074 23364 23130 23420
rect 23130 23364 23134 23420
rect 23070 23360 23134 23364
rect 23150 23420 23214 23424
rect 23150 23364 23154 23420
rect 23154 23364 23210 23420
rect 23210 23364 23214 23420
rect 23150 23360 23214 23364
rect 23230 23420 23294 23424
rect 23230 23364 23234 23420
rect 23234 23364 23290 23420
rect 23290 23364 23294 23420
rect 23230 23360 23294 23364
rect 30879 23420 30943 23424
rect 30879 23364 30883 23420
rect 30883 23364 30939 23420
rect 30939 23364 30943 23420
rect 30879 23360 30943 23364
rect 30959 23420 31023 23424
rect 30959 23364 30963 23420
rect 30963 23364 31019 23420
rect 31019 23364 31023 23420
rect 30959 23360 31023 23364
rect 31039 23420 31103 23424
rect 31039 23364 31043 23420
rect 31043 23364 31099 23420
rect 31099 23364 31103 23420
rect 31039 23360 31103 23364
rect 31119 23420 31183 23424
rect 31119 23364 31123 23420
rect 31123 23364 31179 23420
rect 31179 23364 31183 23420
rect 31119 23360 31183 23364
rect 6552 22876 6616 22880
rect 6552 22820 6556 22876
rect 6556 22820 6612 22876
rect 6612 22820 6616 22876
rect 6552 22816 6616 22820
rect 6632 22876 6696 22880
rect 6632 22820 6636 22876
rect 6636 22820 6692 22876
rect 6692 22820 6696 22876
rect 6632 22816 6696 22820
rect 6712 22876 6776 22880
rect 6712 22820 6716 22876
rect 6716 22820 6772 22876
rect 6772 22820 6776 22876
rect 6712 22816 6776 22820
rect 6792 22876 6856 22880
rect 6792 22820 6796 22876
rect 6796 22820 6852 22876
rect 6852 22820 6856 22876
rect 6792 22816 6856 22820
rect 14441 22876 14505 22880
rect 14441 22820 14445 22876
rect 14445 22820 14501 22876
rect 14501 22820 14505 22876
rect 14441 22816 14505 22820
rect 14521 22876 14585 22880
rect 14521 22820 14525 22876
rect 14525 22820 14581 22876
rect 14581 22820 14585 22876
rect 14521 22816 14585 22820
rect 14601 22876 14665 22880
rect 14601 22820 14605 22876
rect 14605 22820 14661 22876
rect 14661 22820 14665 22876
rect 14601 22816 14665 22820
rect 14681 22876 14745 22880
rect 14681 22820 14685 22876
rect 14685 22820 14741 22876
rect 14741 22820 14745 22876
rect 14681 22816 14745 22820
rect 22330 22876 22394 22880
rect 22330 22820 22334 22876
rect 22334 22820 22390 22876
rect 22390 22820 22394 22876
rect 22330 22816 22394 22820
rect 22410 22876 22474 22880
rect 22410 22820 22414 22876
rect 22414 22820 22470 22876
rect 22470 22820 22474 22876
rect 22410 22816 22474 22820
rect 22490 22876 22554 22880
rect 22490 22820 22494 22876
rect 22494 22820 22550 22876
rect 22550 22820 22554 22876
rect 22490 22816 22554 22820
rect 22570 22876 22634 22880
rect 22570 22820 22574 22876
rect 22574 22820 22630 22876
rect 22630 22820 22634 22876
rect 22570 22816 22634 22820
rect 30219 22876 30283 22880
rect 30219 22820 30223 22876
rect 30223 22820 30279 22876
rect 30279 22820 30283 22876
rect 30219 22816 30283 22820
rect 30299 22876 30363 22880
rect 30299 22820 30303 22876
rect 30303 22820 30359 22876
rect 30359 22820 30363 22876
rect 30299 22816 30363 22820
rect 30379 22876 30443 22880
rect 30379 22820 30383 22876
rect 30383 22820 30439 22876
rect 30439 22820 30443 22876
rect 30379 22816 30443 22820
rect 30459 22876 30523 22880
rect 30459 22820 30463 22876
rect 30463 22820 30519 22876
rect 30519 22820 30523 22876
rect 30459 22816 30523 22820
rect 7212 22332 7276 22336
rect 7212 22276 7216 22332
rect 7216 22276 7272 22332
rect 7272 22276 7276 22332
rect 7212 22272 7276 22276
rect 7292 22332 7356 22336
rect 7292 22276 7296 22332
rect 7296 22276 7352 22332
rect 7352 22276 7356 22332
rect 7292 22272 7356 22276
rect 7372 22332 7436 22336
rect 7372 22276 7376 22332
rect 7376 22276 7432 22332
rect 7432 22276 7436 22332
rect 7372 22272 7436 22276
rect 7452 22332 7516 22336
rect 7452 22276 7456 22332
rect 7456 22276 7512 22332
rect 7512 22276 7516 22332
rect 7452 22272 7516 22276
rect 15101 22332 15165 22336
rect 15101 22276 15105 22332
rect 15105 22276 15161 22332
rect 15161 22276 15165 22332
rect 15101 22272 15165 22276
rect 15181 22332 15245 22336
rect 15181 22276 15185 22332
rect 15185 22276 15241 22332
rect 15241 22276 15245 22332
rect 15181 22272 15245 22276
rect 15261 22332 15325 22336
rect 15261 22276 15265 22332
rect 15265 22276 15321 22332
rect 15321 22276 15325 22332
rect 15261 22272 15325 22276
rect 15341 22332 15405 22336
rect 15341 22276 15345 22332
rect 15345 22276 15401 22332
rect 15401 22276 15405 22332
rect 15341 22272 15405 22276
rect 22990 22332 23054 22336
rect 22990 22276 22994 22332
rect 22994 22276 23050 22332
rect 23050 22276 23054 22332
rect 22990 22272 23054 22276
rect 23070 22332 23134 22336
rect 23070 22276 23074 22332
rect 23074 22276 23130 22332
rect 23130 22276 23134 22332
rect 23070 22272 23134 22276
rect 23150 22332 23214 22336
rect 23150 22276 23154 22332
rect 23154 22276 23210 22332
rect 23210 22276 23214 22332
rect 23150 22272 23214 22276
rect 23230 22332 23294 22336
rect 23230 22276 23234 22332
rect 23234 22276 23290 22332
rect 23290 22276 23294 22332
rect 23230 22272 23294 22276
rect 30879 22332 30943 22336
rect 30879 22276 30883 22332
rect 30883 22276 30939 22332
rect 30939 22276 30943 22332
rect 30879 22272 30943 22276
rect 30959 22332 31023 22336
rect 30959 22276 30963 22332
rect 30963 22276 31019 22332
rect 31019 22276 31023 22332
rect 30959 22272 31023 22276
rect 31039 22332 31103 22336
rect 31039 22276 31043 22332
rect 31043 22276 31099 22332
rect 31099 22276 31103 22332
rect 31039 22272 31103 22276
rect 31119 22332 31183 22336
rect 31119 22276 31123 22332
rect 31123 22276 31179 22332
rect 31179 22276 31183 22332
rect 31119 22272 31183 22276
rect 6552 21788 6616 21792
rect 6552 21732 6556 21788
rect 6556 21732 6612 21788
rect 6612 21732 6616 21788
rect 6552 21728 6616 21732
rect 6632 21788 6696 21792
rect 6632 21732 6636 21788
rect 6636 21732 6692 21788
rect 6692 21732 6696 21788
rect 6632 21728 6696 21732
rect 6712 21788 6776 21792
rect 6712 21732 6716 21788
rect 6716 21732 6772 21788
rect 6772 21732 6776 21788
rect 6712 21728 6776 21732
rect 6792 21788 6856 21792
rect 6792 21732 6796 21788
rect 6796 21732 6852 21788
rect 6852 21732 6856 21788
rect 6792 21728 6856 21732
rect 14441 21788 14505 21792
rect 14441 21732 14445 21788
rect 14445 21732 14501 21788
rect 14501 21732 14505 21788
rect 14441 21728 14505 21732
rect 14521 21788 14585 21792
rect 14521 21732 14525 21788
rect 14525 21732 14581 21788
rect 14581 21732 14585 21788
rect 14521 21728 14585 21732
rect 14601 21788 14665 21792
rect 14601 21732 14605 21788
rect 14605 21732 14661 21788
rect 14661 21732 14665 21788
rect 14601 21728 14665 21732
rect 14681 21788 14745 21792
rect 14681 21732 14685 21788
rect 14685 21732 14741 21788
rect 14741 21732 14745 21788
rect 14681 21728 14745 21732
rect 22330 21788 22394 21792
rect 22330 21732 22334 21788
rect 22334 21732 22390 21788
rect 22390 21732 22394 21788
rect 22330 21728 22394 21732
rect 22410 21788 22474 21792
rect 22410 21732 22414 21788
rect 22414 21732 22470 21788
rect 22470 21732 22474 21788
rect 22410 21728 22474 21732
rect 22490 21788 22554 21792
rect 22490 21732 22494 21788
rect 22494 21732 22550 21788
rect 22550 21732 22554 21788
rect 22490 21728 22554 21732
rect 22570 21788 22634 21792
rect 22570 21732 22574 21788
rect 22574 21732 22630 21788
rect 22630 21732 22634 21788
rect 22570 21728 22634 21732
rect 30219 21788 30283 21792
rect 30219 21732 30223 21788
rect 30223 21732 30279 21788
rect 30279 21732 30283 21788
rect 30219 21728 30283 21732
rect 30299 21788 30363 21792
rect 30299 21732 30303 21788
rect 30303 21732 30359 21788
rect 30359 21732 30363 21788
rect 30299 21728 30363 21732
rect 30379 21788 30443 21792
rect 30379 21732 30383 21788
rect 30383 21732 30439 21788
rect 30439 21732 30443 21788
rect 30379 21728 30443 21732
rect 30459 21788 30523 21792
rect 30459 21732 30463 21788
rect 30463 21732 30519 21788
rect 30519 21732 30523 21788
rect 30459 21728 30523 21732
rect 11836 21660 11900 21724
rect 7212 21244 7276 21248
rect 7212 21188 7216 21244
rect 7216 21188 7272 21244
rect 7272 21188 7276 21244
rect 7212 21184 7276 21188
rect 7292 21244 7356 21248
rect 7292 21188 7296 21244
rect 7296 21188 7352 21244
rect 7352 21188 7356 21244
rect 7292 21184 7356 21188
rect 7372 21244 7436 21248
rect 7372 21188 7376 21244
rect 7376 21188 7432 21244
rect 7432 21188 7436 21244
rect 7372 21184 7436 21188
rect 7452 21244 7516 21248
rect 7452 21188 7456 21244
rect 7456 21188 7512 21244
rect 7512 21188 7516 21244
rect 7452 21184 7516 21188
rect 15101 21244 15165 21248
rect 15101 21188 15105 21244
rect 15105 21188 15161 21244
rect 15161 21188 15165 21244
rect 15101 21184 15165 21188
rect 15181 21244 15245 21248
rect 15181 21188 15185 21244
rect 15185 21188 15241 21244
rect 15241 21188 15245 21244
rect 15181 21184 15245 21188
rect 15261 21244 15325 21248
rect 15261 21188 15265 21244
rect 15265 21188 15321 21244
rect 15321 21188 15325 21244
rect 15261 21184 15325 21188
rect 15341 21244 15405 21248
rect 15341 21188 15345 21244
rect 15345 21188 15401 21244
rect 15401 21188 15405 21244
rect 15341 21184 15405 21188
rect 22990 21244 23054 21248
rect 22990 21188 22994 21244
rect 22994 21188 23050 21244
rect 23050 21188 23054 21244
rect 22990 21184 23054 21188
rect 23070 21244 23134 21248
rect 23070 21188 23074 21244
rect 23074 21188 23130 21244
rect 23130 21188 23134 21244
rect 23070 21184 23134 21188
rect 23150 21244 23214 21248
rect 23150 21188 23154 21244
rect 23154 21188 23210 21244
rect 23210 21188 23214 21244
rect 23150 21184 23214 21188
rect 23230 21244 23294 21248
rect 23230 21188 23234 21244
rect 23234 21188 23290 21244
rect 23290 21188 23294 21244
rect 23230 21184 23294 21188
rect 30879 21244 30943 21248
rect 30879 21188 30883 21244
rect 30883 21188 30939 21244
rect 30939 21188 30943 21244
rect 30879 21184 30943 21188
rect 30959 21244 31023 21248
rect 30959 21188 30963 21244
rect 30963 21188 31019 21244
rect 31019 21188 31023 21244
rect 30959 21184 31023 21188
rect 31039 21244 31103 21248
rect 31039 21188 31043 21244
rect 31043 21188 31099 21244
rect 31099 21188 31103 21244
rect 31039 21184 31103 21188
rect 31119 21244 31183 21248
rect 31119 21188 31123 21244
rect 31123 21188 31179 21244
rect 31179 21188 31183 21244
rect 31119 21184 31183 21188
rect 19380 20708 19444 20772
rect 6552 20700 6616 20704
rect 6552 20644 6556 20700
rect 6556 20644 6612 20700
rect 6612 20644 6616 20700
rect 6552 20640 6616 20644
rect 6632 20700 6696 20704
rect 6632 20644 6636 20700
rect 6636 20644 6692 20700
rect 6692 20644 6696 20700
rect 6632 20640 6696 20644
rect 6712 20700 6776 20704
rect 6712 20644 6716 20700
rect 6716 20644 6772 20700
rect 6772 20644 6776 20700
rect 6712 20640 6776 20644
rect 6792 20700 6856 20704
rect 6792 20644 6796 20700
rect 6796 20644 6852 20700
rect 6852 20644 6856 20700
rect 6792 20640 6856 20644
rect 14441 20700 14505 20704
rect 14441 20644 14445 20700
rect 14445 20644 14501 20700
rect 14501 20644 14505 20700
rect 14441 20640 14505 20644
rect 14521 20700 14585 20704
rect 14521 20644 14525 20700
rect 14525 20644 14581 20700
rect 14581 20644 14585 20700
rect 14521 20640 14585 20644
rect 14601 20700 14665 20704
rect 14601 20644 14605 20700
rect 14605 20644 14661 20700
rect 14661 20644 14665 20700
rect 14601 20640 14665 20644
rect 14681 20700 14745 20704
rect 14681 20644 14685 20700
rect 14685 20644 14741 20700
rect 14741 20644 14745 20700
rect 14681 20640 14745 20644
rect 22330 20700 22394 20704
rect 22330 20644 22334 20700
rect 22334 20644 22390 20700
rect 22390 20644 22394 20700
rect 22330 20640 22394 20644
rect 22410 20700 22474 20704
rect 22410 20644 22414 20700
rect 22414 20644 22470 20700
rect 22470 20644 22474 20700
rect 22410 20640 22474 20644
rect 22490 20700 22554 20704
rect 22490 20644 22494 20700
rect 22494 20644 22550 20700
rect 22550 20644 22554 20700
rect 22490 20640 22554 20644
rect 22570 20700 22634 20704
rect 22570 20644 22574 20700
rect 22574 20644 22630 20700
rect 22630 20644 22634 20700
rect 22570 20640 22634 20644
rect 30219 20700 30283 20704
rect 30219 20644 30223 20700
rect 30223 20644 30279 20700
rect 30279 20644 30283 20700
rect 30219 20640 30283 20644
rect 30299 20700 30363 20704
rect 30299 20644 30303 20700
rect 30303 20644 30359 20700
rect 30359 20644 30363 20700
rect 30299 20640 30363 20644
rect 30379 20700 30443 20704
rect 30379 20644 30383 20700
rect 30383 20644 30439 20700
rect 30439 20644 30443 20700
rect 30379 20640 30443 20644
rect 30459 20700 30523 20704
rect 30459 20644 30463 20700
rect 30463 20644 30519 20700
rect 30519 20644 30523 20700
rect 30459 20640 30523 20644
rect 11836 20496 11900 20500
rect 11836 20440 11886 20496
rect 11886 20440 11900 20496
rect 11836 20436 11900 20440
rect 12204 20436 12268 20500
rect 6132 20164 6196 20228
rect 7212 20156 7276 20160
rect 7212 20100 7216 20156
rect 7216 20100 7272 20156
rect 7272 20100 7276 20156
rect 7212 20096 7276 20100
rect 7292 20156 7356 20160
rect 7292 20100 7296 20156
rect 7296 20100 7352 20156
rect 7352 20100 7356 20156
rect 7292 20096 7356 20100
rect 7372 20156 7436 20160
rect 7372 20100 7376 20156
rect 7376 20100 7432 20156
rect 7432 20100 7436 20156
rect 7372 20096 7436 20100
rect 7452 20156 7516 20160
rect 7452 20100 7456 20156
rect 7456 20100 7512 20156
rect 7512 20100 7516 20156
rect 7452 20096 7516 20100
rect 15101 20156 15165 20160
rect 15101 20100 15105 20156
rect 15105 20100 15161 20156
rect 15161 20100 15165 20156
rect 15101 20096 15165 20100
rect 15181 20156 15245 20160
rect 15181 20100 15185 20156
rect 15185 20100 15241 20156
rect 15241 20100 15245 20156
rect 15181 20096 15245 20100
rect 15261 20156 15325 20160
rect 15261 20100 15265 20156
rect 15265 20100 15321 20156
rect 15321 20100 15325 20156
rect 15261 20096 15325 20100
rect 15341 20156 15405 20160
rect 15341 20100 15345 20156
rect 15345 20100 15401 20156
rect 15401 20100 15405 20156
rect 15341 20096 15405 20100
rect 22990 20156 23054 20160
rect 22990 20100 22994 20156
rect 22994 20100 23050 20156
rect 23050 20100 23054 20156
rect 22990 20096 23054 20100
rect 23070 20156 23134 20160
rect 23070 20100 23074 20156
rect 23074 20100 23130 20156
rect 23130 20100 23134 20156
rect 23070 20096 23134 20100
rect 23150 20156 23214 20160
rect 23150 20100 23154 20156
rect 23154 20100 23210 20156
rect 23210 20100 23214 20156
rect 23150 20096 23214 20100
rect 23230 20156 23294 20160
rect 23230 20100 23234 20156
rect 23234 20100 23290 20156
rect 23290 20100 23294 20156
rect 23230 20096 23294 20100
rect 30879 20156 30943 20160
rect 30879 20100 30883 20156
rect 30883 20100 30939 20156
rect 30939 20100 30943 20156
rect 30879 20096 30943 20100
rect 30959 20156 31023 20160
rect 30959 20100 30963 20156
rect 30963 20100 31019 20156
rect 31019 20100 31023 20156
rect 30959 20096 31023 20100
rect 31039 20156 31103 20160
rect 31039 20100 31043 20156
rect 31043 20100 31099 20156
rect 31099 20100 31103 20156
rect 31039 20096 31103 20100
rect 31119 20156 31183 20160
rect 31119 20100 31123 20156
rect 31123 20100 31179 20156
rect 31179 20100 31183 20156
rect 31119 20096 31183 20100
rect 6552 19612 6616 19616
rect 6552 19556 6556 19612
rect 6556 19556 6612 19612
rect 6612 19556 6616 19612
rect 6552 19552 6616 19556
rect 6632 19612 6696 19616
rect 6632 19556 6636 19612
rect 6636 19556 6692 19612
rect 6692 19556 6696 19612
rect 6632 19552 6696 19556
rect 6712 19612 6776 19616
rect 6712 19556 6716 19612
rect 6716 19556 6772 19612
rect 6772 19556 6776 19612
rect 6712 19552 6776 19556
rect 6792 19612 6856 19616
rect 6792 19556 6796 19612
rect 6796 19556 6852 19612
rect 6852 19556 6856 19612
rect 6792 19552 6856 19556
rect 14441 19612 14505 19616
rect 14441 19556 14445 19612
rect 14445 19556 14501 19612
rect 14501 19556 14505 19612
rect 14441 19552 14505 19556
rect 14521 19612 14585 19616
rect 14521 19556 14525 19612
rect 14525 19556 14581 19612
rect 14581 19556 14585 19612
rect 14521 19552 14585 19556
rect 14601 19612 14665 19616
rect 14601 19556 14605 19612
rect 14605 19556 14661 19612
rect 14661 19556 14665 19612
rect 14601 19552 14665 19556
rect 14681 19612 14745 19616
rect 14681 19556 14685 19612
rect 14685 19556 14741 19612
rect 14741 19556 14745 19612
rect 14681 19552 14745 19556
rect 22330 19612 22394 19616
rect 22330 19556 22334 19612
rect 22334 19556 22390 19612
rect 22390 19556 22394 19612
rect 22330 19552 22394 19556
rect 22410 19612 22474 19616
rect 22410 19556 22414 19612
rect 22414 19556 22470 19612
rect 22470 19556 22474 19612
rect 22410 19552 22474 19556
rect 22490 19612 22554 19616
rect 22490 19556 22494 19612
rect 22494 19556 22550 19612
rect 22550 19556 22554 19612
rect 22490 19552 22554 19556
rect 22570 19612 22634 19616
rect 22570 19556 22574 19612
rect 22574 19556 22630 19612
rect 22630 19556 22634 19612
rect 22570 19552 22634 19556
rect 30219 19612 30283 19616
rect 30219 19556 30223 19612
rect 30223 19556 30279 19612
rect 30279 19556 30283 19612
rect 30219 19552 30283 19556
rect 30299 19612 30363 19616
rect 30299 19556 30303 19612
rect 30303 19556 30359 19612
rect 30359 19556 30363 19612
rect 30299 19552 30363 19556
rect 30379 19612 30443 19616
rect 30379 19556 30383 19612
rect 30383 19556 30439 19612
rect 30439 19556 30443 19612
rect 30379 19552 30443 19556
rect 30459 19612 30523 19616
rect 30459 19556 30463 19612
rect 30463 19556 30519 19612
rect 30519 19556 30523 19612
rect 30459 19552 30523 19556
rect 7212 19068 7276 19072
rect 7212 19012 7216 19068
rect 7216 19012 7272 19068
rect 7272 19012 7276 19068
rect 7212 19008 7276 19012
rect 7292 19068 7356 19072
rect 7292 19012 7296 19068
rect 7296 19012 7352 19068
rect 7352 19012 7356 19068
rect 7292 19008 7356 19012
rect 7372 19068 7436 19072
rect 7372 19012 7376 19068
rect 7376 19012 7432 19068
rect 7432 19012 7436 19068
rect 7372 19008 7436 19012
rect 7452 19068 7516 19072
rect 7452 19012 7456 19068
rect 7456 19012 7512 19068
rect 7512 19012 7516 19068
rect 7452 19008 7516 19012
rect 15101 19068 15165 19072
rect 15101 19012 15105 19068
rect 15105 19012 15161 19068
rect 15161 19012 15165 19068
rect 15101 19008 15165 19012
rect 15181 19068 15245 19072
rect 15181 19012 15185 19068
rect 15185 19012 15241 19068
rect 15241 19012 15245 19068
rect 15181 19008 15245 19012
rect 15261 19068 15325 19072
rect 15261 19012 15265 19068
rect 15265 19012 15321 19068
rect 15321 19012 15325 19068
rect 15261 19008 15325 19012
rect 15341 19068 15405 19072
rect 15341 19012 15345 19068
rect 15345 19012 15401 19068
rect 15401 19012 15405 19068
rect 15341 19008 15405 19012
rect 22990 19068 23054 19072
rect 22990 19012 22994 19068
rect 22994 19012 23050 19068
rect 23050 19012 23054 19068
rect 22990 19008 23054 19012
rect 23070 19068 23134 19072
rect 23070 19012 23074 19068
rect 23074 19012 23130 19068
rect 23130 19012 23134 19068
rect 23070 19008 23134 19012
rect 23150 19068 23214 19072
rect 23150 19012 23154 19068
rect 23154 19012 23210 19068
rect 23210 19012 23214 19068
rect 23150 19008 23214 19012
rect 23230 19068 23294 19072
rect 23230 19012 23234 19068
rect 23234 19012 23290 19068
rect 23290 19012 23294 19068
rect 23230 19008 23294 19012
rect 30879 19068 30943 19072
rect 30879 19012 30883 19068
rect 30883 19012 30939 19068
rect 30939 19012 30943 19068
rect 30879 19008 30943 19012
rect 30959 19068 31023 19072
rect 30959 19012 30963 19068
rect 30963 19012 31019 19068
rect 31019 19012 31023 19068
rect 30959 19008 31023 19012
rect 31039 19068 31103 19072
rect 31039 19012 31043 19068
rect 31043 19012 31099 19068
rect 31099 19012 31103 19068
rect 31039 19008 31103 19012
rect 31119 19068 31183 19072
rect 31119 19012 31123 19068
rect 31123 19012 31179 19068
rect 31179 19012 31183 19068
rect 31119 19008 31183 19012
rect 6552 18524 6616 18528
rect 6552 18468 6556 18524
rect 6556 18468 6612 18524
rect 6612 18468 6616 18524
rect 6552 18464 6616 18468
rect 6632 18524 6696 18528
rect 6632 18468 6636 18524
rect 6636 18468 6692 18524
rect 6692 18468 6696 18524
rect 6632 18464 6696 18468
rect 6712 18524 6776 18528
rect 6712 18468 6716 18524
rect 6716 18468 6772 18524
rect 6772 18468 6776 18524
rect 6712 18464 6776 18468
rect 6792 18524 6856 18528
rect 6792 18468 6796 18524
rect 6796 18468 6852 18524
rect 6852 18468 6856 18524
rect 6792 18464 6856 18468
rect 14441 18524 14505 18528
rect 14441 18468 14445 18524
rect 14445 18468 14501 18524
rect 14501 18468 14505 18524
rect 14441 18464 14505 18468
rect 14521 18524 14585 18528
rect 14521 18468 14525 18524
rect 14525 18468 14581 18524
rect 14581 18468 14585 18524
rect 14521 18464 14585 18468
rect 14601 18524 14665 18528
rect 14601 18468 14605 18524
rect 14605 18468 14661 18524
rect 14661 18468 14665 18524
rect 14601 18464 14665 18468
rect 14681 18524 14745 18528
rect 14681 18468 14685 18524
rect 14685 18468 14741 18524
rect 14741 18468 14745 18524
rect 14681 18464 14745 18468
rect 22330 18524 22394 18528
rect 22330 18468 22334 18524
rect 22334 18468 22390 18524
rect 22390 18468 22394 18524
rect 22330 18464 22394 18468
rect 22410 18524 22474 18528
rect 22410 18468 22414 18524
rect 22414 18468 22470 18524
rect 22470 18468 22474 18524
rect 22410 18464 22474 18468
rect 22490 18524 22554 18528
rect 22490 18468 22494 18524
rect 22494 18468 22550 18524
rect 22550 18468 22554 18524
rect 22490 18464 22554 18468
rect 22570 18524 22634 18528
rect 22570 18468 22574 18524
rect 22574 18468 22630 18524
rect 22630 18468 22634 18524
rect 22570 18464 22634 18468
rect 30219 18524 30283 18528
rect 30219 18468 30223 18524
rect 30223 18468 30279 18524
rect 30279 18468 30283 18524
rect 30219 18464 30283 18468
rect 30299 18524 30363 18528
rect 30299 18468 30303 18524
rect 30303 18468 30359 18524
rect 30359 18468 30363 18524
rect 30299 18464 30363 18468
rect 30379 18524 30443 18528
rect 30379 18468 30383 18524
rect 30383 18468 30439 18524
rect 30439 18468 30443 18524
rect 30379 18464 30443 18468
rect 30459 18524 30523 18528
rect 30459 18468 30463 18524
rect 30463 18468 30519 18524
rect 30519 18468 30523 18524
rect 30459 18464 30523 18468
rect 7212 17980 7276 17984
rect 7212 17924 7216 17980
rect 7216 17924 7272 17980
rect 7272 17924 7276 17980
rect 7212 17920 7276 17924
rect 7292 17980 7356 17984
rect 7292 17924 7296 17980
rect 7296 17924 7352 17980
rect 7352 17924 7356 17980
rect 7292 17920 7356 17924
rect 7372 17980 7436 17984
rect 7372 17924 7376 17980
rect 7376 17924 7432 17980
rect 7432 17924 7436 17980
rect 7372 17920 7436 17924
rect 7452 17980 7516 17984
rect 7452 17924 7456 17980
rect 7456 17924 7512 17980
rect 7512 17924 7516 17980
rect 7452 17920 7516 17924
rect 15101 17980 15165 17984
rect 15101 17924 15105 17980
rect 15105 17924 15161 17980
rect 15161 17924 15165 17980
rect 15101 17920 15165 17924
rect 15181 17980 15245 17984
rect 15181 17924 15185 17980
rect 15185 17924 15241 17980
rect 15241 17924 15245 17980
rect 15181 17920 15245 17924
rect 15261 17980 15325 17984
rect 15261 17924 15265 17980
rect 15265 17924 15321 17980
rect 15321 17924 15325 17980
rect 15261 17920 15325 17924
rect 15341 17980 15405 17984
rect 15341 17924 15345 17980
rect 15345 17924 15401 17980
rect 15401 17924 15405 17980
rect 15341 17920 15405 17924
rect 19564 18048 19628 18052
rect 19564 17992 19578 18048
rect 19578 17992 19628 18048
rect 19564 17988 19628 17992
rect 22990 17980 23054 17984
rect 22990 17924 22994 17980
rect 22994 17924 23050 17980
rect 23050 17924 23054 17980
rect 22990 17920 23054 17924
rect 23070 17980 23134 17984
rect 23070 17924 23074 17980
rect 23074 17924 23130 17980
rect 23130 17924 23134 17980
rect 23070 17920 23134 17924
rect 23150 17980 23214 17984
rect 23150 17924 23154 17980
rect 23154 17924 23210 17980
rect 23210 17924 23214 17980
rect 23150 17920 23214 17924
rect 23230 17980 23294 17984
rect 23230 17924 23234 17980
rect 23234 17924 23290 17980
rect 23290 17924 23294 17980
rect 23230 17920 23294 17924
rect 30879 17980 30943 17984
rect 30879 17924 30883 17980
rect 30883 17924 30939 17980
rect 30939 17924 30943 17980
rect 30879 17920 30943 17924
rect 30959 17980 31023 17984
rect 30959 17924 30963 17980
rect 30963 17924 31019 17980
rect 31019 17924 31023 17980
rect 30959 17920 31023 17924
rect 31039 17980 31103 17984
rect 31039 17924 31043 17980
rect 31043 17924 31099 17980
rect 31099 17924 31103 17980
rect 31039 17920 31103 17924
rect 31119 17980 31183 17984
rect 31119 17924 31123 17980
rect 31123 17924 31179 17980
rect 31179 17924 31183 17980
rect 31119 17920 31183 17924
rect 19748 17912 19812 17916
rect 19748 17856 19762 17912
rect 19762 17856 19812 17912
rect 19748 17852 19812 17856
rect 22140 17716 22204 17780
rect 6552 17436 6616 17440
rect 6552 17380 6556 17436
rect 6556 17380 6612 17436
rect 6612 17380 6616 17436
rect 6552 17376 6616 17380
rect 6632 17436 6696 17440
rect 6632 17380 6636 17436
rect 6636 17380 6692 17436
rect 6692 17380 6696 17436
rect 6632 17376 6696 17380
rect 6712 17436 6776 17440
rect 6712 17380 6716 17436
rect 6716 17380 6772 17436
rect 6772 17380 6776 17436
rect 6712 17376 6776 17380
rect 6792 17436 6856 17440
rect 6792 17380 6796 17436
rect 6796 17380 6852 17436
rect 6852 17380 6856 17436
rect 6792 17376 6856 17380
rect 14441 17436 14505 17440
rect 14441 17380 14445 17436
rect 14445 17380 14501 17436
rect 14501 17380 14505 17436
rect 14441 17376 14505 17380
rect 14521 17436 14585 17440
rect 14521 17380 14525 17436
rect 14525 17380 14581 17436
rect 14581 17380 14585 17436
rect 14521 17376 14585 17380
rect 14601 17436 14665 17440
rect 14601 17380 14605 17436
rect 14605 17380 14661 17436
rect 14661 17380 14665 17436
rect 14601 17376 14665 17380
rect 14681 17436 14745 17440
rect 14681 17380 14685 17436
rect 14685 17380 14741 17436
rect 14741 17380 14745 17436
rect 14681 17376 14745 17380
rect 22330 17436 22394 17440
rect 22330 17380 22334 17436
rect 22334 17380 22390 17436
rect 22390 17380 22394 17436
rect 22330 17376 22394 17380
rect 22410 17436 22474 17440
rect 22410 17380 22414 17436
rect 22414 17380 22470 17436
rect 22470 17380 22474 17436
rect 22410 17376 22474 17380
rect 22490 17436 22554 17440
rect 22490 17380 22494 17436
rect 22494 17380 22550 17436
rect 22550 17380 22554 17436
rect 22490 17376 22554 17380
rect 22570 17436 22634 17440
rect 22570 17380 22574 17436
rect 22574 17380 22630 17436
rect 22630 17380 22634 17436
rect 22570 17376 22634 17380
rect 30219 17436 30283 17440
rect 30219 17380 30223 17436
rect 30223 17380 30279 17436
rect 30279 17380 30283 17436
rect 30219 17376 30283 17380
rect 30299 17436 30363 17440
rect 30299 17380 30303 17436
rect 30303 17380 30359 17436
rect 30359 17380 30363 17436
rect 30299 17376 30363 17380
rect 30379 17436 30443 17440
rect 30379 17380 30383 17436
rect 30383 17380 30439 17436
rect 30439 17380 30443 17436
rect 30379 17376 30443 17380
rect 30459 17436 30523 17440
rect 30459 17380 30463 17436
rect 30463 17380 30519 17436
rect 30519 17380 30523 17436
rect 30459 17376 30523 17380
rect 7212 16892 7276 16896
rect 7212 16836 7216 16892
rect 7216 16836 7272 16892
rect 7272 16836 7276 16892
rect 7212 16832 7276 16836
rect 7292 16892 7356 16896
rect 7292 16836 7296 16892
rect 7296 16836 7352 16892
rect 7352 16836 7356 16892
rect 7292 16832 7356 16836
rect 7372 16892 7436 16896
rect 7372 16836 7376 16892
rect 7376 16836 7432 16892
rect 7432 16836 7436 16892
rect 7372 16832 7436 16836
rect 7452 16892 7516 16896
rect 7452 16836 7456 16892
rect 7456 16836 7512 16892
rect 7512 16836 7516 16892
rect 7452 16832 7516 16836
rect 15101 16892 15165 16896
rect 15101 16836 15105 16892
rect 15105 16836 15161 16892
rect 15161 16836 15165 16892
rect 15101 16832 15165 16836
rect 15181 16892 15245 16896
rect 15181 16836 15185 16892
rect 15185 16836 15241 16892
rect 15241 16836 15245 16892
rect 15181 16832 15245 16836
rect 15261 16892 15325 16896
rect 15261 16836 15265 16892
rect 15265 16836 15321 16892
rect 15321 16836 15325 16892
rect 15261 16832 15325 16836
rect 15341 16892 15405 16896
rect 15341 16836 15345 16892
rect 15345 16836 15401 16892
rect 15401 16836 15405 16892
rect 15341 16832 15405 16836
rect 22990 16892 23054 16896
rect 22990 16836 22994 16892
rect 22994 16836 23050 16892
rect 23050 16836 23054 16892
rect 22990 16832 23054 16836
rect 23070 16892 23134 16896
rect 23070 16836 23074 16892
rect 23074 16836 23130 16892
rect 23130 16836 23134 16892
rect 23070 16832 23134 16836
rect 23150 16892 23214 16896
rect 23150 16836 23154 16892
rect 23154 16836 23210 16892
rect 23210 16836 23214 16892
rect 23150 16832 23214 16836
rect 23230 16892 23294 16896
rect 23230 16836 23234 16892
rect 23234 16836 23290 16892
rect 23290 16836 23294 16892
rect 23230 16832 23294 16836
rect 30879 16892 30943 16896
rect 30879 16836 30883 16892
rect 30883 16836 30939 16892
rect 30939 16836 30943 16892
rect 30879 16832 30943 16836
rect 30959 16892 31023 16896
rect 30959 16836 30963 16892
rect 30963 16836 31019 16892
rect 31019 16836 31023 16892
rect 30959 16832 31023 16836
rect 31039 16892 31103 16896
rect 31039 16836 31043 16892
rect 31043 16836 31099 16892
rect 31099 16836 31103 16892
rect 31039 16832 31103 16836
rect 31119 16892 31183 16896
rect 31119 16836 31123 16892
rect 31123 16836 31179 16892
rect 31179 16836 31183 16892
rect 31119 16832 31183 16836
rect 6552 16348 6616 16352
rect 6552 16292 6556 16348
rect 6556 16292 6612 16348
rect 6612 16292 6616 16348
rect 6552 16288 6616 16292
rect 6632 16348 6696 16352
rect 6632 16292 6636 16348
rect 6636 16292 6692 16348
rect 6692 16292 6696 16348
rect 6632 16288 6696 16292
rect 6712 16348 6776 16352
rect 6712 16292 6716 16348
rect 6716 16292 6772 16348
rect 6772 16292 6776 16348
rect 6712 16288 6776 16292
rect 6792 16348 6856 16352
rect 6792 16292 6796 16348
rect 6796 16292 6852 16348
rect 6852 16292 6856 16348
rect 6792 16288 6856 16292
rect 14441 16348 14505 16352
rect 14441 16292 14445 16348
rect 14445 16292 14501 16348
rect 14501 16292 14505 16348
rect 14441 16288 14505 16292
rect 14521 16348 14585 16352
rect 14521 16292 14525 16348
rect 14525 16292 14581 16348
rect 14581 16292 14585 16348
rect 14521 16288 14585 16292
rect 14601 16348 14665 16352
rect 14601 16292 14605 16348
rect 14605 16292 14661 16348
rect 14661 16292 14665 16348
rect 14601 16288 14665 16292
rect 14681 16348 14745 16352
rect 14681 16292 14685 16348
rect 14685 16292 14741 16348
rect 14741 16292 14745 16348
rect 14681 16288 14745 16292
rect 22330 16348 22394 16352
rect 22330 16292 22334 16348
rect 22334 16292 22390 16348
rect 22390 16292 22394 16348
rect 22330 16288 22394 16292
rect 22410 16348 22474 16352
rect 22410 16292 22414 16348
rect 22414 16292 22470 16348
rect 22470 16292 22474 16348
rect 22410 16288 22474 16292
rect 22490 16348 22554 16352
rect 22490 16292 22494 16348
rect 22494 16292 22550 16348
rect 22550 16292 22554 16348
rect 22490 16288 22554 16292
rect 22570 16348 22634 16352
rect 22570 16292 22574 16348
rect 22574 16292 22630 16348
rect 22630 16292 22634 16348
rect 22570 16288 22634 16292
rect 30219 16348 30283 16352
rect 30219 16292 30223 16348
rect 30223 16292 30279 16348
rect 30279 16292 30283 16348
rect 30219 16288 30283 16292
rect 30299 16348 30363 16352
rect 30299 16292 30303 16348
rect 30303 16292 30359 16348
rect 30359 16292 30363 16348
rect 30299 16288 30363 16292
rect 30379 16348 30443 16352
rect 30379 16292 30383 16348
rect 30383 16292 30439 16348
rect 30439 16292 30443 16348
rect 30379 16288 30443 16292
rect 30459 16348 30523 16352
rect 30459 16292 30463 16348
rect 30463 16292 30519 16348
rect 30519 16292 30523 16348
rect 30459 16288 30523 16292
rect 7212 15804 7276 15808
rect 7212 15748 7216 15804
rect 7216 15748 7272 15804
rect 7272 15748 7276 15804
rect 7212 15744 7276 15748
rect 7292 15804 7356 15808
rect 7292 15748 7296 15804
rect 7296 15748 7352 15804
rect 7352 15748 7356 15804
rect 7292 15744 7356 15748
rect 7372 15804 7436 15808
rect 7372 15748 7376 15804
rect 7376 15748 7432 15804
rect 7432 15748 7436 15804
rect 7372 15744 7436 15748
rect 7452 15804 7516 15808
rect 7452 15748 7456 15804
rect 7456 15748 7512 15804
rect 7512 15748 7516 15804
rect 7452 15744 7516 15748
rect 15101 15804 15165 15808
rect 15101 15748 15105 15804
rect 15105 15748 15161 15804
rect 15161 15748 15165 15804
rect 15101 15744 15165 15748
rect 15181 15804 15245 15808
rect 15181 15748 15185 15804
rect 15185 15748 15241 15804
rect 15241 15748 15245 15804
rect 15181 15744 15245 15748
rect 15261 15804 15325 15808
rect 15261 15748 15265 15804
rect 15265 15748 15321 15804
rect 15321 15748 15325 15804
rect 15261 15744 15325 15748
rect 15341 15804 15405 15808
rect 15341 15748 15345 15804
rect 15345 15748 15401 15804
rect 15401 15748 15405 15804
rect 15341 15744 15405 15748
rect 22990 15804 23054 15808
rect 22990 15748 22994 15804
rect 22994 15748 23050 15804
rect 23050 15748 23054 15804
rect 22990 15744 23054 15748
rect 23070 15804 23134 15808
rect 23070 15748 23074 15804
rect 23074 15748 23130 15804
rect 23130 15748 23134 15804
rect 23070 15744 23134 15748
rect 23150 15804 23214 15808
rect 23150 15748 23154 15804
rect 23154 15748 23210 15804
rect 23210 15748 23214 15804
rect 23150 15744 23214 15748
rect 23230 15804 23294 15808
rect 23230 15748 23234 15804
rect 23234 15748 23290 15804
rect 23290 15748 23294 15804
rect 23230 15744 23294 15748
rect 30879 15804 30943 15808
rect 30879 15748 30883 15804
rect 30883 15748 30939 15804
rect 30939 15748 30943 15804
rect 30879 15744 30943 15748
rect 30959 15804 31023 15808
rect 30959 15748 30963 15804
rect 30963 15748 31019 15804
rect 31019 15748 31023 15804
rect 30959 15744 31023 15748
rect 31039 15804 31103 15808
rect 31039 15748 31043 15804
rect 31043 15748 31099 15804
rect 31099 15748 31103 15804
rect 31039 15744 31103 15748
rect 31119 15804 31183 15808
rect 31119 15748 31123 15804
rect 31123 15748 31179 15804
rect 31179 15748 31183 15804
rect 31119 15744 31183 15748
rect 18828 15268 18892 15332
rect 6552 15260 6616 15264
rect 6552 15204 6556 15260
rect 6556 15204 6612 15260
rect 6612 15204 6616 15260
rect 6552 15200 6616 15204
rect 6632 15260 6696 15264
rect 6632 15204 6636 15260
rect 6636 15204 6692 15260
rect 6692 15204 6696 15260
rect 6632 15200 6696 15204
rect 6712 15260 6776 15264
rect 6712 15204 6716 15260
rect 6716 15204 6772 15260
rect 6772 15204 6776 15260
rect 6712 15200 6776 15204
rect 6792 15260 6856 15264
rect 6792 15204 6796 15260
rect 6796 15204 6852 15260
rect 6852 15204 6856 15260
rect 6792 15200 6856 15204
rect 14441 15260 14505 15264
rect 14441 15204 14445 15260
rect 14445 15204 14501 15260
rect 14501 15204 14505 15260
rect 14441 15200 14505 15204
rect 14521 15260 14585 15264
rect 14521 15204 14525 15260
rect 14525 15204 14581 15260
rect 14581 15204 14585 15260
rect 14521 15200 14585 15204
rect 14601 15260 14665 15264
rect 14601 15204 14605 15260
rect 14605 15204 14661 15260
rect 14661 15204 14665 15260
rect 14601 15200 14665 15204
rect 14681 15260 14745 15264
rect 14681 15204 14685 15260
rect 14685 15204 14741 15260
rect 14741 15204 14745 15260
rect 14681 15200 14745 15204
rect 22330 15260 22394 15264
rect 22330 15204 22334 15260
rect 22334 15204 22390 15260
rect 22390 15204 22394 15260
rect 22330 15200 22394 15204
rect 22410 15260 22474 15264
rect 22410 15204 22414 15260
rect 22414 15204 22470 15260
rect 22470 15204 22474 15260
rect 22410 15200 22474 15204
rect 22490 15260 22554 15264
rect 22490 15204 22494 15260
rect 22494 15204 22550 15260
rect 22550 15204 22554 15260
rect 22490 15200 22554 15204
rect 22570 15260 22634 15264
rect 22570 15204 22574 15260
rect 22574 15204 22630 15260
rect 22630 15204 22634 15260
rect 22570 15200 22634 15204
rect 30219 15260 30283 15264
rect 30219 15204 30223 15260
rect 30223 15204 30279 15260
rect 30279 15204 30283 15260
rect 30219 15200 30283 15204
rect 30299 15260 30363 15264
rect 30299 15204 30303 15260
rect 30303 15204 30359 15260
rect 30359 15204 30363 15260
rect 30299 15200 30363 15204
rect 30379 15260 30443 15264
rect 30379 15204 30383 15260
rect 30383 15204 30439 15260
rect 30439 15204 30443 15260
rect 30379 15200 30443 15204
rect 30459 15260 30523 15264
rect 30459 15204 30463 15260
rect 30463 15204 30519 15260
rect 30519 15204 30523 15260
rect 30459 15200 30523 15204
rect 5580 15132 5644 15196
rect 19748 15132 19812 15196
rect 7212 14716 7276 14720
rect 7212 14660 7216 14716
rect 7216 14660 7272 14716
rect 7272 14660 7276 14716
rect 7212 14656 7276 14660
rect 7292 14716 7356 14720
rect 7292 14660 7296 14716
rect 7296 14660 7352 14716
rect 7352 14660 7356 14716
rect 7292 14656 7356 14660
rect 7372 14716 7436 14720
rect 7372 14660 7376 14716
rect 7376 14660 7432 14716
rect 7432 14660 7436 14716
rect 7372 14656 7436 14660
rect 7452 14716 7516 14720
rect 7452 14660 7456 14716
rect 7456 14660 7512 14716
rect 7512 14660 7516 14716
rect 7452 14656 7516 14660
rect 15101 14716 15165 14720
rect 15101 14660 15105 14716
rect 15105 14660 15161 14716
rect 15161 14660 15165 14716
rect 15101 14656 15165 14660
rect 15181 14716 15245 14720
rect 15181 14660 15185 14716
rect 15185 14660 15241 14716
rect 15241 14660 15245 14716
rect 15181 14656 15245 14660
rect 15261 14716 15325 14720
rect 15261 14660 15265 14716
rect 15265 14660 15321 14716
rect 15321 14660 15325 14716
rect 15261 14656 15325 14660
rect 15341 14716 15405 14720
rect 15341 14660 15345 14716
rect 15345 14660 15401 14716
rect 15401 14660 15405 14716
rect 15341 14656 15405 14660
rect 22990 14716 23054 14720
rect 22990 14660 22994 14716
rect 22994 14660 23050 14716
rect 23050 14660 23054 14716
rect 22990 14656 23054 14660
rect 23070 14716 23134 14720
rect 23070 14660 23074 14716
rect 23074 14660 23130 14716
rect 23130 14660 23134 14716
rect 23070 14656 23134 14660
rect 23150 14716 23214 14720
rect 23150 14660 23154 14716
rect 23154 14660 23210 14716
rect 23210 14660 23214 14716
rect 23150 14656 23214 14660
rect 23230 14716 23294 14720
rect 23230 14660 23234 14716
rect 23234 14660 23290 14716
rect 23290 14660 23294 14716
rect 23230 14656 23294 14660
rect 30879 14716 30943 14720
rect 30879 14660 30883 14716
rect 30883 14660 30939 14716
rect 30939 14660 30943 14716
rect 30879 14656 30943 14660
rect 30959 14716 31023 14720
rect 30959 14660 30963 14716
rect 30963 14660 31019 14716
rect 31019 14660 31023 14716
rect 30959 14656 31023 14660
rect 31039 14716 31103 14720
rect 31039 14660 31043 14716
rect 31043 14660 31099 14716
rect 31099 14660 31103 14716
rect 31039 14656 31103 14660
rect 31119 14716 31183 14720
rect 31119 14660 31123 14716
rect 31123 14660 31179 14716
rect 31179 14660 31183 14716
rect 31119 14656 31183 14660
rect 6552 14172 6616 14176
rect 6552 14116 6556 14172
rect 6556 14116 6612 14172
rect 6612 14116 6616 14172
rect 6552 14112 6616 14116
rect 6632 14172 6696 14176
rect 6632 14116 6636 14172
rect 6636 14116 6692 14172
rect 6692 14116 6696 14172
rect 6632 14112 6696 14116
rect 6712 14172 6776 14176
rect 6712 14116 6716 14172
rect 6716 14116 6772 14172
rect 6772 14116 6776 14172
rect 6712 14112 6776 14116
rect 6792 14172 6856 14176
rect 6792 14116 6796 14172
rect 6796 14116 6852 14172
rect 6852 14116 6856 14172
rect 6792 14112 6856 14116
rect 14441 14172 14505 14176
rect 14441 14116 14445 14172
rect 14445 14116 14501 14172
rect 14501 14116 14505 14172
rect 14441 14112 14505 14116
rect 14521 14172 14585 14176
rect 14521 14116 14525 14172
rect 14525 14116 14581 14172
rect 14581 14116 14585 14172
rect 14521 14112 14585 14116
rect 14601 14172 14665 14176
rect 14601 14116 14605 14172
rect 14605 14116 14661 14172
rect 14661 14116 14665 14172
rect 14601 14112 14665 14116
rect 14681 14172 14745 14176
rect 14681 14116 14685 14172
rect 14685 14116 14741 14172
rect 14741 14116 14745 14172
rect 14681 14112 14745 14116
rect 22330 14172 22394 14176
rect 22330 14116 22334 14172
rect 22334 14116 22390 14172
rect 22390 14116 22394 14172
rect 22330 14112 22394 14116
rect 22410 14172 22474 14176
rect 22410 14116 22414 14172
rect 22414 14116 22470 14172
rect 22470 14116 22474 14172
rect 22410 14112 22474 14116
rect 22490 14172 22554 14176
rect 22490 14116 22494 14172
rect 22494 14116 22550 14172
rect 22550 14116 22554 14172
rect 22490 14112 22554 14116
rect 22570 14172 22634 14176
rect 22570 14116 22574 14172
rect 22574 14116 22630 14172
rect 22630 14116 22634 14172
rect 22570 14112 22634 14116
rect 30219 14172 30283 14176
rect 30219 14116 30223 14172
rect 30223 14116 30279 14172
rect 30279 14116 30283 14172
rect 30219 14112 30283 14116
rect 30299 14172 30363 14176
rect 30299 14116 30303 14172
rect 30303 14116 30359 14172
rect 30359 14116 30363 14172
rect 30299 14112 30363 14116
rect 30379 14172 30443 14176
rect 30379 14116 30383 14172
rect 30383 14116 30439 14172
rect 30439 14116 30443 14172
rect 30379 14112 30443 14116
rect 30459 14172 30523 14176
rect 30459 14116 30463 14172
rect 30463 14116 30519 14172
rect 30519 14116 30523 14172
rect 30459 14112 30523 14116
rect 10916 13908 10980 13972
rect 17356 13772 17420 13836
rect 7212 13628 7276 13632
rect 7212 13572 7216 13628
rect 7216 13572 7272 13628
rect 7272 13572 7276 13628
rect 7212 13568 7276 13572
rect 7292 13628 7356 13632
rect 7292 13572 7296 13628
rect 7296 13572 7352 13628
rect 7352 13572 7356 13628
rect 7292 13568 7356 13572
rect 7372 13628 7436 13632
rect 7372 13572 7376 13628
rect 7376 13572 7432 13628
rect 7432 13572 7436 13628
rect 7372 13568 7436 13572
rect 7452 13628 7516 13632
rect 7452 13572 7456 13628
rect 7456 13572 7512 13628
rect 7512 13572 7516 13628
rect 7452 13568 7516 13572
rect 15101 13628 15165 13632
rect 15101 13572 15105 13628
rect 15105 13572 15161 13628
rect 15161 13572 15165 13628
rect 15101 13568 15165 13572
rect 15181 13628 15245 13632
rect 15181 13572 15185 13628
rect 15185 13572 15241 13628
rect 15241 13572 15245 13628
rect 15181 13568 15245 13572
rect 15261 13628 15325 13632
rect 15261 13572 15265 13628
rect 15265 13572 15321 13628
rect 15321 13572 15325 13628
rect 15261 13568 15325 13572
rect 15341 13628 15405 13632
rect 15341 13572 15345 13628
rect 15345 13572 15401 13628
rect 15401 13572 15405 13628
rect 15341 13568 15405 13572
rect 22990 13628 23054 13632
rect 22990 13572 22994 13628
rect 22994 13572 23050 13628
rect 23050 13572 23054 13628
rect 22990 13568 23054 13572
rect 23070 13628 23134 13632
rect 23070 13572 23074 13628
rect 23074 13572 23130 13628
rect 23130 13572 23134 13628
rect 23070 13568 23134 13572
rect 23150 13628 23214 13632
rect 23150 13572 23154 13628
rect 23154 13572 23210 13628
rect 23210 13572 23214 13628
rect 23150 13568 23214 13572
rect 23230 13628 23294 13632
rect 23230 13572 23234 13628
rect 23234 13572 23290 13628
rect 23290 13572 23294 13628
rect 23230 13568 23294 13572
rect 30879 13628 30943 13632
rect 30879 13572 30883 13628
rect 30883 13572 30939 13628
rect 30939 13572 30943 13628
rect 30879 13568 30943 13572
rect 30959 13628 31023 13632
rect 30959 13572 30963 13628
rect 30963 13572 31019 13628
rect 31019 13572 31023 13628
rect 30959 13568 31023 13572
rect 31039 13628 31103 13632
rect 31039 13572 31043 13628
rect 31043 13572 31099 13628
rect 31099 13572 31103 13628
rect 31039 13568 31103 13572
rect 31119 13628 31183 13632
rect 31119 13572 31123 13628
rect 31123 13572 31179 13628
rect 31179 13572 31183 13628
rect 31119 13568 31183 13572
rect 6552 13084 6616 13088
rect 6552 13028 6556 13084
rect 6556 13028 6612 13084
rect 6612 13028 6616 13084
rect 6552 13024 6616 13028
rect 6632 13084 6696 13088
rect 6632 13028 6636 13084
rect 6636 13028 6692 13084
rect 6692 13028 6696 13084
rect 6632 13024 6696 13028
rect 6712 13084 6776 13088
rect 6712 13028 6716 13084
rect 6716 13028 6772 13084
rect 6772 13028 6776 13084
rect 6712 13024 6776 13028
rect 6792 13084 6856 13088
rect 6792 13028 6796 13084
rect 6796 13028 6852 13084
rect 6852 13028 6856 13084
rect 6792 13024 6856 13028
rect 14441 13084 14505 13088
rect 14441 13028 14445 13084
rect 14445 13028 14501 13084
rect 14501 13028 14505 13084
rect 14441 13024 14505 13028
rect 14521 13084 14585 13088
rect 14521 13028 14525 13084
rect 14525 13028 14581 13084
rect 14581 13028 14585 13084
rect 14521 13024 14585 13028
rect 14601 13084 14665 13088
rect 14601 13028 14605 13084
rect 14605 13028 14661 13084
rect 14661 13028 14665 13084
rect 14601 13024 14665 13028
rect 14681 13084 14745 13088
rect 14681 13028 14685 13084
rect 14685 13028 14741 13084
rect 14741 13028 14745 13084
rect 14681 13024 14745 13028
rect 22330 13084 22394 13088
rect 22330 13028 22334 13084
rect 22334 13028 22390 13084
rect 22390 13028 22394 13084
rect 22330 13024 22394 13028
rect 22410 13084 22474 13088
rect 22410 13028 22414 13084
rect 22414 13028 22470 13084
rect 22470 13028 22474 13084
rect 22410 13024 22474 13028
rect 22490 13084 22554 13088
rect 22490 13028 22494 13084
rect 22494 13028 22550 13084
rect 22550 13028 22554 13084
rect 22490 13024 22554 13028
rect 22570 13084 22634 13088
rect 22570 13028 22574 13084
rect 22574 13028 22630 13084
rect 22630 13028 22634 13084
rect 22570 13024 22634 13028
rect 30219 13084 30283 13088
rect 30219 13028 30223 13084
rect 30223 13028 30279 13084
rect 30279 13028 30283 13084
rect 30219 13024 30283 13028
rect 30299 13084 30363 13088
rect 30299 13028 30303 13084
rect 30303 13028 30359 13084
rect 30359 13028 30363 13084
rect 30299 13024 30363 13028
rect 30379 13084 30443 13088
rect 30379 13028 30383 13084
rect 30383 13028 30439 13084
rect 30439 13028 30443 13084
rect 30379 13024 30443 13028
rect 30459 13084 30523 13088
rect 30459 13028 30463 13084
rect 30463 13028 30519 13084
rect 30519 13028 30523 13084
rect 30459 13024 30523 13028
rect 27844 12820 27908 12884
rect 7212 12540 7276 12544
rect 7212 12484 7216 12540
rect 7216 12484 7272 12540
rect 7272 12484 7276 12540
rect 7212 12480 7276 12484
rect 7292 12540 7356 12544
rect 7292 12484 7296 12540
rect 7296 12484 7352 12540
rect 7352 12484 7356 12540
rect 7292 12480 7356 12484
rect 7372 12540 7436 12544
rect 7372 12484 7376 12540
rect 7376 12484 7432 12540
rect 7432 12484 7436 12540
rect 7372 12480 7436 12484
rect 7452 12540 7516 12544
rect 7452 12484 7456 12540
rect 7456 12484 7512 12540
rect 7512 12484 7516 12540
rect 7452 12480 7516 12484
rect 15101 12540 15165 12544
rect 15101 12484 15105 12540
rect 15105 12484 15161 12540
rect 15161 12484 15165 12540
rect 15101 12480 15165 12484
rect 15181 12540 15245 12544
rect 15181 12484 15185 12540
rect 15185 12484 15241 12540
rect 15241 12484 15245 12540
rect 15181 12480 15245 12484
rect 15261 12540 15325 12544
rect 15261 12484 15265 12540
rect 15265 12484 15321 12540
rect 15321 12484 15325 12540
rect 15261 12480 15325 12484
rect 15341 12540 15405 12544
rect 15341 12484 15345 12540
rect 15345 12484 15401 12540
rect 15401 12484 15405 12540
rect 15341 12480 15405 12484
rect 22990 12540 23054 12544
rect 22990 12484 22994 12540
rect 22994 12484 23050 12540
rect 23050 12484 23054 12540
rect 22990 12480 23054 12484
rect 23070 12540 23134 12544
rect 23070 12484 23074 12540
rect 23074 12484 23130 12540
rect 23130 12484 23134 12540
rect 23070 12480 23134 12484
rect 23150 12540 23214 12544
rect 23150 12484 23154 12540
rect 23154 12484 23210 12540
rect 23210 12484 23214 12540
rect 23150 12480 23214 12484
rect 23230 12540 23294 12544
rect 23230 12484 23234 12540
rect 23234 12484 23290 12540
rect 23290 12484 23294 12540
rect 23230 12480 23294 12484
rect 30879 12540 30943 12544
rect 30879 12484 30883 12540
rect 30883 12484 30939 12540
rect 30939 12484 30943 12540
rect 30879 12480 30943 12484
rect 30959 12540 31023 12544
rect 30959 12484 30963 12540
rect 30963 12484 31019 12540
rect 31019 12484 31023 12540
rect 30959 12480 31023 12484
rect 31039 12540 31103 12544
rect 31039 12484 31043 12540
rect 31043 12484 31099 12540
rect 31099 12484 31103 12540
rect 31039 12480 31103 12484
rect 31119 12540 31183 12544
rect 31119 12484 31123 12540
rect 31123 12484 31179 12540
rect 31179 12484 31183 12540
rect 31119 12480 31183 12484
rect 6552 11996 6616 12000
rect 6552 11940 6556 11996
rect 6556 11940 6612 11996
rect 6612 11940 6616 11996
rect 6552 11936 6616 11940
rect 6632 11996 6696 12000
rect 6632 11940 6636 11996
rect 6636 11940 6692 11996
rect 6692 11940 6696 11996
rect 6632 11936 6696 11940
rect 6712 11996 6776 12000
rect 6712 11940 6716 11996
rect 6716 11940 6772 11996
rect 6772 11940 6776 11996
rect 6712 11936 6776 11940
rect 6792 11996 6856 12000
rect 6792 11940 6796 11996
rect 6796 11940 6852 11996
rect 6852 11940 6856 11996
rect 6792 11936 6856 11940
rect 14441 11996 14505 12000
rect 14441 11940 14445 11996
rect 14445 11940 14501 11996
rect 14501 11940 14505 11996
rect 14441 11936 14505 11940
rect 14521 11996 14585 12000
rect 14521 11940 14525 11996
rect 14525 11940 14581 11996
rect 14581 11940 14585 11996
rect 14521 11936 14585 11940
rect 14601 11996 14665 12000
rect 14601 11940 14605 11996
rect 14605 11940 14661 11996
rect 14661 11940 14665 11996
rect 14601 11936 14665 11940
rect 14681 11996 14745 12000
rect 14681 11940 14685 11996
rect 14685 11940 14741 11996
rect 14741 11940 14745 11996
rect 14681 11936 14745 11940
rect 22330 11996 22394 12000
rect 22330 11940 22334 11996
rect 22334 11940 22390 11996
rect 22390 11940 22394 11996
rect 22330 11936 22394 11940
rect 22410 11996 22474 12000
rect 22410 11940 22414 11996
rect 22414 11940 22470 11996
rect 22470 11940 22474 11996
rect 22410 11936 22474 11940
rect 22490 11996 22554 12000
rect 22490 11940 22494 11996
rect 22494 11940 22550 11996
rect 22550 11940 22554 11996
rect 22490 11936 22554 11940
rect 22570 11996 22634 12000
rect 22570 11940 22574 11996
rect 22574 11940 22630 11996
rect 22630 11940 22634 11996
rect 22570 11936 22634 11940
rect 30219 11996 30283 12000
rect 30219 11940 30223 11996
rect 30223 11940 30279 11996
rect 30279 11940 30283 11996
rect 30219 11936 30283 11940
rect 30299 11996 30363 12000
rect 30299 11940 30303 11996
rect 30303 11940 30359 11996
rect 30359 11940 30363 11996
rect 30299 11936 30363 11940
rect 30379 11996 30443 12000
rect 30379 11940 30383 11996
rect 30383 11940 30439 11996
rect 30439 11940 30443 11996
rect 30379 11936 30443 11940
rect 30459 11996 30523 12000
rect 30459 11940 30463 11996
rect 30463 11940 30519 11996
rect 30519 11940 30523 11996
rect 30459 11936 30523 11940
rect 22140 11656 22204 11660
rect 22140 11600 22190 11656
rect 22190 11600 22204 11656
rect 22140 11596 22204 11600
rect 7212 11452 7276 11456
rect 7212 11396 7216 11452
rect 7216 11396 7272 11452
rect 7272 11396 7276 11452
rect 7212 11392 7276 11396
rect 7292 11452 7356 11456
rect 7292 11396 7296 11452
rect 7296 11396 7352 11452
rect 7352 11396 7356 11452
rect 7292 11392 7356 11396
rect 7372 11452 7436 11456
rect 7372 11396 7376 11452
rect 7376 11396 7432 11452
rect 7432 11396 7436 11452
rect 7372 11392 7436 11396
rect 7452 11452 7516 11456
rect 7452 11396 7456 11452
rect 7456 11396 7512 11452
rect 7512 11396 7516 11452
rect 7452 11392 7516 11396
rect 15101 11452 15165 11456
rect 15101 11396 15105 11452
rect 15105 11396 15161 11452
rect 15161 11396 15165 11452
rect 15101 11392 15165 11396
rect 15181 11452 15245 11456
rect 15181 11396 15185 11452
rect 15185 11396 15241 11452
rect 15241 11396 15245 11452
rect 15181 11392 15245 11396
rect 15261 11452 15325 11456
rect 15261 11396 15265 11452
rect 15265 11396 15321 11452
rect 15321 11396 15325 11452
rect 15261 11392 15325 11396
rect 15341 11452 15405 11456
rect 15341 11396 15345 11452
rect 15345 11396 15401 11452
rect 15401 11396 15405 11452
rect 15341 11392 15405 11396
rect 22990 11452 23054 11456
rect 22990 11396 22994 11452
rect 22994 11396 23050 11452
rect 23050 11396 23054 11452
rect 22990 11392 23054 11396
rect 23070 11452 23134 11456
rect 23070 11396 23074 11452
rect 23074 11396 23130 11452
rect 23130 11396 23134 11452
rect 23070 11392 23134 11396
rect 23150 11452 23214 11456
rect 23150 11396 23154 11452
rect 23154 11396 23210 11452
rect 23210 11396 23214 11452
rect 23150 11392 23214 11396
rect 23230 11452 23294 11456
rect 23230 11396 23234 11452
rect 23234 11396 23290 11452
rect 23290 11396 23294 11452
rect 23230 11392 23294 11396
rect 30879 11452 30943 11456
rect 30879 11396 30883 11452
rect 30883 11396 30939 11452
rect 30939 11396 30943 11452
rect 30879 11392 30943 11396
rect 30959 11452 31023 11456
rect 30959 11396 30963 11452
rect 30963 11396 31019 11452
rect 31019 11396 31023 11452
rect 30959 11392 31023 11396
rect 31039 11452 31103 11456
rect 31039 11396 31043 11452
rect 31043 11396 31099 11452
rect 31099 11396 31103 11452
rect 31039 11392 31103 11396
rect 31119 11452 31183 11456
rect 31119 11396 31123 11452
rect 31123 11396 31179 11452
rect 31179 11396 31183 11452
rect 31119 11392 31183 11396
rect 19564 10916 19628 10980
rect 6552 10908 6616 10912
rect 6552 10852 6556 10908
rect 6556 10852 6612 10908
rect 6612 10852 6616 10908
rect 6552 10848 6616 10852
rect 6632 10908 6696 10912
rect 6632 10852 6636 10908
rect 6636 10852 6692 10908
rect 6692 10852 6696 10908
rect 6632 10848 6696 10852
rect 6712 10908 6776 10912
rect 6712 10852 6716 10908
rect 6716 10852 6772 10908
rect 6772 10852 6776 10908
rect 6712 10848 6776 10852
rect 6792 10908 6856 10912
rect 6792 10852 6796 10908
rect 6796 10852 6852 10908
rect 6852 10852 6856 10908
rect 6792 10848 6856 10852
rect 14441 10908 14505 10912
rect 14441 10852 14445 10908
rect 14445 10852 14501 10908
rect 14501 10852 14505 10908
rect 14441 10848 14505 10852
rect 14521 10908 14585 10912
rect 14521 10852 14525 10908
rect 14525 10852 14581 10908
rect 14581 10852 14585 10908
rect 14521 10848 14585 10852
rect 14601 10908 14665 10912
rect 14601 10852 14605 10908
rect 14605 10852 14661 10908
rect 14661 10852 14665 10908
rect 14601 10848 14665 10852
rect 14681 10908 14745 10912
rect 14681 10852 14685 10908
rect 14685 10852 14741 10908
rect 14741 10852 14745 10908
rect 14681 10848 14745 10852
rect 22330 10908 22394 10912
rect 22330 10852 22334 10908
rect 22334 10852 22390 10908
rect 22390 10852 22394 10908
rect 22330 10848 22394 10852
rect 22410 10908 22474 10912
rect 22410 10852 22414 10908
rect 22414 10852 22470 10908
rect 22470 10852 22474 10908
rect 22410 10848 22474 10852
rect 22490 10908 22554 10912
rect 22490 10852 22494 10908
rect 22494 10852 22550 10908
rect 22550 10852 22554 10908
rect 22490 10848 22554 10852
rect 22570 10908 22634 10912
rect 22570 10852 22574 10908
rect 22574 10852 22630 10908
rect 22630 10852 22634 10908
rect 22570 10848 22634 10852
rect 30219 10908 30283 10912
rect 30219 10852 30223 10908
rect 30223 10852 30279 10908
rect 30279 10852 30283 10908
rect 30219 10848 30283 10852
rect 30299 10908 30363 10912
rect 30299 10852 30303 10908
rect 30303 10852 30359 10908
rect 30359 10852 30363 10908
rect 30299 10848 30363 10852
rect 30379 10908 30443 10912
rect 30379 10852 30383 10908
rect 30383 10852 30439 10908
rect 30439 10852 30443 10908
rect 30379 10848 30443 10852
rect 30459 10908 30523 10912
rect 30459 10852 30463 10908
rect 30463 10852 30519 10908
rect 30519 10852 30523 10908
rect 30459 10848 30523 10852
rect 7212 10364 7276 10368
rect 7212 10308 7216 10364
rect 7216 10308 7272 10364
rect 7272 10308 7276 10364
rect 7212 10304 7276 10308
rect 7292 10364 7356 10368
rect 7292 10308 7296 10364
rect 7296 10308 7352 10364
rect 7352 10308 7356 10364
rect 7292 10304 7356 10308
rect 7372 10364 7436 10368
rect 7372 10308 7376 10364
rect 7376 10308 7432 10364
rect 7432 10308 7436 10364
rect 7372 10304 7436 10308
rect 7452 10364 7516 10368
rect 7452 10308 7456 10364
rect 7456 10308 7512 10364
rect 7512 10308 7516 10364
rect 7452 10304 7516 10308
rect 15101 10364 15165 10368
rect 15101 10308 15105 10364
rect 15105 10308 15161 10364
rect 15161 10308 15165 10364
rect 15101 10304 15165 10308
rect 15181 10364 15245 10368
rect 15181 10308 15185 10364
rect 15185 10308 15241 10364
rect 15241 10308 15245 10364
rect 15181 10304 15245 10308
rect 15261 10364 15325 10368
rect 15261 10308 15265 10364
rect 15265 10308 15321 10364
rect 15321 10308 15325 10364
rect 15261 10304 15325 10308
rect 15341 10364 15405 10368
rect 15341 10308 15345 10364
rect 15345 10308 15401 10364
rect 15401 10308 15405 10364
rect 15341 10304 15405 10308
rect 22990 10364 23054 10368
rect 22990 10308 22994 10364
rect 22994 10308 23050 10364
rect 23050 10308 23054 10364
rect 22990 10304 23054 10308
rect 23070 10364 23134 10368
rect 23070 10308 23074 10364
rect 23074 10308 23130 10364
rect 23130 10308 23134 10364
rect 23070 10304 23134 10308
rect 23150 10364 23214 10368
rect 23150 10308 23154 10364
rect 23154 10308 23210 10364
rect 23210 10308 23214 10364
rect 23150 10304 23214 10308
rect 23230 10364 23294 10368
rect 23230 10308 23234 10364
rect 23234 10308 23290 10364
rect 23290 10308 23294 10364
rect 23230 10304 23294 10308
rect 30879 10364 30943 10368
rect 30879 10308 30883 10364
rect 30883 10308 30939 10364
rect 30939 10308 30943 10364
rect 30879 10304 30943 10308
rect 30959 10364 31023 10368
rect 30959 10308 30963 10364
rect 30963 10308 31019 10364
rect 31019 10308 31023 10364
rect 30959 10304 31023 10308
rect 31039 10364 31103 10368
rect 31039 10308 31043 10364
rect 31043 10308 31099 10364
rect 31099 10308 31103 10364
rect 31039 10304 31103 10308
rect 31119 10364 31183 10368
rect 31119 10308 31123 10364
rect 31123 10308 31179 10364
rect 31179 10308 31183 10364
rect 31119 10304 31183 10308
rect 6552 9820 6616 9824
rect 6552 9764 6556 9820
rect 6556 9764 6612 9820
rect 6612 9764 6616 9820
rect 6552 9760 6616 9764
rect 6632 9820 6696 9824
rect 6632 9764 6636 9820
rect 6636 9764 6692 9820
rect 6692 9764 6696 9820
rect 6632 9760 6696 9764
rect 6712 9820 6776 9824
rect 6712 9764 6716 9820
rect 6716 9764 6772 9820
rect 6772 9764 6776 9820
rect 6712 9760 6776 9764
rect 6792 9820 6856 9824
rect 6792 9764 6796 9820
rect 6796 9764 6852 9820
rect 6852 9764 6856 9820
rect 6792 9760 6856 9764
rect 14441 9820 14505 9824
rect 14441 9764 14445 9820
rect 14445 9764 14501 9820
rect 14501 9764 14505 9820
rect 14441 9760 14505 9764
rect 14521 9820 14585 9824
rect 14521 9764 14525 9820
rect 14525 9764 14581 9820
rect 14581 9764 14585 9820
rect 14521 9760 14585 9764
rect 14601 9820 14665 9824
rect 14601 9764 14605 9820
rect 14605 9764 14661 9820
rect 14661 9764 14665 9820
rect 14601 9760 14665 9764
rect 14681 9820 14745 9824
rect 14681 9764 14685 9820
rect 14685 9764 14741 9820
rect 14741 9764 14745 9820
rect 14681 9760 14745 9764
rect 22330 9820 22394 9824
rect 22330 9764 22334 9820
rect 22334 9764 22390 9820
rect 22390 9764 22394 9820
rect 22330 9760 22394 9764
rect 22410 9820 22474 9824
rect 22410 9764 22414 9820
rect 22414 9764 22470 9820
rect 22470 9764 22474 9820
rect 22410 9760 22474 9764
rect 22490 9820 22554 9824
rect 22490 9764 22494 9820
rect 22494 9764 22550 9820
rect 22550 9764 22554 9820
rect 22490 9760 22554 9764
rect 22570 9820 22634 9824
rect 22570 9764 22574 9820
rect 22574 9764 22630 9820
rect 22630 9764 22634 9820
rect 22570 9760 22634 9764
rect 30219 9820 30283 9824
rect 30219 9764 30223 9820
rect 30223 9764 30279 9820
rect 30279 9764 30283 9820
rect 30219 9760 30283 9764
rect 30299 9820 30363 9824
rect 30299 9764 30303 9820
rect 30303 9764 30359 9820
rect 30359 9764 30363 9820
rect 30299 9760 30363 9764
rect 30379 9820 30443 9824
rect 30379 9764 30383 9820
rect 30383 9764 30439 9820
rect 30439 9764 30443 9820
rect 30379 9760 30443 9764
rect 30459 9820 30523 9824
rect 30459 9764 30463 9820
rect 30463 9764 30519 9820
rect 30519 9764 30523 9820
rect 30459 9760 30523 9764
rect 5764 9616 5828 9620
rect 5764 9560 5778 9616
rect 5778 9560 5828 9616
rect 5764 9556 5828 9560
rect 19196 9556 19260 9620
rect 21588 9420 21652 9484
rect 7212 9276 7276 9280
rect 7212 9220 7216 9276
rect 7216 9220 7272 9276
rect 7272 9220 7276 9276
rect 7212 9216 7276 9220
rect 7292 9276 7356 9280
rect 7292 9220 7296 9276
rect 7296 9220 7352 9276
rect 7352 9220 7356 9276
rect 7292 9216 7356 9220
rect 7372 9276 7436 9280
rect 7372 9220 7376 9276
rect 7376 9220 7432 9276
rect 7432 9220 7436 9276
rect 7372 9216 7436 9220
rect 7452 9276 7516 9280
rect 7452 9220 7456 9276
rect 7456 9220 7512 9276
rect 7512 9220 7516 9276
rect 7452 9216 7516 9220
rect 15101 9276 15165 9280
rect 15101 9220 15105 9276
rect 15105 9220 15161 9276
rect 15161 9220 15165 9276
rect 15101 9216 15165 9220
rect 15181 9276 15245 9280
rect 15181 9220 15185 9276
rect 15185 9220 15241 9276
rect 15241 9220 15245 9276
rect 15181 9216 15245 9220
rect 15261 9276 15325 9280
rect 15261 9220 15265 9276
rect 15265 9220 15321 9276
rect 15321 9220 15325 9276
rect 15261 9216 15325 9220
rect 15341 9276 15405 9280
rect 15341 9220 15345 9276
rect 15345 9220 15401 9276
rect 15401 9220 15405 9276
rect 15341 9216 15405 9220
rect 22990 9276 23054 9280
rect 22990 9220 22994 9276
rect 22994 9220 23050 9276
rect 23050 9220 23054 9276
rect 22990 9216 23054 9220
rect 23070 9276 23134 9280
rect 23070 9220 23074 9276
rect 23074 9220 23130 9276
rect 23130 9220 23134 9276
rect 23070 9216 23134 9220
rect 23150 9276 23214 9280
rect 23150 9220 23154 9276
rect 23154 9220 23210 9276
rect 23210 9220 23214 9276
rect 23150 9216 23214 9220
rect 23230 9276 23294 9280
rect 23230 9220 23234 9276
rect 23234 9220 23290 9276
rect 23290 9220 23294 9276
rect 23230 9216 23294 9220
rect 30879 9276 30943 9280
rect 30879 9220 30883 9276
rect 30883 9220 30939 9276
rect 30939 9220 30943 9276
rect 30879 9216 30943 9220
rect 30959 9276 31023 9280
rect 30959 9220 30963 9276
rect 30963 9220 31019 9276
rect 31019 9220 31023 9276
rect 30959 9216 31023 9220
rect 31039 9276 31103 9280
rect 31039 9220 31043 9276
rect 31043 9220 31099 9276
rect 31099 9220 31103 9276
rect 31039 9216 31103 9220
rect 31119 9276 31183 9280
rect 31119 9220 31123 9276
rect 31123 9220 31179 9276
rect 31179 9220 31183 9276
rect 31119 9216 31183 9220
rect 6552 8732 6616 8736
rect 6552 8676 6556 8732
rect 6556 8676 6612 8732
rect 6612 8676 6616 8732
rect 6552 8672 6616 8676
rect 6632 8732 6696 8736
rect 6632 8676 6636 8732
rect 6636 8676 6692 8732
rect 6692 8676 6696 8732
rect 6632 8672 6696 8676
rect 6712 8732 6776 8736
rect 6712 8676 6716 8732
rect 6716 8676 6772 8732
rect 6772 8676 6776 8732
rect 6712 8672 6776 8676
rect 6792 8732 6856 8736
rect 6792 8676 6796 8732
rect 6796 8676 6852 8732
rect 6852 8676 6856 8732
rect 6792 8672 6856 8676
rect 14441 8732 14505 8736
rect 14441 8676 14445 8732
rect 14445 8676 14501 8732
rect 14501 8676 14505 8732
rect 14441 8672 14505 8676
rect 14521 8732 14585 8736
rect 14521 8676 14525 8732
rect 14525 8676 14581 8732
rect 14581 8676 14585 8732
rect 14521 8672 14585 8676
rect 14601 8732 14665 8736
rect 14601 8676 14605 8732
rect 14605 8676 14661 8732
rect 14661 8676 14665 8732
rect 14601 8672 14665 8676
rect 14681 8732 14745 8736
rect 14681 8676 14685 8732
rect 14685 8676 14741 8732
rect 14741 8676 14745 8732
rect 14681 8672 14745 8676
rect 22330 8732 22394 8736
rect 22330 8676 22334 8732
rect 22334 8676 22390 8732
rect 22390 8676 22394 8732
rect 22330 8672 22394 8676
rect 22410 8732 22474 8736
rect 22410 8676 22414 8732
rect 22414 8676 22470 8732
rect 22470 8676 22474 8732
rect 22410 8672 22474 8676
rect 22490 8732 22554 8736
rect 22490 8676 22494 8732
rect 22494 8676 22550 8732
rect 22550 8676 22554 8732
rect 22490 8672 22554 8676
rect 22570 8732 22634 8736
rect 22570 8676 22574 8732
rect 22574 8676 22630 8732
rect 22630 8676 22634 8732
rect 22570 8672 22634 8676
rect 30219 8732 30283 8736
rect 30219 8676 30223 8732
rect 30223 8676 30279 8732
rect 30279 8676 30283 8732
rect 30219 8672 30283 8676
rect 30299 8732 30363 8736
rect 30299 8676 30303 8732
rect 30303 8676 30359 8732
rect 30359 8676 30363 8732
rect 30299 8672 30363 8676
rect 30379 8732 30443 8736
rect 30379 8676 30383 8732
rect 30383 8676 30439 8732
rect 30439 8676 30443 8732
rect 30379 8672 30443 8676
rect 30459 8732 30523 8736
rect 30459 8676 30463 8732
rect 30463 8676 30519 8732
rect 30519 8676 30523 8732
rect 30459 8672 30523 8676
rect 18828 8256 18892 8260
rect 18828 8200 18842 8256
rect 18842 8200 18892 8256
rect 18828 8196 18892 8200
rect 7212 8188 7276 8192
rect 7212 8132 7216 8188
rect 7216 8132 7272 8188
rect 7272 8132 7276 8188
rect 7212 8128 7276 8132
rect 7292 8188 7356 8192
rect 7292 8132 7296 8188
rect 7296 8132 7352 8188
rect 7352 8132 7356 8188
rect 7292 8128 7356 8132
rect 7372 8188 7436 8192
rect 7372 8132 7376 8188
rect 7376 8132 7432 8188
rect 7432 8132 7436 8188
rect 7372 8128 7436 8132
rect 7452 8188 7516 8192
rect 7452 8132 7456 8188
rect 7456 8132 7512 8188
rect 7512 8132 7516 8188
rect 7452 8128 7516 8132
rect 15101 8188 15165 8192
rect 15101 8132 15105 8188
rect 15105 8132 15161 8188
rect 15161 8132 15165 8188
rect 15101 8128 15165 8132
rect 15181 8188 15245 8192
rect 15181 8132 15185 8188
rect 15185 8132 15241 8188
rect 15241 8132 15245 8188
rect 15181 8128 15245 8132
rect 15261 8188 15325 8192
rect 15261 8132 15265 8188
rect 15265 8132 15321 8188
rect 15321 8132 15325 8188
rect 15261 8128 15325 8132
rect 15341 8188 15405 8192
rect 15341 8132 15345 8188
rect 15345 8132 15401 8188
rect 15401 8132 15405 8188
rect 15341 8128 15405 8132
rect 22990 8188 23054 8192
rect 22990 8132 22994 8188
rect 22994 8132 23050 8188
rect 23050 8132 23054 8188
rect 22990 8128 23054 8132
rect 23070 8188 23134 8192
rect 23070 8132 23074 8188
rect 23074 8132 23130 8188
rect 23130 8132 23134 8188
rect 23070 8128 23134 8132
rect 23150 8188 23214 8192
rect 23150 8132 23154 8188
rect 23154 8132 23210 8188
rect 23210 8132 23214 8188
rect 23150 8128 23214 8132
rect 23230 8188 23294 8192
rect 23230 8132 23234 8188
rect 23234 8132 23290 8188
rect 23290 8132 23294 8188
rect 23230 8128 23294 8132
rect 30879 8188 30943 8192
rect 30879 8132 30883 8188
rect 30883 8132 30939 8188
rect 30939 8132 30943 8188
rect 30879 8128 30943 8132
rect 30959 8188 31023 8192
rect 30959 8132 30963 8188
rect 30963 8132 31019 8188
rect 31019 8132 31023 8188
rect 30959 8128 31023 8132
rect 31039 8188 31103 8192
rect 31039 8132 31043 8188
rect 31043 8132 31099 8188
rect 31099 8132 31103 8188
rect 31039 8128 31103 8132
rect 31119 8188 31183 8192
rect 31119 8132 31123 8188
rect 31123 8132 31179 8188
rect 31179 8132 31183 8188
rect 31119 8128 31183 8132
rect 19380 8060 19444 8124
rect 26556 7924 26620 7988
rect 6552 7644 6616 7648
rect 6552 7588 6556 7644
rect 6556 7588 6612 7644
rect 6612 7588 6616 7644
rect 6552 7584 6616 7588
rect 6632 7644 6696 7648
rect 6632 7588 6636 7644
rect 6636 7588 6692 7644
rect 6692 7588 6696 7644
rect 6632 7584 6696 7588
rect 6712 7644 6776 7648
rect 6712 7588 6716 7644
rect 6716 7588 6772 7644
rect 6772 7588 6776 7644
rect 6712 7584 6776 7588
rect 6792 7644 6856 7648
rect 6792 7588 6796 7644
rect 6796 7588 6852 7644
rect 6852 7588 6856 7644
rect 6792 7584 6856 7588
rect 14441 7644 14505 7648
rect 14441 7588 14445 7644
rect 14445 7588 14501 7644
rect 14501 7588 14505 7644
rect 14441 7584 14505 7588
rect 14521 7644 14585 7648
rect 14521 7588 14525 7644
rect 14525 7588 14581 7644
rect 14581 7588 14585 7644
rect 14521 7584 14585 7588
rect 14601 7644 14665 7648
rect 14601 7588 14605 7644
rect 14605 7588 14661 7644
rect 14661 7588 14665 7644
rect 14601 7584 14665 7588
rect 14681 7644 14745 7648
rect 14681 7588 14685 7644
rect 14685 7588 14741 7644
rect 14741 7588 14745 7644
rect 14681 7584 14745 7588
rect 22330 7644 22394 7648
rect 22330 7588 22334 7644
rect 22334 7588 22390 7644
rect 22390 7588 22394 7644
rect 22330 7584 22394 7588
rect 22410 7644 22474 7648
rect 22410 7588 22414 7644
rect 22414 7588 22470 7644
rect 22470 7588 22474 7644
rect 22410 7584 22474 7588
rect 22490 7644 22554 7648
rect 22490 7588 22494 7644
rect 22494 7588 22550 7644
rect 22550 7588 22554 7644
rect 22490 7584 22554 7588
rect 22570 7644 22634 7648
rect 22570 7588 22574 7644
rect 22574 7588 22630 7644
rect 22630 7588 22634 7644
rect 22570 7584 22634 7588
rect 30219 7644 30283 7648
rect 30219 7588 30223 7644
rect 30223 7588 30279 7644
rect 30279 7588 30283 7644
rect 30219 7584 30283 7588
rect 30299 7644 30363 7648
rect 30299 7588 30303 7644
rect 30303 7588 30359 7644
rect 30359 7588 30363 7644
rect 30299 7584 30363 7588
rect 30379 7644 30443 7648
rect 30379 7588 30383 7644
rect 30383 7588 30439 7644
rect 30439 7588 30443 7644
rect 30379 7584 30443 7588
rect 30459 7644 30523 7648
rect 30459 7588 30463 7644
rect 30463 7588 30519 7644
rect 30519 7588 30523 7644
rect 30459 7584 30523 7588
rect 7212 7100 7276 7104
rect 7212 7044 7216 7100
rect 7216 7044 7272 7100
rect 7272 7044 7276 7100
rect 7212 7040 7276 7044
rect 7292 7100 7356 7104
rect 7292 7044 7296 7100
rect 7296 7044 7352 7100
rect 7352 7044 7356 7100
rect 7292 7040 7356 7044
rect 7372 7100 7436 7104
rect 7372 7044 7376 7100
rect 7376 7044 7432 7100
rect 7432 7044 7436 7100
rect 7372 7040 7436 7044
rect 7452 7100 7516 7104
rect 7452 7044 7456 7100
rect 7456 7044 7512 7100
rect 7512 7044 7516 7100
rect 7452 7040 7516 7044
rect 15101 7100 15165 7104
rect 15101 7044 15105 7100
rect 15105 7044 15161 7100
rect 15161 7044 15165 7100
rect 15101 7040 15165 7044
rect 15181 7100 15245 7104
rect 15181 7044 15185 7100
rect 15185 7044 15241 7100
rect 15241 7044 15245 7100
rect 15181 7040 15245 7044
rect 15261 7100 15325 7104
rect 15261 7044 15265 7100
rect 15265 7044 15321 7100
rect 15321 7044 15325 7100
rect 15261 7040 15325 7044
rect 15341 7100 15405 7104
rect 15341 7044 15345 7100
rect 15345 7044 15401 7100
rect 15401 7044 15405 7100
rect 15341 7040 15405 7044
rect 22990 7100 23054 7104
rect 22990 7044 22994 7100
rect 22994 7044 23050 7100
rect 23050 7044 23054 7100
rect 22990 7040 23054 7044
rect 23070 7100 23134 7104
rect 23070 7044 23074 7100
rect 23074 7044 23130 7100
rect 23130 7044 23134 7100
rect 23070 7040 23134 7044
rect 23150 7100 23214 7104
rect 23150 7044 23154 7100
rect 23154 7044 23210 7100
rect 23210 7044 23214 7100
rect 23150 7040 23214 7044
rect 23230 7100 23294 7104
rect 23230 7044 23234 7100
rect 23234 7044 23290 7100
rect 23290 7044 23294 7100
rect 23230 7040 23294 7044
rect 30879 7100 30943 7104
rect 30879 7044 30883 7100
rect 30883 7044 30939 7100
rect 30939 7044 30943 7100
rect 30879 7040 30943 7044
rect 30959 7100 31023 7104
rect 30959 7044 30963 7100
rect 30963 7044 31019 7100
rect 31019 7044 31023 7100
rect 30959 7040 31023 7044
rect 31039 7100 31103 7104
rect 31039 7044 31043 7100
rect 31043 7044 31099 7100
rect 31099 7044 31103 7100
rect 31039 7040 31103 7044
rect 31119 7100 31183 7104
rect 31119 7044 31123 7100
rect 31123 7044 31179 7100
rect 31179 7044 31183 7100
rect 31119 7040 31183 7044
rect 6552 6556 6616 6560
rect 6552 6500 6556 6556
rect 6556 6500 6612 6556
rect 6612 6500 6616 6556
rect 6552 6496 6616 6500
rect 6632 6556 6696 6560
rect 6632 6500 6636 6556
rect 6636 6500 6692 6556
rect 6692 6500 6696 6556
rect 6632 6496 6696 6500
rect 6712 6556 6776 6560
rect 6712 6500 6716 6556
rect 6716 6500 6772 6556
rect 6772 6500 6776 6556
rect 6712 6496 6776 6500
rect 6792 6556 6856 6560
rect 6792 6500 6796 6556
rect 6796 6500 6852 6556
rect 6852 6500 6856 6556
rect 6792 6496 6856 6500
rect 14441 6556 14505 6560
rect 14441 6500 14445 6556
rect 14445 6500 14501 6556
rect 14501 6500 14505 6556
rect 14441 6496 14505 6500
rect 14521 6556 14585 6560
rect 14521 6500 14525 6556
rect 14525 6500 14581 6556
rect 14581 6500 14585 6556
rect 14521 6496 14585 6500
rect 14601 6556 14665 6560
rect 14601 6500 14605 6556
rect 14605 6500 14661 6556
rect 14661 6500 14665 6556
rect 14601 6496 14665 6500
rect 14681 6556 14745 6560
rect 14681 6500 14685 6556
rect 14685 6500 14741 6556
rect 14741 6500 14745 6556
rect 14681 6496 14745 6500
rect 22330 6556 22394 6560
rect 22330 6500 22334 6556
rect 22334 6500 22390 6556
rect 22390 6500 22394 6556
rect 22330 6496 22394 6500
rect 22410 6556 22474 6560
rect 22410 6500 22414 6556
rect 22414 6500 22470 6556
rect 22470 6500 22474 6556
rect 22410 6496 22474 6500
rect 22490 6556 22554 6560
rect 22490 6500 22494 6556
rect 22494 6500 22550 6556
rect 22550 6500 22554 6556
rect 22490 6496 22554 6500
rect 22570 6556 22634 6560
rect 22570 6500 22574 6556
rect 22574 6500 22630 6556
rect 22630 6500 22634 6556
rect 22570 6496 22634 6500
rect 30219 6556 30283 6560
rect 30219 6500 30223 6556
rect 30223 6500 30279 6556
rect 30279 6500 30283 6556
rect 30219 6496 30283 6500
rect 30299 6556 30363 6560
rect 30299 6500 30303 6556
rect 30303 6500 30359 6556
rect 30359 6500 30363 6556
rect 30299 6496 30363 6500
rect 30379 6556 30443 6560
rect 30379 6500 30383 6556
rect 30383 6500 30439 6556
rect 30439 6500 30443 6556
rect 30379 6496 30443 6500
rect 30459 6556 30523 6560
rect 30459 6500 30463 6556
rect 30463 6500 30519 6556
rect 30519 6500 30523 6556
rect 30459 6496 30523 6500
rect 7212 6012 7276 6016
rect 7212 5956 7216 6012
rect 7216 5956 7272 6012
rect 7272 5956 7276 6012
rect 7212 5952 7276 5956
rect 7292 6012 7356 6016
rect 7292 5956 7296 6012
rect 7296 5956 7352 6012
rect 7352 5956 7356 6012
rect 7292 5952 7356 5956
rect 7372 6012 7436 6016
rect 7372 5956 7376 6012
rect 7376 5956 7432 6012
rect 7432 5956 7436 6012
rect 7372 5952 7436 5956
rect 7452 6012 7516 6016
rect 7452 5956 7456 6012
rect 7456 5956 7512 6012
rect 7512 5956 7516 6012
rect 7452 5952 7516 5956
rect 15101 6012 15165 6016
rect 15101 5956 15105 6012
rect 15105 5956 15161 6012
rect 15161 5956 15165 6012
rect 15101 5952 15165 5956
rect 15181 6012 15245 6016
rect 15181 5956 15185 6012
rect 15185 5956 15241 6012
rect 15241 5956 15245 6012
rect 15181 5952 15245 5956
rect 15261 6012 15325 6016
rect 15261 5956 15265 6012
rect 15265 5956 15321 6012
rect 15321 5956 15325 6012
rect 15261 5952 15325 5956
rect 15341 6012 15405 6016
rect 15341 5956 15345 6012
rect 15345 5956 15401 6012
rect 15401 5956 15405 6012
rect 15341 5952 15405 5956
rect 22990 6012 23054 6016
rect 22990 5956 22994 6012
rect 22994 5956 23050 6012
rect 23050 5956 23054 6012
rect 22990 5952 23054 5956
rect 23070 6012 23134 6016
rect 23070 5956 23074 6012
rect 23074 5956 23130 6012
rect 23130 5956 23134 6012
rect 23070 5952 23134 5956
rect 23150 6012 23214 6016
rect 23150 5956 23154 6012
rect 23154 5956 23210 6012
rect 23210 5956 23214 6012
rect 23150 5952 23214 5956
rect 23230 6012 23294 6016
rect 23230 5956 23234 6012
rect 23234 5956 23290 6012
rect 23290 5956 23294 6012
rect 23230 5952 23294 5956
rect 30879 6012 30943 6016
rect 30879 5956 30883 6012
rect 30883 5956 30939 6012
rect 30939 5956 30943 6012
rect 30879 5952 30943 5956
rect 30959 6012 31023 6016
rect 30959 5956 30963 6012
rect 30963 5956 31019 6012
rect 31019 5956 31023 6012
rect 30959 5952 31023 5956
rect 31039 6012 31103 6016
rect 31039 5956 31043 6012
rect 31043 5956 31099 6012
rect 31099 5956 31103 6012
rect 31039 5952 31103 5956
rect 31119 6012 31183 6016
rect 31119 5956 31123 6012
rect 31123 5956 31179 6012
rect 31179 5956 31183 6012
rect 31119 5952 31183 5956
rect 6552 5468 6616 5472
rect 6552 5412 6556 5468
rect 6556 5412 6612 5468
rect 6612 5412 6616 5468
rect 6552 5408 6616 5412
rect 6632 5468 6696 5472
rect 6632 5412 6636 5468
rect 6636 5412 6692 5468
rect 6692 5412 6696 5468
rect 6632 5408 6696 5412
rect 6712 5468 6776 5472
rect 6712 5412 6716 5468
rect 6716 5412 6772 5468
rect 6772 5412 6776 5468
rect 6712 5408 6776 5412
rect 6792 5468 6856 5472
rect 6792 5412 6796 5468
rect 6796 5412 6852 5468
rect 6852 5412 6856 5468
rect 6792 5408 6856 5412
rect 14441 5468 14505 5472
rect 14441 5412 14445 5468
rect 14445 5412 14501 5468
rect 14501 5412 14505 5468
rect 14441 5408 14505 5412
rect 14521 5468 14585 5472
rect 14521 5412 14525 5468
rect 14525 5412 14581 5468
rect 14581 5412 14585 5468
rect 14521 5408 14585 5412
rect 14601 5468 14665 5472
rect 14601 5412 14605 5468
rect 14605 5412 14661 5468
rect 14661 5412 14665 5468
rect 14601 5408 14665 5412
rect 14681 5468 14745 5472
rect 14681 5412 14685 5468
rect 14685 5412 14741 5468
rect 14741 5412 14745 5468
rect 14681 5408 14745 5412
rect 22330 5468 22394 5472
rect 22330 5412 22334 5468
rect 22334 5412 22390 5468
rect 22390 5412 22394 5468
rect 22330 5408 22394 5412
rect 22410 5468 22474 5472
rect 22410 5412 22414 5468
rect 22414 5412 22470 5468
rect 22470 5412 22474 5468
rect 22410 5408 22474 5412
rect 22490 5468 22554 5472
rect 22490 5412 22494 5468
rect 22494 5412 22550 5468
rect 22550 5412 22554 5468
rect 22490 5408 22554 5412
rect 22570 5468 22634 5472
rect 22570 5412 22574 5468
rect 22574 5412 22630 5468
rect 22630 5412 22634 5468
rect 22570 5408 22634 5412
rect 30219 5468 30283 5472
rect 30219 5412 30223 5468
rect 30223 5412 30279 5468
rect 30279 5412 30283 5468
rect 30219 5408 30283 5412
rect 30299 5468 30363 5472
rect 30299 5412 30303 5468
rect 30303 5412 30359 5468
rect 30359 5412 30363 5468
rect 30299 5408 30363 5412
rect 30379 5468 30443 5472
rect 30379 5412 30383 5468
rect 30383 5412 30439 5468
rect 30439 5412 30443 5468
rect 30379 5408 30443 5412
rect 30459 5468 30523 5472
rect 30459 5412 30463 5468
rect 30463 5412 30519 5468
rect 30519 5412 30523 5468
rect 30459 5408 30523 5412
rect 7212 4924 7276 4928
rect 7212 4868 7216 4924
rect 7216 4868 7272 4924
rect 7272 4868 7276 4924
rect 7212 4864 7276 4868
rect 7292 4924 7356 4928
rect 7292 4868 7296 4924
rect 7296 4868 7352 4924
rect 7352 4868 7356 4924
rect 7292 4864 7356 4868
rect 7372 4924 7436 4928
rect 7372 4868 7376 4924
rect 7376 4868 7432 4924
rect 7432 4868 7436 4924
rect 7372 4864 7436 4868
rect 7452 4924 7516 4928
rect 7452 4868 7456 4924
rect 7456 4868 7512 4924
rect 7512 4868 7516 4924
rect 7452 4864 7516 4868
rect 15101 4924 15165 4928
rect 15101 4868 15105 4924
rect 15105 4868 15161 4924
rect 15161 4868 15165 4924
rect 15101 4864 15165 4868
rect 15181 4924 15245 4928
rect 15181 4868 15185 4924
rect 15185 4868 15241 4924
rect 15241 4868 15245 4924
rect 15181 4864 15245 4868
rect 15261 4924 15325 4928
rect 15261 4868 15265 4924
rect 15265 4868 15321 4924
rect 15321 4868 15325 4924
rect 15261 4864 15325 4868
rect 15341 4924 15405 4928
rect 15341 4868 15345 4924
rect 15345 4868 15401 4924
rect 15401 4868 15405 4924
rect 15341 4864 15405 4868
rect 22990 4924 23054 4928
rect 22990 4868 22994 4924
rect 22994 4868 23050 4924
rect 23050 4868 23054 4924
rect 22990 4864 23054 4868
rect 23070 4924 23134 4928
rect 23070 4868 23074 4924
rect 23074 4868 23130 4924
rect 23130 4868 23134 4924
rect 23070 4864 23134 4868
rect 23150 4924 23214 4928
rect 23150 4868 23154 4924
rect 23154 4868 23210 4924
rect 23210 4868 23214 4924
rect 23150 4864 23214 4868
rect 23230 4924 23294 4928
rect 23230 4868 23234 4924
rect 23234 4868 23290 4924
rect 23290 4868 23294 4924
rect 23230 4864 23294 4868
rect 30879 4924 30943 4928
rect 30879 4868 30883 4924
rect 30883 4868 30939 4924
rect 30939 4868 30943 4924
rect 30879 4864 30943 4868
rect 30959 4924 31023 4928
rect 30959 4868 30963 4924
rect 30963 4868 31019 4924
rect 31019 4868 31023 4924
rect 30959 4864 31023 4868
rect 31039 4924 31103 4928
rect 31039 4868 31043 4924
rect 31043 4868 31099 4924
rect 31099 4868 31103 4924
rect 31039 4864 31103 4868
rect 31119 4924 31183 4928
rect 31119 4868 31123 4924
rect 31123 4868 31179 4924
rect 31179 4868 31183 4924
rect 31119 4864 31183 4868
rect 6552 4380 6616 4384
rect 6552 4324 6556 4380
rect 6556 4324 6612 4380
rect 6612 4324 6616 4380
rect 6552 4320 6616 4324
rect 6632 4380 6696 4384
rect 6632 4324 6636 4380
rect 6636 4324 6692 4380
rect 6692 4324 6696 4380
rect 6632 4320 6696 4324
rect 6712 4380 6776 4384
rect 6712 4324 6716 4380
rect 6716 4324 6772 4380
rect 6772 4324 6776 4380
rect 6712 4320 6776 4324
rect 6792 4380 6856 4384
rect 6792 4324 6796 4380
rect 6796 4324 6852 4380
rect 6852 4324 6856 4380
rect 6792 4320 6856 4324
rect 14441 4380 14505 4384
rect 14441 4324 14445 4380
rect 14445 4324 14501 4380
rect 14501 4324 14505 4380
rect 14441 4320 14505 4324
rect 14521 4380 14585 4384
rect 14521 4324 14525 4380
rect 14525 4324 14581 4380
rect 14581 4324 14585 4380
rect 14521 4320 14585 4324
rect 14601 4380 14665 4384
rect 14601 4324 14605 4380
rect 14605 4324 14661 4380
rect 14661 4324 14665 4380
rect 14601 4320 14665 4324
rect 14681 4380 14745 4384
rect 14681 4324 14685 4380
rect 14685 4324 14741 4380
rect 14741 4324 14745 4380
rect 14681 4320 14745 4324
rect 22330 4380 22394 4384
rect 22330 4324 22334 4380
rect 22334 4324 22390 4380
rect 22390 4324 22394 4380
rect 22330 4320 22394 4324
rect 22410 4380 22474 4384
rect 22410 4324 22414 4380
rect 22414 4324 22470 4380
rect 22470 4324 22474 4380
rect 22410 4320 22474 4324
rect 22490 4380 22554 4384
rect 22490 4324 22494 4380
rect 22494 4324 22550 4380
rect 22550 4324 22554 4380
rect 22490 4320 22554 4324
rect 22570 4380 22634 4384
rect 22570 4324 22574 4380
rect 22574 4324 22630 4380
rect 22630 4324 22634 4380
rect 22570 4320 22634 4324
rect 30219 4380 30283 4384
rect 30219 4324 30223 4380
rect 30223 4324 30279 4380
rect 30279 4324 30283 4380
rect 30219 4320 30283 4324
rect 30299 4380 30363 4384
rect 30299 4324 30303 4380
rect 30303 4324 30359 4380
rect 30359 4324 30363 4380
rect 30299 4320 30363 4324
rect 30379 4380 30443 4384
rect 30379 4324 30383 4380
rect 30383 4324 30439 4380
rect 30439 4324 30443 4380
rect 30379 4320 30443 4324
rect 30459 4380 30523 4384
rect 30459 4324 30463 4380
rect 30463 4324 30519 4380
rect 30519 4324 30523 4380
rect 30459 4320 30523 4324
rect 7212 3836 7276 3840
rect 7212 3780 7216 3836
rect 7216 3780 7272 3836
rect 7272 3780 7276 3836
rect 7212 3776 7276 3780
rect 7292 3836 7356 3840
rect 7292 3780 7296 3836
rect 7296 3780 7352 3836
rect 7352 3780 7356 3836
rect 7292 3776 7356 3780
rect 7372 3836 7436 3840
rect 7372 3780 7376 3836
rect 7376 3780 7432 3836
rect 7432 3780 7436 3836
rect 7372 3776 7436 3780
rect 7452 3836 7516 3840
rect 7452 3780 7456 3836
rect 7456 3780 7512 3836
rect 7512 3780 7516 3836
rect 7452 3776 7516 3780
rect 15101 3836 15165 3840
rect 15101 3780 15105 3836
rect 15105 3780 15161 3836
rect 15161 3780 15165 3836
rect 15101 3776 15165 3780
rect 15181 3836 15245 3840
rect 15181 3780 15185 3836
rect 15185 3780 15241 3836
rect 15241 3780 15245 3836
rect 15181 3776 15245 3780
rect 15261 3836 15325 3840
rect 15261 3780 15265 3836
rect 15265 3780 15321 3836
rect 15321 3780 15325 3836
rect 15261 3776 15325 3780
rect 15341 3836 15405 3840
rect 15341 3780 15345 3836
rect 15345 3780 15401 3836
rect 15401 3780 15405 3836
rect 15341 3776 15405 3780
rect 22990 3836 23054 3840
rect 22990 3780 22994 3836
rect 22994 3780 23050 3836
rect 23050 3780 23054 3836
rect 22990 3776 23054 3780
rect 23070 3836 23134 3840
rect 23070 3780 23074 3836
rect 23074 3780 23130 3836
rect 23130 3780 23134 3836
rect 23070 3776 23134 3780
rect 23150 3836 23214 3840
rect 23150 3780 23154 3836
rect 23154 3780 23210 3836
rect 23210 3780 23214 3836
rect 23150 3776 23214 3780
rect 23230 3836 23294 3840
rect 23230 3780 23234 3836
rect 23234 3780 23290 3836
rect 23290 3780 23294 3836
rect 23230 3776 23294 3780
rect 30879 3836 30943 3840
rect 30879 3780 30883 3836
rect 30883 3780 30939 3836
rect 30939 3780 30943 3836
rect 30879 3776 30943 3780
rect 30959 3836 31023 3840
rect 30959 3780 30963 3836
rect 30963 3780 31019 3836
rect 31019 3780 31023 3836
rect 30959 3776 31023 3780
rect 31039 3836 31103 3840
rect 31039 3780 31043 3836
rect 31043 3780 31099 3836
rect 31099 3780 31103 3836
rect 31039 3776 31103 3780
rect 31119 3836 31183 3840
rect 31119 3780 31123 3836
rect 31123 3780 31179 3836
rect 31179 3780 31183 3836
rect 31119 3776 31183 3780
rect 6552 3292 6616 3296
rect 6552 3236 6556 3292
rect 6556 3236 6612 3292
rect 6612 3236 6616 3292
rect 6552 3232 6616 3236
rect 6632 3292 6696 3296
rect 6632 3236 6636 3292
rect 6636 3236 6692 3292
rect 6692 3236 6696 3292
rect 6632 3232 6696 3236
rect 6712 3292 6776 3296
rect 6712 3236 6716 3292
rect 6716 3236 6772 3292
rect 6772 3236 6776 3292
rect 6712 3232 6776 3236
rect 6792 3292 6856 3296
rect 6792 3236 6796 3292
rect 6796 3236 6852 3292
rect 6852 3236 6856 3292
rect 6792 3232 6856 3236
rect 14441 3292 14505 3296
rect 14441 3236 14445 3292
rect 14445 3236 14501 3292
rect 14501 3236 14505 3292
rect 14441 3232 14505 3236
rect 14521 3292 14585 3296
rect 14521 3236 14525 3292
rect 14525 3236 14581 3292
rect 14581 3236 14585 3292
rect 14521 3232 14585 3236
rect 14601 3292 14665 3296
rect 14601 3236 14605 3292
rect 14605 3236 14661 3292
rect 14661 3236 14665 3292
rect 14601 3232 14665 3236
rect 14681 3292 14745 3296
rect 14681 3236 14685 3292
rect 14685 3236 14741 3292
rect 14741 3236 14745 3292
rect 14681 3232 14745 3236
rect 22330 3292 22394 3296
rect 22330 3236 22334 3292
rect 22334 3236 22390 3292
rect 22390 3236 22394 3292
rect 22330 3232 22394 3236
rect 22410 3292 22474 3296
rect 22410 3236 22414 3292
rect 22414 3236 22470 3292
rect 22470 3236 22474 3292
rect 22410 3232 22474 3236
rect 22490 3292 22554 3296
rect 22490 3236 22494 3292
rect 22494 3236 22550 3292
rect 22550 3236 22554 3292
rect 22490 3232 22554 3236
rect 22570 3292 22634 3296
rect 22570 3236 22574 3292
rect 22574 3236 22630 3292
rect 22630 3236 22634 3292
rect 22570 3232 22634 3236
rect 30219 3292 30283 3296
rect 30219 3236 30223 3292
rect 30223 3236 30279 3292
rect 30279 3236 30283 3292
rect 30219 3232 30283 3236
rect 30299 3292 30363 3296
rect 30299 3236 30303 3292
rect 30303 3236 30359 3292
rect 30359 3236 30363 3292
rect 30299 3232 30363 3236
rect 30379 3292 30443 3296
rect 30379 3236 30383 3292
rect 30383 3236 30439 3292
rect 30439 3236 30443 3292
rect 30379 3232 30443 3236
rect 30459 3292 30523 3296
rect 30459 3236 30463 3292
rect 30463 3236 30519 3292
rect 30519 3236 30523 3292
rect 30459 3232 30523 3236
rect 15700 3028 15764 3092
rect 7212 2748 7276 2752
rect 7212 2692 7216 2748
rect 7216 2692 7272 2748
rect 7272 2692 7276 2748
rect 7212 2688 7276 2692
rect 7292 2748 7356 2752
rect 7292 2692 7296 2748
rect 7296 2692 7352 2748
rect 7352 2692 7356 2748
rect 7292 2688 7356 2692
rect 7372 2748 7436 2752
rect 7372 2692 7376 2748
rect 7376 2692 7432 2748
rect 7432 2692 7436 2748
rect 7372 2688 7436 2692
rect 7452 2748 7516 2752
rect 7452 2692 7456 2748
rect 7456 2692 7512 2748
rect 7512 2692 7516 2748
rect 7452 2688 7516 2692
rect 15101 2748 15165 2752
rect 15101 2692 15105 2748
rect 15105 2692 15161 2748
rect 15161 2692 15165 2748
rect 15101 2688 15165 2692
rect 15181 2748 15245 2752
rect 15181 2692 15185 2748
rect 15185 2692 15241 2748
rect 15241 2692 15245 2748
rect 15181 2688 15245 2692
rect 15261 2748 15325 2752
rect 15261 2692 15265 2748
rect 15265 2692 15321 2748
rect 15321 2692 15325 2748
rect 15261 2688 15325 2692
rect 15341 2748 15405 2752
rect 15341 2692 15345 2748
rect 15345 2692 15401 2748
rect 15401 2692 15405 2748
rect 15341 2688 15405 2692
rect 22990 2748 23054 2752
rect 22990 2692 22994 2748
rect 22994 2692 23050 2748
rect 23050 2692 23054 2748
rect 22990 2688 23054 2692
rect 23070 2748 23134 2752
rect 23070 2692 23074 2748
rect 23074 2692 23130 2748
rect 23130 2692 23134 2748
rect 23070 2688 23134 2692
rect 23150 2748 23214 2752
rect 23150 2692 23154 2748
rect 23154 2692 23210 2748
rect 23210 2692 23214 2748
rect 23150 2688 23214 2692
rect 23230 2748 23294 2752
rect 23230 2692 23234 2748
rect 23234 2692 23290 2748
rect 23290 2692 23294 2748
rect 23230 2688 23294 2692
rect 30879 2748 30943 2752
rect 30879 2692 30883 2748
rect 30883 2692 30939 2748
rect 30939 2692 30943 2748
rect 30879 2688 30943 2692
rect 30959 2748 31023 2752
rect 30959 2692 30963 2748
rect 30963 2692 31019 2748
rect 31019 2692 31023 2748
rect 30959 2688 31023 2692
rect 31039 2748 31103 2752
rect 31039 2692 31043 2748
rect 31043 2692 31099 2748
rect 31099 2692 31103 2748
rect 31039 2688 31103 2692
rect 31119 2748 31183 2752
rect 31119 2692 31123 2748
rect 31123 2692 31179 2748
rect 31179 2692 31183 2748
rect 31119 2688 31183 2692
<< metal4 >>
rect 6544 33760 6864 34320
rect 6544 33696 6552 33760
rect 6616 33696 6632 33760
rect 6696 33696 6712 33760
rect 6776 33696 6792 33760
rect 6856 33696 6864 33760
rect 6544 32672 6864 33696
rect 6544 32608 6552 32672
rect 6616 32608 6632 32672
rect 6696 32608 6712 32672
rect 6776 32608 6792 32672
rect 6856 32608 6864 32672
rect 6544 31584 6864 32608
rect 6544 31520 6552 31584
rect 6616 31520 6632 31584
rect 6696 31520 6712 31584
rect 6776 31520 6792 31584
rect 6856 31520 6864 31584
rect 6544 30496 6864 31520
rect 6544 30432 6552 30496
rect 6616 30432 6632 30496
rect 6696 30432 6712 30496
rect 6776 30432 6792 30496
rect 6856 30432 6864 30496
rect 6544 29408 6864 30432
rect 6544 29344 6552 29408
rect 6616 29344 6632 29408
rect 6696 29344 6712 29408
rect 6776 29344 6792 29408
rect 6856 29344 6864 29408
rect 6544 28320 6864 29344
rect 6544 28256 6552 28320
rect 6616 28256 6632 28320
rect 6696 28256 6712 28320
rect 6776 28256 6792 28320
rect 6856 28256 6864 28320
rect 6544 27232 6864 28256
rect 6544 27168 6552 27232
rect 6616 27168 6632 27232
rect 6696 27168 6712 27232
rect 6776 27168 6792 27232
rect 6856 27168 6864 27232
rect 6544 26144 6864 27168
rect 6544 26080 6552 26144
rect 6616 26080 6632 26144
rect 6696 26080 6712 26144
rect 6776 26080 6792 26144
rect 6856 26080 6864 26144
rect 6544 25056 6864 26080
rect 6544 24992 6552 25056
rect 6616 24992 6632 25056
rect 6696 24992 6712 25056
rect 6776 24992 6792 25056
rect 6856 24992 6864 25056
rect 5579 24988 5645 24989
rect 5579 24924 5580 24988
rect 5644 24924 5645 24988
rect 5579 24923 5645 24924
rect 5582 15197 5642 24923
rect 6544 23968 6864 24992
rect 6544 23904 6552 23968
rect 6616 23904 6632 23968
rect 6696 23904 6712 23968
rect 6776 23904 6792 23968
rect 6856 23904 6864 23968
rect 6131 23628 6197 23629
rect 6131 23564 6132 23628
rect 6196 23564 6197 23628
rect 6131 23563 6197 23564
rect 5763 23492 5829 23493
rect 5763 23428 5764 23492
rect 5828 23428 5829 23492
rect 5763 23427 5829 23428
rect 5579 15196 5645 15197
rect 5579 15132 5580 15196
rect 5644 15132 5645 15196
rect 5579 15131 5645 15132
rect 5766 9621 5826 23427
rect 6134 20229 6194 23563
rect 6544 22880 6864 23904
rect 6544 22816 6552 22880
rect 6616 22816 6632 22880
rect 6696 22816 6712 22880
rect 6776 22816 6792 22880
rect 6856 22816 6864 22880
rect 6544 21792 6864 22816
rect 6544 21728 6552 21792
rect 6616 21728 6632 21792
rect 6696 21728 6712 21792
rect 6776 21728 6792 21792
rect 6856 21728 6864 21792
rect 6544 20704 6864 21728
rect 6544 20640 6552 20704
rect 6616 20640 6632 20704
rect 6696 20640 6712 20704
rect 6776 20640 6792 20704
rect 6856 20640 6864 20704
rect 6131 20228 6197 20229
rect 6131 20164 6132 20228
rect 6196 20164 6197 20228
rect 6131 20163 6197 20164
rect 6544 19616 6864 20640
rect 6544 19552 6552 19616
rect 6616 19552 6632 19616
rect 6696 19552 6712 19616
rect 6776 19552 6792 19616
rect 6856 19552 6864 19616
rect 6544 18528 6864 19552
rect 6544 18464 6552 18528
rect 6616 18464 6632 18528
rect 6696 18464 6712 18528
rect 6776 18464 6792 18528
rect 6856 18464 6864 18528
rect 6544 17440 6864 18464
rect 6544 17376 6552 17440
rect 6616 17376 6632 17440
rect 6696 17376 6712 17440
rect 6776 17376 6792 17440
rect 6856 17376 6864 17440
rect 6544 16352 6864 17376
rect 6544 16288 6552 16352
rect 6616 16288 6632 16352
rect 6696 16288 6712 16352
rect 6776 16288 6792 16352
rect 6856 16288 6864 16352
rect 6544 15264 6864 16288
rect 6544 15200 6552 15264
rect 6616 15200 6632 15264
rect 6696 15200 6712 15264
rect 6776 15200 6792 15264
rect 6856 15200 6864 15264
rect 6544 14176 6864 15200
rect 6544 14112 6552 14176
rect 6616 14112 6632 14176
rect 6696 14112 6712 14176
rect 6776 14112 6792 14176
rect 6856 14112 6864 14176
rect 6544 13088 6864 14112
rect 6544 13024 6552 13088
rect 6616 13024 6632 13088
rect 6696 13024 6712 13088
rect 6776 13024 6792 13088
rect 6856 13024 6864 13088
rect 6544 12000 6864 13024
rect 6544 11936 6552 12000
rect 6616 11936 6632 12000
rect 6696 11936 6712 12000
rect 6776 11936 6792 12000
rect 6856 11936 6864 12000
rect 6544 10912 6864 11936
rect 6544 10848 6552 10912
rect 6616 10848 6632 10912
rect 6696 10848 6712 10912
rect 6776 10848 6792 10912
rect 6856 10848 6864 10912
rect 6544 9824 6864 10848
rect 6544 9760 6552 9824
rect 6616 9760 6632 9824
rect 6696 9760 6712 9824
rect 6776 9760 6792 9824
rect 6856 9760 6864 9824
rect 5763 9620 5829 9621
rect 5763 9556 5764 9620
rect 5828 9556 5829 9620
rect 5763 9555 5829 9556
rect 6544 8736 6864 9760
rect 6544 8672 6552 8736
rect 6616 8672 6632 8736
rect 6696 8672 6712 8736
rect 6776 8672 6792 8736
rect 6856 8672 6864 8736
rect 6544 7648 6864 8672
rect 6544 7584 6552 7648
rect 6616 7584 6632 7648
rect 6696 7584 6712 7648
rect 6776 7584 6792 7648
rect 6856 7584 6864 7648
rect 6544 6560 6864 7584
rect 6544 6496 6552 6560
rect 6616 6496 6632 6560
rect 6696 6496 6712 6560
rect 6776 6496 6792 6560
rect 6856 6496 6864 6560
rect 6544 5472 6864 6496
rect 6544 5408 6552 5472
rect 6616 5408 6632 5472
rect 6696 5408 6712 5472
rect 6776 5408 6792 5472
rect 6856 5408 6864 5472
rect 6544 4384 6864 5408
rect 6544 4320 6552 4384
rect 6616 4320 6632 4384
rect 6696 4320 6712 4384
rect 6776 4320 6792 4384
rect 6856 4320 6864 4384
rect 6544 3296 6864 4320
rect 6544 3232 6552 3296
rect 6616 3232 6632 3296
rect 6696 3232 6712 3296
rect 6776 3232 6792 3296
rect 6856 3232 6864 3296
rect 6544 2672 6864 3232
rect 7204 34304 7524 34320
rect 7204 34240 7212 34304
rect 7276 34240 7292 34304
rect 7356 34240 7372 34304
rect 7436 34240 7452 34304
rect 7516 34240 7524 34304
rect 7204 33216 7524 34240
rect 14433 33760 14753 34320
rect 14433 33696 14441 33760
rect 14505 33696 14521 33760
rect 14585 33696 14601 33760
rect 14665 33696 14681 33760
rect 14745 33696 14753 33760
rect 10915 33284 10981 33285
rect 10915 33220 10916 33284
rect 10980 33220 10981 33284
rect 10915 33219 10981 33220
rect 7204 33152 7212 33216
rect 7276 33152 7292 33216
rect 7356 33152 7372 33216
rect 7436 33152 7452 33216
rect 7516 33152 7524 33216
rect 7204 32128 7524 33152
rect 7204 32064 7212 32128
rect 7276 32064 7292 32128
rect 7356 32064 7372 32128
rect 7436 32064 7452 32128
rect 7516 32064 7524 32128
rect 7204 31040 7524 32064
rect 7204 30976 7212 31040
rect 7276 30976 7292 31040
rect 7356 30976 7372 31040
rect 7436 30976 7452 31040
rect 7516 30976 7524 31040
rect 7204 29952 7524 30976
rect 7204 29888 7212 29952
rect 7276 29888 7292 29952
rect 7356 29888 7372 29952
rect 7436 29888 7452 29952
rect 7516 29888 7524 29952
rect 7204 28864 7524 29888
rect 7204 28800 7212 28864
rect 7276 28800 7292 28864
rect 7356 28800 7372 28864
rect 7436 28800 7452 28864
rect 7516 28800 7524 28864
rect 7204 27776 7524 28800
rect 7204 27712 7212 27776
rect 7276 27712 7292 27776
rect 7356 27712 7372 27776
rect 7436 27712 7452 27776
rect 7516 27712 7524 27776
rect 7204 26688 7524 27712
rect 7204 26624 7212 26688
rect 7276 26624 7292 26688
rect 7356 26624 7372 26688
rect 7436 26624 7452 26688
rect 7516 26624 7524 26688
rect 7204 25600 7524 26624
rect 7204 25536 7212 25600
rect 7276 25536 7292 25600
rect 7356 25536 7372 25600
rect 7436 25536 7452 25600
rect 7516 25536 7524 25600
rect 7204 24512 7524 25536
rect 7204 24448 7212 24512
rect 7276 24448 7292 24512
rect 7356 24448 7372 24512
rect 7436 24448 7452 24512
rect 7516 24448 7524 24512
rect 7204 23424 7524 24448
rect 7204 23360 7212 23424
rect 7276 23360 7292 23424
rect 7356 23360 7372 23424
rect 7436 23360 7452 23424
rect 7516 23360 7524 23424
rect 7204 22336 7524 23360
rect 7204 22272 7212 22336
rect 7276 22272 7292 22336
rect 7356 22272 7372 22336
rect 7436 22272 7452 22336
rect 7516 22272 7524 22336
rect 7204 21248 7524 22272
rect 7204 21184 7212 21248
rect 7276 21184 7292 21248
rect 7356 21184 7372 21248
rect 7436 21184 7452 21248
rect 7516 21184 7524 21248
rect 7204 20160 7524 21184
rect 7204 20096 7212 20160
rect 7276 20096 7292 20160
rect 7356 20096 7372 20160
rect 7436 20096 7452 20160
rect 7516 20096 7524 20160
rect 7204 19072 7524 20096
rect 7204 19008 7212 19072
rect 7276 19008 7292 19072
rect 7356 19008 7372 19072
rect 7436 19008 7452 19072
rect 7516 19008 7524 19072
rect 7204 17984 7524 19008
rect 7204 17920 7212 17984
rect 7276 17920 7292 17984
rect 7356 17920 7372 17984
rect 7436 17920 7452 17984
rect 7516 17920 7524 17984
rect 7204 16896 7524 17920
rect 7204 16832 7212 16896
rect 7276 16832 7292 16896
rect 7356 16832 7372 16896
rect 7436 16832 7452 16896
rect 7516 16832 7524 16896
rect 7204 15808 7524 16832
rect 7204 15744 7212 15808
rect 7276 15744 7292 15808
rect 7356 15744 7372 15808
rect 7436 15744 7452 15808
rect 7516 15744 7524 15808
rect 7204 14720 7524 15744
rect 7204 14656 7212 14720
rect 7276 14656 7292 14720
rect 7356 14656 7372 14720
rect 7436 14656 7452 14720
rect 7516 14656 7524 14720
rect 7204 13632 7524 14656
rect 10918 13973 10978 33219
rect 12203 33148 12269 33149
rect 12203 33084 12204 33148
rect 12268 33084 12269 33148
rect 12203 33083 12269 33084
rect 11835 21724 11901 21725
rect 11835 21660 11836 21724
rect 11900 21660 11901 21724
rect 11835 21659 11901 21660
rect 11838 20501 11898 21659
rect 12206 20501 12266 33083
rect 14433 32672 14753 33696
rect 14433 32608 14441 32672
rect 14505 32608 14521 32672
rect 14585 32608 14601 32672
rect 14665 32608 14681 32672
rect 14745 32608 14753 32672
rect 14433 31584 14753 32608
rect 14433 31520 14441 31584
rect 14505 31520 14521 31584
rect 14585 31520 14601 31584
rect 14665 31520 14681 31584
rect 14745 31520 14753 31584
rect 14433 30496 14753 31520
rect 14433 30432 14441 30496
rect 14505 30432 14521 30496
rect 14585 30432 14601 30496
rect 14665 30432 14681 30496
rect 14745 30432 14753 30496
rect 14433 29408 14753 30432
rect 14433 29344 14441 29408
rect 14505 29344 14521 29408
rect 14585 29344 14601 29408
rect 14665 29344 14681 29408
rect 14745 29344 14753 29408
rect 14433 28320 14753 29344
rect 14433 28256 14441 28320
rect 14505 28256 14521 28320
rect 14585 28256 14601 28320
rect 14665 28256 14681 28320
rect 14745 28256 14753 28320
rect 14433 27232 14753 28256
rect 14433 27168 14441 27232
rect 14505 27168 14521 27232
rect 14585 27168 14601 27232
rect 14665 27168 14681 27232
rect 14745 27168 14753 27232
rect 14433 26144 14753 27168
rect 14433 26080 14441 26144
rect 14505 26080 14521 26144
rect 14585 26080 14601 26144
rect 14665 26080 14681 26144
rect 14745 26080 14753 26144
rect 14433 25056 14753 26080
rect 14433 24992 14441 25056
rect 14505 24992 14521 25056
rect 14585 24992 14601 25056
rect 14665 24992 14681 25056
rect 14745 24992 14753 25056
rect 14433 23968 14753 24992
rect 14433 23904 14441 23968
rect 14505 23904 14521 23968
rect 14585 23904 14601 23968
rect 14665 23904 14681 23968
rect 14745 23904 14753 23968
rect 14433 22880 14753 23904
rect 14433 22816 14441 22880
rect 14505 22816 14521 22880
rect 14585 22816 14601 22880
rect 14665 22816 14681 22880
rect 14745 22816 14753 22880
rect 14433 21792 14753 22816
rect 14433 21728 14441 21792
rect 14505 21728 14521 21792
rect 14585 21728 14601 21792
rect 14665 21728 14681 21792
rect 14745 21728 14753 21792
rect 14433 20704 14753 21728
rect 14433 20640 14441 20704
rect 14505 20640 14521 20704
rect 14585 20640 14601 20704
rect 14665 20640 14681 20704
rect 14745 20640 14753 20704
rect 11835 20500 11901 20501
rect 11835 20436 11836 20500
rect 11900 20436 11901 20500
rect 11835 20435 11901 20436
rect 12203 20500 12269 20501
rect 12203 20436 12204 20500
rect 12268 20436 12269 20500
rect 12203 20435 12269 20436
rect 14433 19616 14753 20640
rect 14433 19552 14441 19616
rect 14505 19552 14521 19616
rect 14585 19552 14601 19616
rect 14665 19552 14681 19616
rect 14745 19552 14753 19616
rect 14433 18528 14753 19552
rect 14433 18464 14441 18528
rect 14505 18464 14521 18528
rect 14585 18464 14601 18528
rect 14665 18464 14681 18528
rect 14745 18464 14753 18528
rect 14433 17440 14753 18464
rect 14433 17376 14441 17440
rect 14505 17376 14521 17440
rect 14585 17376 14601 17440
rect 14665 17376 14681 17440
rect 14745 17376 14753 17440
rect 14433 16352 14753 17376
rect 14433 16288 14441 16352
rect 14505 16288 14521 16352
rect 14585 16288 14601 16352
rect 14665 16288 14681 16352
rect 14745 16288 14753 16352
rect 14433 15264 14753 16288
rect 14433 15200 14441 15264
rect 14505 15200 14521 15264
rect 14585 15200 14601 15264
rect 14665 15200 14681 15264
rect 14745 15200 14753 15264
rect 14433 14176 14753 15200
rect 14433 14112 14441 14176
rect 14505 14112 14521 14176
rect 14585 14112 14601 14176
rect 14665 14112 14681 14176
rect 14745 14112 14753 14176
rect 10915 13972 10981 13973
rect 10915 13908 10916 13972
rect 10980 13908 10981 13972
rect 10915 13907 10981 13908
rect 7204 13568 7212 13632
rect 7276 13568 7292 13632
rect 7356 13568 7372 13632
rect 7436 13568 7452 13632
rect 7516 13568 7524 13632
rect 7204 12544 7524 13568
rect 7204 12480 7212 12544
rect 7276 12480 7292 12544
rect 7356 12480 7372 12544
rect 7436 12480 7452 12544
rect 7516 12480 7524 12544
rect 7204 11456 7524 12480
rect 7204 11392 7212 11456
rect 7276 11392 7292 11456
rect 7356 11392 7372 11456
rect 7436 11392 7452 11456
rect 7516 11392 7524 11456
rect 7204 10368 7524 11392
rect 7204 10304 7212 10368
rect 7276 10304 7292 10368
rect 7356 10304 7372 10368
rect 7436 10304 7452 10368
rect 7516 10304 7524 10368
rect 7204 9280 7524 10304
rect 7204 9216 7212 9280
rect 7276 9216 7292 9280
rect 7356 9216 7372 9280
rect 7436 9216 7452 9280
rect 7516 9216 7524 9280
rect 7204 8192 7524 9216
rect 7204 8128 7212 8192
rect 7276 8128 7292 8192
rect 7356 8128 7372 8192
rect 7436 8128 7452 8192
rect 7516 8128 7524 8192
rect 7204 7104 7524 8128
rect 7204 7040 7212 7104
rect 7276 7040 7292 7104
rect 7356 7040 7372 7104
rect 7436 7040 7452 7104
rect 7516 7040 7524 7104
rect 7204 6016 7524 7040
rect 7204 5952 7212 6016
rect 7276 5952 7292 6016
rect 7356 5952 7372 6016
rect 7436 5952 7452 6016
rect 7516 5952 7524 6016
rect 7204 4928 7524 5952
rect 7204 4864 7212 4928
rect 7276 4864 7292 4928
rect 7356 4864 7372 4928
rect 7436 4864 7452 4928
rect 7516 4864 7524 4928
rect 7204 3840 7524 4864
rect 7204 3776 7212 3840
rect 7276 3776 7292 3840
rect 7356 3776 7372 3840
rect 7436 3776 7452 3840
rect 7516 3776 7524 3840
rect 7204 2752 7524 3776
rect 7204 2688 7212 2752
rect 7276 2688 7292 2752
rect 7356 2688 7372 2752
rect 7436 2688 7452 2752
rect 7516 2688 7524 2752
rect 7204 2672 7524 2688
rect 14433 13088 14753 14112
rect 14433 13024 14441 13088
rect 14505 13024 14521 13088
rect 14585 13024 14601 13088
rect 14665 13024 14681 13088
rect 14745 13024 14753 13088
rect 14433 12000 14753 13024
rect 14433 11936 14441 12000
rect 14505 11936 14521 12000
rect 14585 11936 14601 12000
rect 14665 11936 14681 12000
rect 14745 11936 14753 12000
rect 14433 10912 14753 11936
rect 14433 10848 14441 10912
rect 14505 10848 14521 10912
rect 14585 10848 14601 10912
rect 14665 10848 14681 10912
rect 14745 10848 14753 10912
rect 14433 9824 14753 10848
rect 14433 9760 14441 9824
rect 14505 9760 14521 9824
rect 14585 9760 14601 9824
rect 14665 9760 14681 9824
rect 14745 9760 14753 9824
rect 14433 8736 14753 9760
rect 14433 8672 14441 8736
rect 14505 8672 14521 8736
rect 14585 8672 14601 8736
rect 14665 8672 14681 8736
rect 14745 8672 14753 8736
rect 14433 7648 14753 8672
rect 14433 7584 14441 7648
rect 14505 7584 14521 7648
rect 14585 7584 14601 7648
rect 14665 7584 14681 7648
rect 14745 7584 14753 7648
rect 14433 6560 14753 7584
rect 14433 6496 14441 6560
rect 14505 6496 14521 6560
rect 14585 6496 14601 6560
rect 14665 6496 14681 6560
rect 14745 6496 14753 6560
rect 14433 5472 14753 6496
rect 14433 5408 14441 5472
rect 14505 5408 14521 5472
rect 14585 5408 14601 5472
rect 14665 5408 14681 5472
rect 14745 5408 14753 5472
rect 14433 4384 14753 5408
rect 14433 4320 14441 4384
rect 14505 4320 14521 4384
rect 14585 4320 14601 4384
rect 14665 4320 14681 4384
rect 14745 4320 14753 4384
rect 14433 3296 14753 4320
rect 14433 3232 14441 3296
rect 14505 3232 14521 3296
rect 14585 3232 14601 3296
rect 14665 3232 14681 3296
rect 14745 3232 14753 3296
rect 14433 2672 14753 3232
rect 15093 34304 15413 34320
rect 15093 34240 15101 34304
rect 15165 34240 15181 34304
rect 15245 34240 15261 34304
rect 15325 34240 15341 34304
rect 15405 34240 15413 34304
rect 15093 33216 15413 34240
rect 22322 33760 22642 34320
rect 22322 33696 22330 33760
rect 22394 33696 22410 33760
rect 22474 33696 22490 33760
rect 22554 33696 22570 33760
rect 22634 33696 22642 33760
rect 19195 33284 19261 33285
rect 19195 33220 19196 33284
rect 19260 33220 19261 33284
rect 19195 33219 19261 33220
rect 21587 33284 21653 33285
rect 21587 33220 21588 33284
rect 21652 33220 21653 33284
rect 21587 33219 21653 33220
rect 15093 33152 15101 33216
rect 15165 33152 15181 33216
rect 15245 33152 15261 33216
rect 15325 33152 15341 33216
rect 15405 33152 15413 33216
rect 15093 32128 15413 33152
rect 15093 32064 15101 32128
rect 15165 32064 15181 32128
rect 15245 32064 15261 32128
rect 15325 32064 15341 32128
rect 15405 32064 15413 32128
rect 15093 31040 15413 32064
rect 15093 30976 15101 31040
rect 15165 30976 15181 31040
rect 15245 30976 15261 31040
rect 15325 30976 15341 31040
rect 15405 30976 15413 31040
rect 15093 29952 15413 30976
rect 15093 29888 15101 29952
rect 15165 29888 15181 29952
rect 15245 29888 15261 29952
rect 15325 29888 15341 29952
rect 15405 29888 15413 29952
rect 15093 28864 15413 29888
rect 15093 28800 15101 28864
rect 15165 28800 15181 28864
rect 15245 28800 15261 28864
rect 15325 28800 15341 28864
rect 15405 28800 15413 28864
rect 15093 27776 15413 28800
rect 15093 27712 15101 27776
rect 15165 27712 15181 27776
rect 15245 27712 15261 27776
rect 15325 27712 15341 27776
rect 15405 27712 15413 27776
rect 15093 26688 15413 27712
rect 15093 26624 15101 26688
rect 15165 26624 15181 26688
rect 15245 26624 15261 26688
rect 15325 26624 15341 26688
rect 15405 26624 15413 26688
rect 15093 25600 15413 26624
rect 17355 26348 17421 26349
rect 17355 26284 17356 26348
rect 17420 26284 17421 26348
rect 17355 26283 17421 26284
rect 15093 25536 15101 25600
rect 15165 25536 15181 25600
rect 15245 25536 15261 25600
rect 15325 25536 15341 25600
rect 15405 25536 15413 25600
rect 15093 24512 15413 25536
rect 15093 24448 15101 24512
rect 15165 24448 15181 24512
rect 15245 24448 15261 24512
rect 15325 24448 15341 24512
rect 15405 24448 15413 24512
rect 15093 23424 15413 24448
rect 15699 23764 15765 23765
rect 15699 23700 15700 23764
rect 15764 23700 15765 23764
rect 15699 23699 15765 23700
rect 15093 23360 15101 23424
rect 15165 23360 15181 23424
rect 15245 23360 15261 23424
rect 15325 23360 15341 23424
rect 15405 23360 15413 23424
rect 15093 22336 15413 23360
rect 15093 22272 15101 22336
rect 15165 22272 15181 22336
rect 15245 22272 15261 22336
rect 15325 22272 15341 22336
rect 15405 22272 15413 22336
rect 15093 21248 15413 22272
rect 15093 21184 15101 21248
rect 15165 21184 15181 21248
rect 15245 21184 15261 21248
rect 15325 21184 15341 21248
rect 15405 21184 15413 21248
rect 15093 20160 15413 21184
rect 15093 20096 15101 20160
rect 15165 20096 15181 20160
rect 15245 20096 15261 20160
rect 15325 20096 15341 20160
rect 15405 20096 15413 20160
rect 15093 19072 15413 20096
rect 15093 19008 15101 19072
rect 15165 19008 15181 19072
rect 15245 19008 15261 19072
rect 15325 19008 15341 19072
rect 15405 19008 15413 19072
rect 15093 17984 15413 19008
rect 15093 17920 15101 17984
rect 15165 17920 15181 17984
rect 15245 17920 15261 17984
rect 15325 17920 15341 17984
rect 15405 17920 15413 17984
rect 15093 16896 15413 17920
rect 15093 16832 15101 16896
rect 15165 16832 15181 16896
rect 15245 16832 15261 16896
rect 15325 16832 15341 16896
rect 15405 16832 15413 16896
rect 15093 15808 15413 16832
rect 15093 15744 15101 15808
rect 15165 15744 15181 15808
rect 15245 15744 15261 15808
rect 15325 15744 15341 15808
rect 15405 15744 15413 15808
rect 15093 14720 15413 15744
rect 15093 14656 15101 14720
rect 15165 14656 15181 14720
rect 15245 14656 15261 14720
rect 15325 14656 15341 14720
rect 15405 14656 15413 14720
rect 15093 13632 15413 14656
rect 15093 13568 15101 13632
rect 15165 13568 15181 13632
rect 15245 13568 15261 13632
rect 15325 13568 15341 13632
rect 15405 13568 15413 13632
rect 15093 12544 15413 13568
rect 15093 12480 15101 12544
rect 15165 12480 15181 12544
rect 15245 12480 15261 12544
rect 15325 12480 15341 12544
rect 15405 12480 15413 12544
rect 15093 11456 15413 12480
rect 15093 11392 15101 11456
rect 15165 11392 15181 11456
rect 15245 11392 15261 11456
rect 15325 11392 15341 11456
rect 15405 11392 15413 11456
rect 15093 10368 15413 11392
rect 15093 10304 15101 10368
rect 15165 10304 15181 10368
rect 15245 10304 15261 10368
rect 15325 10304 15341 10368
rect 15405 10304 15413 10368
rect 15093 9280 15413 10304
rect 15093 9216 15101 9280
rect 15165 9216 15181 9280
rect 15245 9216 15261 9280
rect 15325 9216 15341 9280
rect 15405 9216 15413 9280
rect 15093 8192 15413 9216
rect 15093 8128 15101 8192
rect 15165 8128 15181 8192
rect 15245 8128 15261 8192
rect 15325 8128 15341 8192
rect 15405 8128 15413 8192
rect 15093 7104 15413 8128
rect 15093 7040 15101 7104
rect 15165 7040 15181 7104
rect 15245 7040 15261 7104
rect 15325 7040 15341 7104
rect 15405 7040 15413 7104
rect 15093 6016 15413 7040
rect 15093 5952 15101 6016
rect 15165 5952 15181 6016
rect 15245 5952 15261 6016
rect 15325 5952 15341 6016
rect 15405 5952 15413 6016
rect 15093 4928 15413 5952
rect 15093 4864 15101 4928
rect 15165 4864 15181 4928
rect 15245 4864 15261 4928
rect 15325 4864 15341 4928
rect 15405 4864 15413 4928
rect 15093 3840 15413 4864
rect 15093 3776 15101 3840
rect 15165 3776 15181 3840
rect 15245 3776 15261 3840
rect 15325 3776 15341 3840
rect 15405 3776 15413 3840
rect 15093 2752 15413 3776
rect 15702 3093 15762 23699
rect 17358 13837 17418 26283
rect 18827 15332 18893 15333
rect 18827 15268 18828 15332
rect 18892 15268 18893 15332
rect 18827 15267 18893 15268
rect 17355 13836 17421 13837
rect 17355 13772 17356 13836
rect 17420 13772 17421 13836
rect 17355 13771 17421 13772
rect 18830 8261 18890 15267
rect 19198 9621 19258 33219
rect 19379 20772 19445 20773
rect 19379 20708 19380 20772
rect 19444 20708 19445 20772
rect 19379 20707 19445 20708
rect 19195 9620 19261 9621
rect 19195 9556 19196 9620
rect 19260 9556 19261 9620
rect 19195 9555 19261 9556
rect 18827 8260 18893 8261
rect 18827 8196 18828 8260
rect 18892 8196 18893 8260
rect 18827 8195 18893 8196
rect 19382 8125 19442 20707
rect 19563 18052 19629 18053
rect 19563 17988 19564 18052
rect 19628 17988 19629 18052
rect 19563 17987 19629 17988
rect 19566 10981 19626 17987
rect 19747 17916 19813 17917
rect 19747 17852 19748 17916
rect 19812 17852 19813 17916
rect 19747 17851 19813 17852
rect 19750 15197 19810 17851
rect 19747 15196 19813 15197
rect 19747 15132 19748 15196
rect 19812 15132 19813 15196
rect 19747 15131 19813 15132
rect 19563 10980 19629 10981
rect 19563 10916 19564 10980
rect 19628 10916 19629 10980
rect 19563 10915 19629 10916
rect 21590 9485 21650 33219
rect 22322 32672 22642 33696
rect 22322 32608 22330 32672
rect 22394 32608 22410 32672
rect 22474 32608 22490 32672
rect 22554 32608 22570 32672
rect 22634 32608 22642 32672
rect 22322 31584 22642 32608
rect 22322 31520 22330 31584
rect 22394 31520 22410 31584
rect 22474 31520 22490 31584
rect 22554 31520 22570 31584
rect 22634 31520 22642 31584
rect 22322 30496 22642 31520
rect 22322 30432 22330 30496
rect 22394 30432 22410 30496
rect 22474 30432 22490 30496
rect 22554 30432 22570 30496
rect 22634 30432 22642 30496
rect 22322 29408 22642 30432
rect 22322 29344 22330 29408
rect 22394 29344 22410 29408
rect 22474 29344 22490 29408
rect 22554 29344 22570 29408
rect 22634 29344 22642 29408
rect 22322 28320 22642 29344
rect 22322 28256 22330 28320
rect 22394 28256 22410 28320
rect 22474 28256 22490 28320
rect 22554 28256 22570 28320
rect 22634 28256 22642 28320
rect 22322 27232 22642 28256
rect 22322 27168 22330 27232
rect 22394 27168 22410 27232
rect 22474 27168 22490 27232
rect 22554 27168 22570 27232
rect 22634 27168 22642 27232
rect 22322 26144 22642 27168
rect 22322 26080 22330 26144
rect 22394 26080 22410 26144
rect 22474 26080 22490 26144
rect 22554 26080 22570 26144
rect 22634 26080 22642 26144
rect 22322 25056 22642 26080
rect 22322 24992 22330 25056
rect 22394 24992 22410 25056
rect 22474 24992 22490 25056
rect 22554 24992 22570 25056
rect 22634 24992 22642 25056
rect 22322 23968 22642 24992
rect 22322 23904 22330 23968
rect 22394 23904 22410 23968
rect 22474 23904 22490 23968
rect 22554 23904 22570 23968
rect 22634 23904 22642 23968
rect 22322 22880 22642 23904
rect 22322 22816 22330 22880
rect 22394 22816 22410 22880
rect 22474 22816 22490 22880
rect 22554 22816 22570 22880
rect 22634 22816 22642 22880
rect 22322 21792 22642 22816
rect 22322 21728 22330 21792
rect 22394 21728 22410 21792
rect 22474 21728 22490 21792
rect 22554 21728 22570 21792
rect 22634 21728 22642 21792
rect 22322 20704 22642 21728
rect 22322 20640 22330 20704
rect 22394 20640 22410 20704
rect 22474 20640 22490 20704
rect 22554 20640 22570 20704
rect 22634 20640 22642 20704
rect 22322 19616 22642 20640
rect 22322 19552 22330 19616
rect 22394 19552 22410 19616
rect 22474 19552 22490 19616
rect 22554 19552 22570 19616
rect 22634 19552 22642 19616
rect 22322 18528 22642 19552
rect 22322 18464 22330 18528
rect 22394 18464 22410 18528
rect 22474 18464 22490 18528
rect 22554 18464 22570 18528
rect 22634 18464 22642 18528
rect 22139 17780 22205 17781
rect 22139 17716 22140 17780
rect 22204 17716 22205 17780
rect 22139 17715 22205 17716
rect 22142 11661 22202 17715
rect 22322 17440 22642 18464
rect 22322 17376 22330 17440
rect 22394 17376 22410 17440
rect 22474 17376 22490 17440
rect 22554 17376 22570 17440
rect 22634 17376 22642 17440
rect 22322 16352 22642 17376
rect 22322 16288 22330 16352
rect 22394 16288 22410 16352
rect 22474 16288 22490 16352
rect 22554 16288 22570 16352
rect 22634 16288 22642 16352
rect 22322 15264 22642 16288
rect 22322 15200 22330 15264
rect 22394 15200 22410 15264
rect 22474 15200 22490 15264
rect 22554 15200 22570 15264
rect 22634 15200 22642 15264
rect 22322 14176 22642 15200
rect 22322 14112 22330 14176
rect 22394 14112 22410 14176
rect 22474 14112 22490 14176
rect 22554 14112 22570 14176
rect 22634 14112 22642 14176
rect 22322 13088 22642 14112
rect 22322 13024 22330 13088
rect 22394 13024 22410 13088
rect 22474 13024 22490 13088
rect 22554 13024 22570 13088
rect 22634 13024 22642 13088
rect 22322 12000 22642 13024
rect 22322 11936 22330 12000
rect 22394 11936 22410 12000
rect 22474 11936 22490 12000
rect 22554 11936 22570 12000
rect 22634 11936 22642 12000
rect 22139 11660 22205 11661
rect 22139 11596 22140 11660
rect 22204 11596 22205 11660
rect 22139 11595 22205 11596
rect 22322 10912 22642 11936
rect 22322 10848 22330 10912
rect 22394 10848 22410 10912
rect 22474 10848 22490 10912
rect 22554 10848 22570 10912
rect 22634 10848 22642 10912
rect 22322 9824 22642 10848
rect 22322 9760 22330 9824
rect 22394 9760 22410 9824
rect 22474 9760 22490 9824
rect 22554 9760 22570 9824
rect 22634 9760 22642 9824
rect 21587 9484 21653 9485
rect 21587 9420 21588 9484
rect 21652 9420 21653 9484
rect 21587 9419 21653 9420
rect 22322 8736 22642 9760
rect 22322 8672 22330 8736
rect 22394 8672 22410 8736
rect 22474 8672 22490 8736
rect 22554 8672 22570 8736
rect 22634 8672 22642 8736
rect 19379 8124 19445 8125
rect 19379 8060 19380 8124
rect 19444 8060 19445 8124
rect 19379 8059 19445 8060
rect 22322 7648 22642 8672
rect 22322 7584 22330 7648
rect 22394 7584 22410 7648
rect 22474 7584 22490 7648
rect 22554 7584 22570 7648
rect 22634 7584 22642 7648
rect 22322 6560 22642 7584
rect 22322 6496 22330 6560
rect 22394 6496 22410 6560
rect 22474 6496 22490 6560
rect 22554 6496 22570 6560
rect 22634 6496 22642 6560
rect 22322 5472 22642 6496
rect 22322 5408 22330 5472
rect 22394 5408 22410 5472
rect 22474 5408 22490 5472
rect 22554 5408 22570 5472
rect 22634 5408 22642 5472
rect 22322 4384 22642 5408
rect 22322 4320 22330 4384
rect 22394 4320 22410 4384
rect 22474 4320 22490 4384
rect 22554 4320 22570 4384
rect 22634 4320 22642 4384
rect 22322 3296 22642 4320
rect 22322 3232 22330 3296
rect 22394 3232 22410 3296
rect 22474 3232 22490 3296
rect 22554 3232 22570 3296
rect 22634 3232 22642 3296
rect 15699 3092 15765 3093
rect 15699 3028 15700 3092
rect 15764 3028 15765 3092
rect 15699 3027 15765 3028
rect 15093 2688 15101 2752
rect 15165 2688 15181 2752
rect 15245 2688 15261 2752
rect 15325 2688 15341 2752
rect 15405 2688 15413 2752
rect 15093 2672 15413 2688
rect 22322 2672 22642 3232
rect 22982 34304 23302 34320
rect 22982 34240 22990 34304
rect 23054 34240 23070 34304
rect 23134 34240 23150 34304
rect 23214 34240 23230 34304
rect 23294 34240 23302 34304
rect 22982 33216 23302 34240
rect 22982 33152 22990 33216
rect 23054 33152 23070 33216
rect 23134 33152 23150 33216
rect 23214 33152 23230 33216
rect 23294 33152 23302 33216
rect 22982 32128 23302 33152
rect 22982 32064 22990 32128
rect 23054 32064 23070 32128
rect 23134 32064 23150 32128
rect 23214 32064 23230 32128
rect 23294 32064 23302 32128
rect 22982 31040 23302 32064
rect 22982 30976 22990 31040
rect 23054 30976 23070 31040
rect 23134 30976 23150 31040
rect 23214 30976 23230 31040
rect 23294 30976 23302 31040
rect 22982 29952 23302 30976
rect 22982 29888 22990 29952
rect 23054 29888 23070 29952
rect 23134 29888 23150 29952
rect 23214 29888 23230 29952
rect 23294 29888 23302 29952
rect 22982 28864 23302 29888
rect 30211 33760 30531 34320
rect 30211 33696 30219 33760
rect 30283 33696 30299 33760
rect 30363 33696 30379 33760
rect 30443 33696 30459 33760
rect 30523 33696 30531 33760
rect 30211 32672 30531 33696
rect 30211 32608 30219 32672
rect 30283 32608 30299 32672
rect 30363 32608 30379 32672
rect 30443 32608 30459 32672
rect 30523 32608 30531 32672
rect 30211 31584 30531 32608
rect 30211 31520 30219 31584
rect 30283 31520 30299 31584
rect 30363 31520 30379 31584
rect 30443 31520 30459 31584
rect 30523 31520 30531 31584
rect 30211 30496 30531 31520
rect 30211 30432 30219 30496
rect 30283 30432 30299 30496
rect 30363 30432 30379 30496
rect 30443 30432 30459 30496
rect 30523 30432 30531 30496
rect 30211 29408 30531 30432
rect 30211 29344 30219 29408
rect 30283 29344 30299 29408
rect 30363 29344 30379 29408
rect 30443 29344 30459 29408
rect 30523 29344 30531 29408
rect 27843 29068 27909 29069
rect 27843 29004 27844 29068
rect 27908 29004 27909 29068
rect 27843 29003 27909 29004
rect 22982 28800 22990 28864
rect 23054 28800 23070 28864
rect 23134 28800 23150 28864
rect 23214 28800 23230 28864
rect 23294 28800 23302 28864
rect 22982 27776 23302 28800
rect 22982 27712 22990 27776
rect 23054 27712 23070 27776
rect 23134 27712 23150 27776
rect 23214 27712 23230 27776
rect 23294 27712 23302 27776
rect 22982 26688 23302 27712
rect 22982 26624 22990 26688
rect 23054 26624 23070 26688
rect 23134 26624 23150 26688
rect 23214 26624 23230 26688
rect 23294 26624 23302 26688
rect 22982 25600 23302 26624
rect 22982 25536 22990 25600
rect 23054 25536 23070 25600
rect 23134 25536 23150 25600
rect 23214 25536 23230 25600
rect 23294 25536 23302 25600
rect 22982 24512 23302 25536
rect 22982 24448 22990 24512
rect 23054 24448 23070 24512
rect 23134 24448 23150 24512
rect 23214 24448 23230 24512
rect 23294 24448 23302 24512
rect 22982 23424 23302 24448
rect 26555 24036 26621 24037
rect 26555 23972 26556 24036
rect 26620 23972 26621 24036
rect 26555 23971 26621 23972
rect 22982 23360 22990 23424
rect 23054 23360 23070 23424
rect 23134 23360 23150 23424
rect 23214 23360 23230 23424
rect 23294 23360 23302 23424
rect 22982 22336 23302 23360
rect 22982 22272 22990 22336
rect 23054 22272 23070 22336
rect 23134 22272 23150 22336
rect 23214 22272 23230 22336
rect 23294 22272 23302 22336
rect 22982 21248 23302 22272
rect 22982 21184 22990 21248
rect 23054 21184 23070 21248
rect 23134 21184 23150 21248
rect 23214 21184 23230 21248
rect 23294 21184 23302 21248
rect 22982 20160 23302 21184
rect 22982 20096 22990 20160
rect 23054 20096 23070 20160
rect 23134 20096 23150 20160
rect 23214 20096 23230 20160
rect 23294 20096 23302 20160
rect 22982 19072 23302 20096
rect 22982 19008 22990 19072
rect 23054 19008 23070 19072
rect 23134 19008 23150 19072
rect 23214 19008 23230 19072
rect 23294 19008 23302 19072
rect 22982 17984 23302 19008
rect 22982 17920 22990 17984
rect 23054 17920 23070 17984
rect 23134 17920 23150 17984
rect 23214 17920 23230 17984
rect 23294 17920 23302 17984
rect 22982 16896 23302 17920
rect 22982 16832 22990 16896
rect 23054 16832 23070 16896
rect 23134 16832 23150 16896
rect 23214 16832 23230 16896
rect 23294 16832 23302 16896
rect 22982 15808 23302 16832
rect 22982 15744 22990 15808
rect 23054 15744 23070 15808
rect 23134 15744 23150 15808
rect 23214 15744 23230 15808
rect 23294 15744 23302 15808
rect 22982 14720 23302 15744
rect 22982 14656 22990 14720
rect 23054 14656 23070 14720
rect 23134 14656 23150 14720
rect 23214 14656 23230 14720
rect 23294 14656 23302 14720
rect 22982 13632 23302 14656
rect 22982 13568 22990 13632
rect 23054 13568 23070 13632
rect 23134 13568 23150 13632
rect 23214 13568 23230 13632
rect 23294 13568 23302 13632
rect 22982 12544 23302 13568
rect 22982 12480 22990 12544
rect 23054 12480 23070 12544
rect 23134 12480 23150 12544
rect 23214 12480 23230 12544
rect 23294 12480 23302 12544
rect 22982 11456 23302 12480
rect 22982 11392 22990 11456
rect 23054 11392 23070 11456
rect 23134 11392 23150 11456
rect 23214 11392 23230 11456
rect 23294 11392 23302 11456
rect 22982 10368 23302 11392
rect 22982 10304 22990 10368
rect 23054 10304 23070 10368
rect 23134 10304 23150 10368
rect 23214 10304 23230 10368
rect 23294 10304 23302 10368
rect 22982 9280 23302 10304
rect 22982 9216 22990 9280
rect 23054 9216 23070 9280
rect 23134 9216 23150 9280
rect 23214 9216 23230 9280
rect 23294 9216 23302 9280
rect 22982 8192 23302 9216
rect 22982 8128 22990 8192
rect 23054 8128 23070 8192
rect 23134 8128 23150 8192
rect 23214 8128 23230 8192
rect 23294 8128 23302 8192
rect 22982 7104 23302 8128
rect 26558 7989 26618 23971
rect 27846 12885 27906 29003
rect 30211 28320 30531 29344
rect 30211 28256 30219 28320
rect 30283 28256 30299 28320
rect 30363 28256 30379 28320
rect 30443 28256 30459 28320
rect 30523 28256 30531 28320
rect 30211 27232 30531 28256
rect 30211 27168 30219 27232
rect 30283 27168 30299 27232
rect 30363 27168 30379 27232
rect 30443 27168 30459 27232
rect 30523 27168 30531 27232
rect 30211 26144 30531 27168
rect 30211 26080 30219 26144
rect 30283 26080 30299 26144
rect 30363 26080 30379 26144
rect 30443 26080 30459 26144
rect 30523 26080 30531 26144
rect 30211 25056 30531 26080
rect 30211 24992 30219 25056
rect 30283 24992 30299 25056
rect 30363 24992 30379 25056
rect 30443 24992 30459 25056
rect 30523 24992 30531 25056
rect 30211 23968 30531 24992
rect 30211 23904 30219 23968
rect 30283 23904 30299 23968
rect 30363 23904 30379 23968
rect 30443 23904 30459 23968
rect 30523 23904 30531 23968
rect 30211 22880 30531 23904
rect 30211 22816 30219 22880
rect 30283 22816 30299 22880
rect 30363 22816 30379 22880
rect 30443 22816 30459 22880
rect 30523 22816 30531 22880
rect 30211 21792 30531 22816
rect 30211 21728 30219 21792
rect 30283 21728 30299 21792
rect 30363 21728 30379 21792
rect 30443 21728 30459 21792
rect 30523 21728 30531 21792
rect 30211 20704 30531 21728
rect 30211 20640 30219 20704
rect 30283 20640 30299 20704
rect 30363 20640 30379 20704
rect 30443 20640 30459 20704
rect 30523 20640 30531 20704
rect 30211 19616 30531 20640
rect 30211 19552 30219 19616
rect 30283 19552 30299 19616
rect 30363 19552 30379 19616
rect 30443 19552 30459 19616
rect 30523 19552 30531 19616
rect 30211 18528 30531 19552
rect 30211 18464 30219 18528
rect 30283 18464 30299 18528
rect 30363 18464 30379 18528
rect 30443 18464 30459 18528
rect 30523 18464 30531 18528
rect 30211 17440 30531 18464
rect 30211 17376 30219 17440
rect 30283 17376 30299 17440
rect 30363 17376 30379 17440
rect 30443 17376 30459 17440
rect 30523 17376 30531 17440
rect 30211 16352 30531 17376
rect 30211 16288 30219 16352
rect 30283 16288 30299 16352
rect 30363 16288 30379 16352
rect 30443 16288 30459 16352
rect 30523 16288 30531 16352
rect 30211 15264 30531 16288
rect 30211 15200 30219 15264
rect 30283 15200 30299 15264
rect 30363 15200 30379 15264
rect 30443 15200 30459 15264
rect 30523 15200 30531 15264
rect 30211 14176 30531 15200
rect 30211 14112 30219 14176
rect 30283 14112 30299 14176
rect 30363 14112 30379 14176
rect 30443 14112 30459 14176
rect 30523 14112 30531 14176
rect 30211 13088 30531 14112
rect 30211 13024 30219 13088
rect 30283 13024 30299 13088
rect 30363 13024 30379 13088
rect 30443 13024 30459 13088
rect 30523 13024 30531 13088
rect 27843 12884 27909 12885
rect 27843 12820 27844 12884
rect 27908 12820 27909 12884
rect 27843 12819 27909 12820
rect 30211 12000 30531 13024
rect 30211 11936 30219 12000
rect 30283 11936 30299 12000
rect 30363 11936 30379 12000
rect 30443 11936 30459 12000
rect 30523 11936 30531 12000
rect 30211 10912 30531 11936
rect 30211 10848 30219 10912
rect 30283 10848 30299 10912
rect 30363 10848 30379 10912
rect 30443 10848 30459 10912
rect 30523 10848 30531 10912
rect 30211 9824 30531 10848
rect 30211 9760 30219 9824
rect 30283 9760 30299 9824
rect 30363 9760 30379 9824
rect 30443 9760 30459 9824
rect 30523 9760 30531 9824
rect 30211 8736 30531 9760
rect 30211 8672 30219 8736
rect 30283 8672 30299 8736
rect 30363 8672 30379 8736
rect 30443 8672 30459 8736
rect 30523 8672 30531 8736
rect 26555 7988 26621 7989
rect 26555 7924 26556 7988
rect 26620 7924 26621 7988
rect 26555 7923 26621 7924
rect 22982 7040 22990 7104
rect 23054 7040 23070 7104
rect 23134 7040 23150 7104
rect 23214 7040 23230 7104
rect 23294 7040 23302 7104
rect 22982 6016 23302 7040
rect 22982 5952 22990 6016
rect 23054 5952 23070 6016
rect 23134 5952 23150 6016
rect 23214 5952 23230 6016
rect 23294 5952 23302 6016
rect 22982 4928 23302 5952
rect 22982 4864 22990 4928
rect 23054 4864 23070 4928
rect 23134 4864 23150 4928
rect 23214 4864 23230 4928
rect 23294 4864 23302 4928
rect 22982 3840 23302 4864
rect 22982 3776 22990 3840
rect 23054 3776 23070 3840
rect 23134 3776 23150 3840
rect 23214 3776 23230 3840
rect 23294 3776 23302 3840
rect 22982 2752 23302 3776
rect 22982 2688 22990 2752
rect 23054 2688 23070 2752
rect 23134 2688 23150 2752
rect 23214 2688 23230 2752
rect 23294 2688 23302 2752
rect 22982 2672 23302 2688
rect 30211 7648 30531 8672
rect 30211 7584 30219 7648
rect 30283 7584 30299 7648
rect 30363 7584 30379 7648
rect 30443 7584 30459 7648
rect 30523 7584 30531 7648
rect 30211 6560 30531 7584
rect 30211 6496 30219 6560
rect 30283 6496 30299 6560
rect 30363 6496 30379 6560
rect 30443 6496 30459 6560
rect 30523 6496 30531 6560
rect 30211 5472 30531 6496
rect 30211 5408 30219 5472
rect 30283 5408 30299 5472
rect 30363 5408 30379 5472
rect 30443 5408 30459 5472
rect 30523 5408 30531 5472
rect 30211 4384 30531 5408
rect 30211 4320 30219 4384
rect 30283 4320 30299 4384
rect 30363 4320 30379 4384
rect 30443 4320 30459 4384
rect 30523 4320 30531 4384
rect 30211 3296 30531 4320
rect 30211 3232 30219 3296
rect 30283 3232 30299 3296
rect 30363 3232 30379 3296
rect 30443 3232 30459 3296
rect 30523 3232 30531 3296
rect 30211 2672 30531 3232
rect 30871 34304 31191 34320
rect 30871 34240 30879 34304
rect 30943 34240 30959 34304
rect 31023 34240 31039 34304
rect 31103 34240 31119 34304
rect 31183 34240 31191 34304
rect 30871 33216 31191 34240
rect 30871 33152 30879 33216
rect 30943 33152 30959 33216
rect 31023 33152 31039 33216
rect 31103 33152 31119 33216
rect 31183 33152 31191 33216
rect 30871 32128 31191 33152
rect 30871 32064 30879 32128
rect 30943 32064 30959 32128
rect 31023 32064 31039 32128
rect 31103 32064 31119 32128
rect 31183 32064 31191 32128
rect 30871 31040 31191 32064
rect 30871 30976 30879 31040
rect 30943 30976 30959 31040
rect 31023 30976 31039 31040
rect 31103 30976 31119 31040
rect 31183 30976 31191 31040
rect 30871 29952 31191 30976
rect 30871 29888 30879 29952
rect 30943 29888 30959 29952
rect 31023 29888 31039 29952
rect 31103 29888 31119 29952
rect 31183 29888 31191 29952
rect 30871 28864 31191 29888
rect 30871 28800 30879 28864
rect 30943 28800 30959 28864
rect 31023 28800 31039 28864
rect 31103 28800 31119 28864
rect 31183 28800 31191 28864
rect 30871 27776 31191 28800
rect 30871 27712 30879 27776
rect 30943 27712 30959 27776
rect 31023 27712 31039 27776
rect 31103 27712 31119 27776
rect 31183 27712 31191 27776
rect 30871 26688 31191 27712
rect 30871 26624 30879 26688
rect 30943 26624 30959 26688
rect 31023 26624 31039 26688
rect 31103 26624 31119 26688
rect 31183 26624 31191 26688
rect 30871 25600 31191 26624
rect 30871 25536 30879 25600
rect 30943 25536 30959 25600
rect 31023 25536 31039 25600
rect 31103 25536 31119 25600
rect 31183 25536 31191 25600
rect 30871 24512 31191 25536
rect 30871 24448 30879 24512
rect 30943 24448 30959 24512
rect 31023 24448 31039 24512
rect 31103 24448 31119 24512
rect 31183 24448 31191 24512
rect 30871 23424 31191 24448
rect 30871 23360 30879 23424
rect 30943 23360 30959 23424
rect 31023 23360 31039 23424
rect 31103 23360 31119 23424
rect 31183 23360 31191 23424
rect 30871 22336 31191 23360
rect 30871 22272 30879 22336
rect 30943 22272 30959 22336
rect 31023 22272 31039 22336
rect 31103 22272 31119 22336
rect 31183 22272 31191 22336
rect 30871 21248 31191 22272
rect 30871 21184 30879 21248
rect 30943 21184 30959 21248
rect 31023 21184 31039 21248
rect 31103 21184 31119 21248
rect 31183 21184 31191 21248
rect 30871 20160 31191 21184
rect 30871 20096 30879 20160
rect 30943 20096 30959 20160
rect 31023 20096 31039 20160
rect 31103 20096 31119 20160
rect 31183 20096 31191 20160
rect 30871 19072 31191 20096
rect 30871 19008 30879 19072
rect 30943 19008 30959 19072
rect 31023 19008 31039 19072
rect 31103 19008 31119 19072
rect 31183 19008 31191 19072
rect 30871 17984 31191 19008
rect 30871 17920 30879 17984
rect 30943 17920 30959 17984
rect 31023 17920 31039 17984
rect 31103 17920 31119 17984
rect 31183 17920 31191 17984
rect 30871 16896 31191 17920
rect 30871 16832 30879 16896
rect 30943 16832 30959 16896
rect 31023 16832 31039 16896
rect 31103 16832 31119 16896
rect 31183 16832 31191 16896
rect 30871 15808 31191 16832
rect 30871 15744 30879 15808
rect 30943 15744 30959 15808
rect 31023 15744 31039 15808
rect 31103 15744 31119 15808
rect 31183 15744 31191 15808
rect 30871 14720 31191 15744
rect 30871 14656 30879 14720
rect 30943 14656 30959 14720
rect 31023 14656 31039 14720
rect 31103 14656 31119 14720
rect 31183 14656 31191 14720
rect 30871 13632 31191 14656
rect 30871 13568 30879 13632
rect 30943 13568 30959 13632
rect 31023 13568 31039 13632
rect 31103 13568 31119 13632
rect 31183 13568 31191 13632
rect 30871 12544 31191 13568
rect 30871 12480 30879 12544
rect 30943 12480 30959 12544
rect 31023 12480 31039 12544
rect 31103 12480 31119 12544
rect 31183 12480 31191 12544
rect 30871 11456 31191 12480
rect 30871 11392 30879 11456
rect 30943 11392 30959 11456
rect 31023 11392 31039 11456
rect 31103 11392 31119 11456
rect 31183 11392 31191 11456
rect 30871 10368 31191 11392
rect 30871 10304 30879 10368
rect 30943 10304 30959 10368
rect 31023 10304 31039 10368
rect 31103 10304 31119 10368
rect 31183 10304 31191 10368
rect 30871 9280 31191 10304
rect 30871 9216 30879 9280
rect 30943 9216 30959 9280
rect 31023 9216 31039 9280
rect 31103 9216 31119 9280
rect 31183 9216 31191 9280
rect 30871 8192 31191 9216
rect 30871 8128 30879 8192
rect 30943 8128 30959 8192
rect 31023 8128 31039 8192
rect 31103 8128 31119 8192
rect 31183 8128 31191 8192
rect 30871 7104 31191 8128
rect 30871 7040 30879 7104
rect 30943 7040 30959 7104
rect 31023 7040 31039 7104
rect 31103 7040 31119 7104
rect 31183 7040 31191 7104
rect 30871 6016 31191 7040
rect 30871 5952 30879 6016
rect 30943 5952 30959 6016
rect 31023 5952 31039 6016
rect 31103 5952 31119 6016
rect 31183 5952 31191 6016
rect 30871 4928 31191 5952
rect 30871 4864 30879 4928
rect 30943 4864 30959 4928
rect 31023 4864 31039 4928
rect 31103 4864 31119 4928
rect 31183 4864 31191 4928
rect 30871 3840 31191 4864
rect 30871 3776 30879 3840
rect 30943 3776 30959 3840
rect 31023 3776 31039 3840
rect 31103 3776 31119 3840
rect 31183 3776 31191 3840
rect 30871 2752 31191 3776
rect 30871 2688 30879 2752
rect 30943 2688 30959 2752
rect 31023 2688 31039 2752
rect 31103 2688 31119 2752
rect 31183 2688 31191 2752
rect 30871 2672 31191 2688
use sky130_fd_sc_hd__inv_2  _0709_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25392 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1688980957
transform 1 0 18952 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0711_
timestamp 1688980957
transform 1 0 10580 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1688980957
transform 1 0 13156 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1688980957
transform -1 0 11868 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1688980957
transform -1 0 12052 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1688980957
transform -1 0 15364 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0716_
timestamp 1688980957
transform 1 0 14260 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1688980957
transform -1 0 10212 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1688980957
transform 1 0 27048 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1688980957
transform -1 0 16560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1688980957
transform -1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1688980957
transform -1 0 15548 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0722_
timestamp 1688980957
transform 1 0 15088 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0723_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0724_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0725_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0726_
timestamp 1688980957
transform -1 0 11132 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0727_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10212 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1688980957
transform 1 0 10212 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0729_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0730_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0731_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12328 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0732_
timestamp 1688980957
transform -1 0 14352 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0733_
timestamp 1688980957
transform -1 0 13064 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0734_
timestamp 1688980957
transform -1 0 11868 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0735_
timestamp 1688980957
transform 1 0 10028 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0736_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11960 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0737_
timestamp 1688980957
transform -1 0 14168 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_1  _0738_
timestamp 1688980957
transform 1 0 11316 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _0739_
timestamp 1688980957
transform -1 0 13892 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0740_
timestamp 1688980957
transform -1 0 13616 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0741_
timestamp 1688980957
transform -1 0 11960 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0742_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9936 0 1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0743_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9752 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0744_
timestamp 1688980957
transform -1 0 11684 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0745_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10488 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0746_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0747_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0748_
timestamp 1688980957
transform -1 0 10120 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0749_
timestamp 1688980957
transform -1 0 10396 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0750_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9016 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and4bb_1  _0751_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9752 0 -1 20128
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _0752_
timestamp 1688980957
transform -1 0 9016 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0753_
timestamp 1688980957
transform -1 0 11592 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0754_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12052 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0755_
timestamp 1688980957
transform -1 0 11132 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0756_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9936 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0757_
timestamp 1688980957
transform 1 0 11868 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0758_
timestamp 1688980957
transform 1 0 10856 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0759_
timestamp 1688980957
transform -1 0 11868 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0760_
timestamp 1688980957
transform 1 0 11868 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0761_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12604 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _0762_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _0763_
timestamp 1688980957
transform -1 0 11684 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0764_
timestamp 1688980957
transform 1 0 12052 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0765_
timestamp 1688980957
transform 1 0 11868 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0766_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29072 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0767_
timestamp 1688980957
transform -1 0 28428 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0768_
timestamp 1688980957
transform 1 0 30360 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0769_
timestamp 1688980957
transform -1 0 30084 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0770_
timestamp 1688980957
transform 1 0 26864 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0771_
timestamp 1688980957
transform 1 0 28612 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0772_
timestamp 1688980957
transform -1 0 29624 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0773_
timestamp 1688980957
transform 1 0 27968 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0774_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0775_
timestamp 1688980957
transform -1 0 23368 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _0776_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27324 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0777_
timestamp 1688980957
transform -1 0 29716 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or4bb_1  _0778_
timestamp 1688980957
transform -1 0 28428 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _0779_
timestamp 1688980957
transform -1 0 28520 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0780_
timestamp 1688980957
transform -1 0 27784 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0781_
timestamp 1688980957
transform 1 0 27416 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0782_
timestamp 1688980957
transform -1 0 27416 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0783_
timestamp 1688980957
transform -1 0 28244 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0784_
timestamp 1688980957
transform -1 0 31648 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0785_
timestamp 1688980957
transform -1 0 29624 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0786_
timestamp 1688980957
transform -1 0 28888 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0787_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30360 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0788_
timestamp 1688980957
transform 1 0 29532 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0789_
timestamp 1688980957
transform -1 0 29072 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0790_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27416 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0791_
timestamp 1688980957
transform 1 0 26864 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1688980957
transform 1 0 26956 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0793_
timestamp 1688980957
transform -1 0 27600 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0794_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26864 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _0795_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27876 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1688980957
transform -1 0 28612 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0797_
timestamp 1688980957
transform -1 0 29900 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0798_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29716 0 1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0799_
timestamp 1688980957
transform 1 0 29532 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0800_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27324 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_2  _0801_
timestamp 1688980957
transform 1 0 26036 0 1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0802_
timestamp 1688980957
transform 1 0 23092 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0803_
timestamp 1688980957
transform 1 0 28888 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0804_
timestamp 1688980957
transform -1 0 29716 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0805_
timestamp 1688980957
transform 1 0 26220 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0806_
timestamp 1688980957
transform -1 0 28152 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0807_
timestamp 1688980957
transform -1 0 25944 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0808_
timestamp 1688980957
transform -1 0 24380 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0809_
timestamp 1688980957
transform 1 0 26036 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0810_
timestamp 1688980957
transform -1 0 25852 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _0811_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28612 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0812_
timestamp 1688980957
transform -1 0 27048 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0813_
timestamp 1688980957
transform 1 0 29716 0 1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0814_
timestamp 1688980957
transform 1 0 26772 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0815_
timestamp 1688980957
transform 1 0 30084 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0816_
timestamp 1688980957
transform -1 0 30636 0 -1 16864
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0817_
timestamp 1688980957
transform 1 0 29532 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0818_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29348 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0819_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29716 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0820_
timestamp 1688980957
transform -1 0 29624 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0821_
timestamp 1688980957
transform 1 0 27968 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1688980957
transform -1 0 32016 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0823_
timestamp 1688980957
transform 1 0 30636 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _0824_
timestamp 1688980957
transform -1 0 30820 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0825_
timestamp 1688980957
transform 1 0 30452 0 1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0826_
timestamp 1688980957
transform 1 0 30084 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0827_
timestamp 1688980957
transform 1 0 30636 0 -1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0828_
timestamp 1688980957
transform 1 0 30544 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0829_
timestamp 1688980957
transform -1 0 32016 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1688980957
transform -1 0 31096 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0831_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29256 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1688980957
transform 1 0 31648 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0833_
timestamp 1688980957
transform -1 0 30360 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0834_
timestamp 1688980957
transform 1 0 29440 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0835_
timestamp 1688980957
transform 1 0 31188 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1688980957
transform -1 0 32660 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0837_
timestamp 1688980957
transform -1 0 30360 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0838_
timestamp 1688980957
transform 1 0 29348 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0839_
timestamp 1688980957
transform 1 0 27784 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0840_
timestamp 1688980957
transform -1 0 28336 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0841_
timestamp 1688980957
transform 1 0 26864 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0842_
timestamp 1688980957
transform 1 0 26128 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0843_
timestamp 1688980957
transform -1 0 27324 0 -1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0844_
timestamp 1688980957
transform 1 0 26128 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0845_
timestamp 1688980957
transform -1 0 27048 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0846_
timestamp 1688980957
transform -1 0 26128 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0847_
timestamp 1688980957
transform 1 0 25668 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0848_
timestamp 1688980957
transform 1 0 25852 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0849_
timestamp 1688980957
transform 1 0 25392 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0850_
timestamp 1688980957
transform -1 0 26956 0 -1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1688980957
transform 1 0 28336 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0852_
timestamp 1688980957
transform -1 0 28152 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _0853_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 -1 12512
box -38 -48 1970 592
use sky130_fd_sc_hd__a22o_1  _0854_
timestamp 1688980957
transform -1 0 26680 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0855_
timestamp 1688980957
transform -1 0 26036 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0856_
timestamp 1688980957
transform -1 0 26680 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0857_
timestamp 1688980957
transform 1 0 28612 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1688980957
transform -1 0 29624 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1688980957
transform -1 0 24380 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1688980957
transform -1 0 25300 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1688980957
transform 1 0 21988 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 1688980957
transform -1 0 26956 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp 1688980957
transform -1 0 24196 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1688980957
transform -1 0 25116 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0865_
timestamp 1688980957
transform -1 0 23368 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0866_
timestamp 1688980957
transform 1 0 10304 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0867_
timestamp 1688980957
transform 1 0 8004 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0868_
timestamp 1688980957
transform -1 0 9568 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0869_
timestamp 1688980957
transform -1 0 9108 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0870_
timestamp 1688980957
transform -1 0 13248 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0871_
timestamp 1688980957
transform -1 0 15180 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0872_
timestamp 1688980957
transform -1 0 14904 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0873_
timestamp 1688980957
transform 1 0 13340 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0874_
timestamp 1688980957
transform 1 0 14536 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1688980957
transform 1 0 11868 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1688980957
transform -1 0 12604 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0877_
timestamp 1688980957
transform 1 0 10764 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0878_
timestamp 1688980957
transform 1 0 8280 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0879_
timestamp 1688980957
transform 1 0 8004 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0880_
timestamp 1688980957
transform 1 0 8004 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0881_
timestamp 1688980957
transform 1 0 8832 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0882_
timestamp 1688980957
transform -1 0 10120 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _0883_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0884_
timestamp 1688980957
transform 1 0 9200 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _0885_
timestamp 1688980957
transform -1 0 11040 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__and4_2  _0886_
timestamp 1688980957
transform 1 0 10580 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0887_
timestamp 1688980957
transform 1 0 13616 0 1 26656
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1688980957
transform 1 0 14076 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0889_
timestamp 1688980957
transform -1 0 16744 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0890_
timestamp 1688980957
transform 1 0 13892 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0891_
timestamp 1688980957
transform 1 0 14536 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _0892_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14352 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0893_
timestamp 1688980957
transform -1 0 12328 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0894_
timestamp 1688980957
transform 1 0 12328 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0895_
timestamp 1688980957
transform -1 0 11684 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0896_
timestamp 1688980957
transform 1 0 11868 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0897_
timestamp 1688980957
transform -1 0 12328 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0898_
timestamp 1688980957
transform 1 0 12236 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0899_
timestamp 1688980957
transform -1 0 11040 0 1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0900_
timestamp 1688980957
transform 1 0 11316 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0901_
timestamp 1688980957
transform 1 0 10580 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0902_
timestamp 1688980957
transform -1 0 11500 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0903_
timestamp 1688980957
transform 1 0 13156 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0904_
timestamp 1688980957
transform 1 0 11592 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0905_
timestamp 1688980957
transform -1 0 11040 0 1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0906_
timestamp 1688980957
transform -1 0 12328 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0907_
timestamp 1688980957
transform 1 0 9752 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0908_
timestamp 1688980957
transform 1 0 15548 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0909_
timestamp 1688980957
transform 1 0 13800 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1688980957
transform -1 0 14996 0 -1 32096
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _0911_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0912_
timestamp 1688980957
transform 1 0 14720 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0913_
timestamp 1688980957
transform -1 0 15640 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0914_
timestamp 1688980957
transform -1 0 16560 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _0915_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14444 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1688980957
transform 1 0 15732 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0917_
timestamp 1688980957
transform 1 0 12788 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0918_
timestamp 1688980957
transform 1 0 13984 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0919_
timestamp 1688980957
transform 1 0 13432 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0920_
timestamp 1688980957
transform -1 0 15088 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1688980957
transform 1 0 16100 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0922_
timestamp 1688980957
transform -1 0 11960 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0923_
timestamp 1688980957
transform 1 0 11960 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0924_
timestamp 1688980957
transform 1 0 15272 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0925_
timestamp 1688980957
transform -1 0 14812 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0926_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14168 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0927_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15272 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0928_
timestamp 1688980957
transform 1 0 10580 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0929_
timestamp 1688980957
transform 1 0 9568 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0930_
timestamp 1688980957
transform 1 0 10212 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0931_
timestamp 1688980957
transform 1 0 9936 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0932_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11868 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0933_
timestamp 1688980957
transform 1 0 10672 0 -1 27744
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_1  _0934_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0935_
timestamp 1688980957
transform 1 0 9384 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1688980957
transform -1 0 8372 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_2  _0937_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0938_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21344 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0939_
timestamp 1688980957
transform 1 0 19044 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0940_
timestamp 1688980957
transform 1 0 19412 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0941_
timestamp 1688980957
transform 1 0 18308 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0942_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17572 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0943_
timestamp 1688980957
transform 1 0 16468 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1688980957
transform -1 0 16836 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0945_
timestamp 1688980957
transform 1 0 16928 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0946_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_2  _0947_
timestamp 1688980957
transform -1 0 18308 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0948_
timestamp 1688980957
transform 1 0 14444 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0949_
timestamp 1688980957
transform -1 0 18032 0 -1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__nor3b_1  _0950_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _0951_
timestamp 1688980957
transform -1 0 16376 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _0952_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1688980957
transform 1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0954_
timestamp 1688980957
transform 1 0 17112 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0955_
timestamp 1688980957
transform 1 0 16744 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0956_
timestamp 1688980957
transform 1 0 17480 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__and4bb_2  _0957_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16100 0 -1 11424
box -38 -48 958 592
use sky130_fd_sc_hd__or3b_1  _0958_
timestamp 1688980957
transform -1 0 17664 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0959_
timestamp 1688980957
transform 1 0 17020 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0960_
timestamp 1688980957
transform 1 0 16652 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0961_
timestamp 1688980957
transform -1 0 18216 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0962_
timestamp 1688980957
transform 1 0 14904 0 1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0963_
timestamp 1688980957
transform 1 0 15180 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0964_
timestamp 1688980957
transform 1 0 15732 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0965_
timestamp 1688980957
transform 1 0 15732 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0966_
timestamp 1688980957
transform 1 0 14812 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _0967_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18584 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0968_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20884 0 -1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0969_
timestamp 1688980957
transform 1 0 18952 0 -1 20128
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0970_
timestamp 1688980957
transform 1 0 16928 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_4  _0971_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_1  _0972_
timestamp 1688980957
transform 1 0 21344 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _0973_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19688 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0974_
timestamp 1688980957
transform 1 0 22632 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _0975_
timestamp 1688980957
transform -1 0 9936 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0976_
timestamp 1688980957
transform 1 0 7912 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _0977_
timestamp 1688980957
transform 1 0 10580 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0978_
timestamp 1688980957
transform -1 0 10488 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _0979_
timestamp 1688980957
transform 1 0 5704 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0980_
timestamp 1688980957
transform 1 0 5428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0981_
timestamp 1688980957
transform 1 0 18308 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0982_
timestamp 1688980957
transform 1 0 16652 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0983_
timestamp 1688980957
transform 1 0 4692 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0984_
timestamp 1688980957
transform 1 0 5428 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0985_
timestamp 1688980957
transform 1 0 19136 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0986_
timestamp 1688980957
transform 1 0 19596 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1688980957
transform 1 0 19136 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0988_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19688 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0989_
timestamp 1688980957
transform 1 0 6256 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0990_
timestamp 1688980957
transform -1 0 7636 0 1 12512
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0991_
timestamp 1688980957
transform -1 0 4416 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0992_
timestamp 1688980957
transform 1 0 7084 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0993_
timestamp 1688980957
transform -1 0 8464 0 -1 15776
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0994_
timestamp 1688980957
transform 1 0 5612 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0995_
timestamp 1688980957
transform 1 0 17572 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0996_
timestamp 1688980957
transform 1 0 18676 0 1 24480
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0997_
timestamp 1688980957
transform -1 0 19688 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0998_
timestamp 1688980957
transform 1 0 10764 0 -1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0999_
timestamp 1688980957
transform -1 0 12696 0 -1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1000_
timestamp 1688980957
transform 1 0 11592 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1001_
timestamp 1688980957
transform 1 0 18032 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1002_
timestamp 1688980957
transform -1 0 19044 0 -1 25568
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1003_
timestamp 1688980957
transform 1 0 22724 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1004_
timestamp 1688980957
transform 1 0 17572 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1688980957
transform 1 0 19044 0 -1 22304
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1006_
timestamp 1688980957
transform 1 0 26404 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1007_
timestamp 1688980957
transform -1 0 7268 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1008_
timestamp 1688980957
transform -1 0 8464 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1009_
timestamp 1688980957
transform 1 0 6256 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1010_
timestamp 1688980957
transform 1 0 19044 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1011_
timestamp 1688980957
transform 1 0 19688 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1012_
timestamp 1688980957
transform -1 0 24104 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1688980957
transform -1 0 21252 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1014_
timestamp 1688980957
transform -1 0 21528 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1015_
timestamp 1688980957
transform 1 0 23828 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1016_
timestamp 1688980957
transform 1 0 24380 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1017_
timestamp 1688980957
transform -1 0 27140 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1688980957
transform -1 0 28060 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1019_
timestamp 1688980957
transform -1 0 27324 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1020_
timestamp 1688980957
transform -1 0 27968 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1021_
timestamp 1688980957
transform -1 0 6164 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1022_
timestamp 1688980957
transform -1 0 12052 0 -1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1023_
timestamp 1688980957
transform 1 0 19136 0 1 21216
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1024_
timestamp 1688980957
transform 1 0 12512 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1025_
timestamp 1688980957
transform -1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1026_
timestamp 1688980957
transform -1 0 7360 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1027_
timestamp 1688980957
transform -1 0 19136 0 -1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1028_
timestamp 1688980957
transform 1 0 20148 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _1029_
timestamp 1688980957
transform -1 0 13432 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_4  _1030_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18952 0 1 10336
box -38 -48 958 592
use sky130_fd_sc_hd__nand3b_4  _1031_
timestamp 1688980957
transform 1 0 20884 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _1032_
timestamp 1688980957
transform -1 0 8740 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1033_
timestamp 1688980957
transform -1 0 7544 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1034_
timestamp 1688980957
transform 1 0 18676 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1035_
timestamp 1688980957
transform 1 0 10764 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1036_
timestamp 1688980957
transform 1 0 19044 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1037_
timestamp 1688980957
transform -1 0 18952 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1038_
timestamp 1688980957
transform -1 0 6716 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1039_
timestamp 1688980957
transform 1 0 19596 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1040_
timestamp 1688980957
transform 1 0 21344 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1041_
timestamp 1688980957
transform 1 0 27784 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1042_
timestamp 1688980957
transform -1 0 29072 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1043_
timestamp 1688980957
transform 1 0 27784 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1044_
timestamp 1688980957
transform 1 0 5888 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1045_
timestamp 1688980957
transform 1 0 19412 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1046_
timestamp 1688980957
transform 1 0 5428 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _1047_
timestamp 1688980957
transform 1 0 20884 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1048_
timestamp 1688980957
transform -1 0 6256 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1049_
timestamp 1688980957
transform -1 0 6900 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1050_
timestamp 1688980957
transform -1 0 26680 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1051_
timestamp 1688980957
transform 1 0 9200 0 1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1052_
timestamp 1688980957
transform -1 0 18216 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1053_
timestamp 1688980957
transform -1 0 22908 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1054_
timestamp 1688980957
transform -1 0 9200 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1055_
timestamp 1688980957
transform 1 0 29164 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1056_
timestamp 1688980957
transform -1 0 22264 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1057_
timestamp 1688980957
transform 1 0 28980 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1058_
timestamp 1688980957
transform -1 0 29256 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1059_
timestamp 1688980957
transform 1 0 28888 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1060_
timestamp 1688980957
transform 1 0 6164 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1061_
timestamp 1688980957
transform -1 0 26680 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1062_
timestamp 1688980957
transform -1 0 5980 0 -1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1063_
timestamp 1688980957
transform -1 0 6072 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1064_
timestamp 1688980957
transform 1 0 11040 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1065_
timestamp 1688980957
transform 1 0 10856 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1066_
timestamp 1688980957
transform 1 0 13156 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1067_
timestamp 1688980957
transform 1 0 13156 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1068_
timestamp 1688980957
transform 1 0 13800 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1069_
timestamp 1688980957
transform -1 0 16376 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1070_
timestamp 1688980957
transform 1 0 16284 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1071_
timestamp 1688980957
transform 1 0 16744 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1072_
timestamp 1688980957
transform -1 0 20608 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1073_
timestamp 1688980957
transform -1 0 20792 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1074_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22172 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_4  _1075_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19412 0 1 11424
box -38 -48 1418 592
use sky130_fd_sc_hd__mux4_1  _1076_
timestamp 1688980957
transform 1 0 25668 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1077_
timestamp 1688980957
transform -1 0 27784 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1078_
timestamp 1688980957
transform 1 0 27048 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1079_
timestamp 1688980957
transform 1 0 21068 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1080_
timestamp 1688980957
transform -1 0 23460 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1081_
timestamp 1688980957
transform 1 0 22540 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1082_
timestamp 1688980957
transform -1 0 25484 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1083_
timestamp 1688980957
transform -1 0 25760 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1084_
timestamp 1688980957
transform 1 0 24472 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1085_
timestamp 1688980957
transform 1 0 18584 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1086_
timestamp 1688980957
transform 1 0 20148 0 1 9248
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1087_
timestamp 1688980957
transform 1 0 20884 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1088_
timestamp 1688980957
transform 1 0 25484 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1089_
timestamp 1688980957
transform -1 0 28244 0 -1 7072
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1090_
timestamp 1688980957
transform -1 0 27048 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1091_
timestamp 1688980957
transform 1 0 15732 0 1 24480
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1092_
timestamp 1688980957
transform 1 0 20976 0 -1 19040
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1093_
timestamp 1688980957
transform 1 0 21436 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1094_
timestamp 1688980957
transform -1 0 24196 0 1 13600
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1095_
timestamp 1688980957
transform -1 0 24656 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1096_
timestamp 1688980957
transform 1 0 23460 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux4_1  _1097_
timestamp 1688980957
transform 1 0 5520 0 1 17952
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_1  _1098_
timestamp 1688980957
transform 1 0 19320 0 -1 17952
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1099_
timestamp 1688980957
transform 1 0 19780 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1100_
timestamp 1688980957
transform 1 0 21712 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1101_
timestamp 1688980957
transform -1 0 22356 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1102_
timestamp 1688980957
transform 1 0 20240 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _1103_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14444 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1104_
timestamp 1688980957
transform 1 0 18584 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1105_
timestamp 1688980957
transform 1 0 18768 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1106_
timestamp 1688980957
transform 1 0 8096 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1107_
timestamp 1688980957
transform 1 0 9108 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1108_
timestamp 1688980957
transform 1 0 3772 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1109_
timestamp 1688980957
transform 1 0 18400 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1110_
timestamp 1688980957
transform -1 0 18216 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1111_
timestamp 1688980957
transform 1 0 14812 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1112_
timestamp 1688980957
transform -1 0 24012 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1113_
timestamp 1688980957
transform -1 0 25392 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1114_
timestamp 1688980957
transform -1 0 8924 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1115_
timestamp 1688980957
transform 1 0 9844 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1116_
timestamp 1688980957
transform -1 0 6256 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1117_
timestamp 1688980957
transform 1 0 17296 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1118_
timestamp 1688980957
transform 1 0 5520 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1119_
timestamp 1688980957
transform -1 0 21712 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1120_
timestamp 1688980957
transform 1 0 3772 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1121_
timestamp 1688980957
transform 1 0 3864 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1122_
timestamp 1688980957
transform 1 0 18308 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1123_
timestamp 1688980957
transform 1 0 13708 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1124_
timestamp 1688980957
transform -1 0 25300 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1125_
timestamp 1688980957
transform 1 0 28612 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1126_
timestamp 1688980957
transform 1 0 5428 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1127_
timestamp 1688980957
transform -1 0 24196 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1128_
timestamp 1688980957
transform 1 0 8372 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1129_
timestamp 1688980957
transform -1 0 24288 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1130_
timestamp 1688980957
transform 1 0 27140 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1131_
timestamp 1688980957
transform -1 0 29256 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1132_
timestamp 1688980957
transform 1 0 16284 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1133_
timestamp 1688980957
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1134_
timestamp 1688980957
transform 1 0 5428 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1135_
timestamp 1688980957
transform 1 0 22172 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _1136_
timestamp 1688980957
transform 1 0 13156 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__and4b_1  _1137_
timestamp 1688980957
transform -1 0 18308 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1138_
timestamp 1688980957
transform -1 0 14904 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1139_
timestamp 1688980957
transform 1 0 15732 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1140_
timestamp 1688980957
transform -1 0 14536 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1141_
timestamp 1688980957
transform 1 0 14904 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1142_
timestamp 1688980957
transform -1 0 6992 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1143_
timestamp 1688980957
transform 1 0 7084 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1144_
timestamp 1688980957
transform 1 0 31464 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1145_
timestamp 1688980957
transform -1 0 13984 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1146_
timestamp 1688980957
transform 1 0 21528 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1147_
timestamp 1688980957
transform 1 0 3404 0 -1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1148_
timestamp 1688980957
transform 1 0 5428 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1149_
timestamp 1688980957
transform 1 0 32660 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1150_
timestamp 1688980957
transform 1 0 32660 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1151_
timestamp 1688980957
transform 1 0 30452 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1152_
timestamp 1688980957
transform -1 0 31280 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1153_
timestamp 1688980957
transform 1 0 29532 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1154_
timestamp 1688980957
transform -1 0 6256 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1155_
timestamp 1688980957
transform 1 0 33028 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1156_
timestamp 1688980957
transform 1 0 4508 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1157_
timestamp 1688980957
transform 1 0 32016 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1158_
timestamp 1688980957
transform 1 0 3772 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1159_
timestamp 1688980957
transform 1 0 3956 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1160_
timestamp 1688980957
transform 1 0 31188 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1161_
timestamp 1688980957
transform 1 0 3588 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1162_
timestamp 1688980957
transform -1 0 4784 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1163_
timestamp 1688980957
transform -1 0 23644 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1164_
timestamp 1688980957
transform 1 0 32108 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1165_
timestamp 1688980957
transform 1 0 32384 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1166_
timestamp 1688980957
transform -1 0 25944 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1167_
timestamp 1688980957
transform -1 0 32844 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1168_
timestamp 1688980957
transform -1 0 30268 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1169_
timestamp 1688980957
transform 1 0 31096 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1170_
timestamp 1688980957
transform -1 0 4232 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1171_
timestamp 1688980957
transform 1 0 32660 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1172_
timestamp 1688980957
transform 1 0 3680 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1173_
timestamp 1688980957
transform 1 0 4508 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _1174_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1175_
timestamp 1688980957
transform 1 0 18768 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1176_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1177_
timestamp 1688980957
transform -1 0 21620 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1178_
timestamp 1688980957
transform -1 0 14904 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__or3_2  _1179_
timestamp 1688980957
transform -1 0 18032 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1180_
timestamp 1688980957
transform -1 0 14904 0 1 14688
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1181_
timestamp 1688980957
transform -1 0 14628 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1182_
timestamp 1688980957
transform -1 0 26772 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1183_
timestamp 1688980957
transform 1 0 17572 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1184_
timestamp 1688980957
transform -1 0 14720 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1185_
timestamp 1688980957
transform 1 0 16468 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1186_
timestamp 1688980957
transform 1 0 17296 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__and4bb_1  _1187_
timestamp 1688980957
transform -1 0 17940 0 -1 17952
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _1188_
timestamp 1688980957
transform 1 0 12788 0 1 13600
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _1189_
timestamp 1688980957
transform -1 0 16928 0 1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _1190_
timestamp 1688980957
transform -1 0 19044 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1191_
timestamp 1688980957
transform 1 0 18400 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1192_
timestamp 1688980957
transform 1 0 17664 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1193_
timestamp 1688980957
transform 1 0 18308 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _1194_
timestamp 1688980957
transform 1 0 16928 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1195_
timestamp 1688980957
transform 1 0 16284 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1196_
timestamp 1688980957
transform 1 0 14904 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1197_
timestamp 1688980957
transform 1 0 14720 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _1198_
timestamp 1688980957
transform 1 0 11960 0 1 23392
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1199_
timestamp 1688980957
transform -1 0 12972 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _1200_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26680 0 1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1688980957
transform -1 0 20516 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1688980957
transform 1 0 18676 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1688980957
transform -1 0 24932 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1688980957
transform -1 0 13432 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1688980957
transform -1 0 23736 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1206_
timestamp 1688980957
transform -1 0 5428 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1207_
timestamp 1688980957
transform -1 0 5428 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1208_
timestamp 1688980957
transform 1 0 33764 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1209_
timestamp 1688980957
transform -1 0 3404 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1210_
timestamp 1688980957
transform -1 0 32568 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1211_
timestamp 1688980957
transform -1 0 31832 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1212_
timestamp 1688980957
transform 1 0 33764 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1213_
timestamp 1688980957
transform -1 0 27048 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1214_
timestamp 1688980957
transform 1 0 33764 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1215_
timestamp 1688980957
transform 1 0 33764 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1216_
timestamp 1688980957
transform -1 0 23920 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1217_
timestamp 1688980957
transform -1 0 4048 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1218_
timestamp 1688980957
transform 1 0 3312 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1688980957
transform 1 0 32016 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1220_
timestamp 1688980957
transform -1 0 5152 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1221_
timestamp 1688980957
transform -1 0 5152 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1222_
timestamp 1688980957
transform -1 0 33856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1223_
timestamp 1688980957
transform 1 0 3312 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1224_
timestamp 1688980957
transform 1 0 33764 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1688980957
transform -1 0 5152 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1226_
timestamp 1688980957
transform -1 0 30912 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1227_
timestamp 1688980957
transform -1 0 32200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1228_
timestamp 1688980957
transform -1 0 31464 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1229_
timestamp 1688980957
transform 1 0 33764 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1230_
timestamp 1688980957
transform 1 0 33764 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1231_
timestamp 1688980957
transform -1 0 7268 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1232_
timestamp 1688980957
transform -1 0 5152 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1233_
timestamp 1688980957
transform -1 0 22632 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1234_
timestamp 1688980957
transform -1 0 14996 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1235_
timestamp 1688980957
transform -1 0 33304 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1236_
timestamp 1688980957
transform -1 0 8280 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1237_
timestamp 1688980957
transform -1 0 7912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1238_
timestamp 1688980957
transform -1 0 23736 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1239_
timestamp 1688980957
transform -1 0 7268 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1240_
timestamp 1688980957
transform -1 0 14720 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1241_
timestamp 1688980957
transform -1 0 18124 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1242_
timestamp 1688980957
transform -1 0 31464 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1243_
timestamp 1688980957
transform -1 0 27968 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1244_
timestamp 1688980957
transform -1 0 24840 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1245_
timestamp 1688980957
transform -1 0 9384 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1246_
timestamp 1688980957
transform 1 0 23644 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1247_
timestamp 1688980957
transform -1 0 6532 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1248_
timestamp 1688980957
transform -1 0 29716 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1249_
timestamp 1688980957
transform -1 0 25576 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1250_
timestamp 1688980957
transform -1 0 15456 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1251_
timestamp 1688980957
transform -1 0 18860 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1252_
timestamp 1688980957
transform -1 0 5152 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1688980957
transform -1 0 4600 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1254_
timestamp 1688980957
transform -1 0 23276 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1688980957
transform -1 0 6992 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1256_
timestamp 1688980957
transform -1 0 18584 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1257_
timestamp 1688980957
transform 1 0 3496 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1258_
timestamp 1688980957
transform -1 0 10856 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1259_
timestamp 1688980957
transform 1 0 7636 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1260_
timestamp 1688980957
transform -1 0 26312 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1261_
timestamp 1688980957
transform -1 0 25024 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1262_
timestamp 1688980957
transform -1 0 17572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1263_
timestamp 1688980957
transform -1 0 18768 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1264_
timestamp 1688980957
transform 1 0 19044 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1265_
timestamp 1688980957
transform -1 0 5152 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1266_
timestamp 1688980957
transform -1 0 10212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1267_
timestamp 1688980957
transform -1 0 10764 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1268_
timestamp 1688980957
transform 1 0 17848 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1269_
timestamp 1688980957
transform -1 0 21160 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1270_
timestamp 1688980957
transform -1 0 23000 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1271_
timestamp 1688980957
transform -1 0 21160 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1272_
timestamp 1688980957
transform 1 0 23828 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1273_
timestamp 1688980957
transform -1 0 23368 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1274_
timestamp 1688980957
transform -1 0 27140 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1275_
timestamp 1688980957
transform 1 0 20516 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1276_
timestamp 1688980957
transform 1 0 25300 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1688980957
transform -1 0 23736 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1278_
timestamp 1688980957
transform -1 0 28888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1279_
timestamp 1688980957
transform 1 0 17388 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1280_
timestamp 1688980957
transform -1 0 18584 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1281_
timestamp 1688980957
transform 1 0 14812 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1282_
timestamp 1688980957
transform 1 0 15732 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1283_
timestamp 1688980957
transform 1 0 12788 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1284_
timestamp 1688980957
transform -1 0 14260 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1285_
timestamp 1688980957
transform -1 0 11960 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1688980957
transform -1 0 11684 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1287_
timestamp 1688980957
transform -1 0 6440 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1688980957
transform -1 0 3404 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 1688980957
transform 1 0 26772 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1290_
timestamp 1688980957
transform -1 0 7636 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1688980957
transform 1 0 31188 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1292_
timestamp 1688980957
transform 1 0 28704 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1688980957
transform -1 0 31740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1294_
timestamp 1688980957
transform -1 0 23276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1295_
timestamp 1688980957
transform -1 0 31740 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1296_
timestamp 1688980957
transform -1 0 9752 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1297_
timestamp 1688980957
transform -1 0 23184 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 1688980957
transform -1 0 18492 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1299_
timestamp 1688980957
transform -1 0 10120 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1688980957
transform 1 0 26680 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1301_
timestamp 1688980957
transform 1 0 5428 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 1688980957
transform -1 0 5704 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1688980957
transform 1 0 20516 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1688980957
transform -1 0 5704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1305_
timestamp 1688980957
transform -1 0 21160 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1306_
timestamp 1688980957
transform 1 0 5060 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1307_
timestamp 1688980957
transform 1 0 28612 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1688980957
transform -1 0 30268 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1309_
timestamp 1688980957
transform 1 0 28060 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1310_
timestamp 1688980957
transform 1 0 21988 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1311_
timestamp 1688980957
transform 1 0 20976 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1312_
timestamp 1688980957
transform -1 0 7820 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1313_
timestamp 1688980957
transform -1 0 19136 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1688980957
transform -1 0 21160 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1315_
timestamp 1688980957
transform -1 0 13432 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1316_
timestamp 1688980957
transform -1 0 21068 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1317_
timestamp 1688980957
transform -1 0 8280 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1318_
timestamp 1688980957
transform -1 0 9016 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1319_
timestamp 1688980957
transform -1 0 21160 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1688980957
transform -1 0 7912 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1321_
timestamp 1688980957
transform 1 0 14168 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1322_
timestamp 1688980957
transform -1 0 12328 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1323_
timestamp 1688980957
transform -1 0 28888 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1324_
timestamp 1688980957
transform 1 0 26864 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1325_
timestamp 1688980957
transform 1 0 23092 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1326_
timestamp 1688980957
transform -1 0 21160 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1688980957
transform -1 0 25300 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1328_
timestamp 1688980957
transform -1 0 8280 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1329_
timestamp 1688980957
transform -1 0 27692 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1330_
timestamp 1688980957
transform 1 0 24288 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1331_
timestamp 1688980957
transform -1 0 14720 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1332_
timestamp 1688980957
transform -1 0 19780 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1333_
timestamp 1688980957
transform 1 0 5888 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1334_
timestamp 1688980957
transform 1 0 5612 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1335_
timestamp 1688980957
transform -1 0 21160 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1336_
timestamp 1688980957
transform -1 0 6348 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1337_
timestamp 1688980957
transform -1 0 18952 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1338_
timestamp 1688980957
transform 1 0 5060 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1339_
timestamp 1688980957
transform 1 0 11316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1340_
timestamp 1688980957
transform -1 0 9660 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1341_
timestamp 1688980957
transform 1 0 23736 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1342_
timestamp 1688980957
transform 1 0 21896 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1343_
timestamp 1688980957
transform 1 0 15272 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1344_
timestamp 1688980957
transform -1 0 16836 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1345_
timestamp 1688980957
transform 1 0 18676 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1346_
timestamp 1688980957
transform 1 0 18308 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1347_
timestamp 1688980957
transform 1 0 31464 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1688980957
transform 1 0 13892 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1349_
timestamp 1688980957
transform 1 0 8740 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1350_
timestamp 1688980957
transform 1 0 8280 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1351_
timestamp 1688980957
transform 1 0 8188 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 1688980957
transform 1 0 9476 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1353_
timestamp 1688980957
transform -1 0 16652 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 1688980957
transform -1 0 15916 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1355_
timestamp 1688980957
transform -1 0 13800 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1356_
timestamp 1688980957
transform 1 0 16652 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1357_
timestamp 1688980957
transform -1 0 16928 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1688980957
transform -1 0 17296 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1359_
timestamp 1688980957
transform 1 0 15364 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1360_
timestamp 1688980957
transform -1 0 15640 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1361_
timestamp 1688980957
transform -1 0 10856 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1362_
timestamp 1688980957
transform -1 0 12604 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1363_
timestamp 1688980957
transform 1 0 11040 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1364_
timestamp 1688980957
transform -1 0 13432 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1365_
timestamp 1688980957
transform 1 0 8464 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1366_
timestamp 1688980957
transform 1 0 7636 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1367_
timestamp 1688980957
transform 1 0 7636 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1368_
timestamp 1688980957
transform 1 0 6900 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1369_
timestamp 1688980957
transform 1 0 15272 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1370_
timestamp 1688980957
transform -1 0 16008 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1371_
timestamp 1688980957
transform -1 0 16744 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1372_
timestamp 1688980957
transform -1 0 16008 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1373_
timestamp 1688980957
transform -1 0 12144 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1374_
timestamp 1688980957
transform -1 0 9752 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1375_
timestamp 1688980957
transform 1 0 10580 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1376_
timestamp 1688980957
transform -1 0 7084 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1377_
timestamp 1688980957
transform 1 0 13892 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1378_
timestamp 1688980957
transform 1 0 23736 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1379_
timestamp 1688980957
transform -1 0 25024 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1380_
timestamp 1688980957
transform 1 0 23828 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1381_
timestamp 1688980957
transform -1 0 26128 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1382_
timestamp 1688980957
transform -1 0 23276 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1383_
timestamp 1688980957
transform 1 0 25300 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1384_
timestamp 1688980957
transform 1 0 23092 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1385_
timestamp 1688980957
transform -1 0 30912 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1688980957
transform -1 0 31188 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1387_
timestamp 1688980957
transform -1 0 11684 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1388_
timestamp 1688980957
transform 1 0 28060 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1389_
timestamp 1688980957
transform -1 0 25300 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1390_
timestamp 1688980957
transform -1 0 25944 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1391_
timestamp 1688980957
transform 1 0 24932 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1392_
timestamp 1688980957
transform -1 0 25668 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1393_
timestamp 1688980957
transform -1 0 28888 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1394_
timestamp 1688980957
transform -1 0 30360 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1395_
timestamp 1688980957
transform -1 0 33396 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1396_
timestamp 1688980957
transform 1 0 30176 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1397_
timestamp 1688980957
transform -1 0 32660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1398_
timestamp 1688980957
transform 1 0 31924 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1399_
timestamp 1688980957
transform -1 0 32200 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1400_
timestamp 1688980957
transform 1 0 28612 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1401_
timestamp 1688980957
transform -1 0 31464 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1402_
timestamp 1688980957
transform 1 0 25668 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1403_
timestamp 1688980957
transform -1 0 28888 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1404_
timestamp 1688980957
transform 1 0 26036 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1405_
timestamp 1688980957
transform 1 0 23644 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1406_
timestamp 1688980957
transform -1 0 28336 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1407_
timestamp 1688980957
transform -1 0 29164 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1408_
timestamp 1688980957
transform -1 0 31464 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1409_
timestamp 1688980957
transform -1 0 32936 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1410_
timestamp 1688980957
transform -1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1411_
timestamp 1688980957
transform -1 0 13064 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1412_
timestamp 1688980957
transform 1 0 13616 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1413_
timestamp 1688980957
transform -1 0 14168 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1414_
timestamp 1688980957
transform 1 0 10212 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1415_
timestamp 1688980957
transform 1 0 7636 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1416_
timestamp 1688980957
transform 1 0 7636 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1417_
timestamp 1688980957
transform 1 0 8924 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1419_
timestamp 1688980957
transform 1 0 17664 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1420_
timestamp 1688980957
transform -1 0 20424 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1421_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25668 0 1 14688
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1422_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13984 0 1 14688
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _1423_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1424_
timestamp 1688980957
transform -1 0 5152 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1425_
timestamp 1688980957
transform -1 0 4876 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1426_
timestamp 1688980957
transform 1 0 32108 0 1 27744
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1427_
timestamp 1688980957
transform -1 0 4876 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1428_
timestamp 1688980957
transform 1 0 31188 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1429_
timestamp 1688980957
transform 1 0 28980 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1430_
timestamp 1688980957
transform 1 0 31740 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1431_
timestamp 1688980957
transform 1 0 25300 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1432_
timestamp 1688980957
transform 1 0 31832 0 1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1433_
timestamp 1688980957
transform 1 0 31832 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1434_
timestamp 1688980957
transform 1 0 22264 0 1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1435_
timestamp 1688980957
transform -1 0 4876 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1436_
timestamp 1688980957
transform -1 0 4876 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1437_
timestamp 1688980957
transform 1 0 31004 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1438_
timestamp 1688980957
transform -1 0 4876 0 -1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1439_
timestamp 1688980957
transform 1 0 3036 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1440_
timestamp 1688980957
transform 1 0 31740 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1441_
timestamp 1688980957
transform -1 0 4876 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1442_
timestamp 1688980957
transform 1 0 31832 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1443_
timestamp 1688980957
transform -1 0 4876 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1444_
timestamp 1688980957
transform 1 0 29256 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1445_
timestamp 1688980957
transform 1 0 30084 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1446_
timestamp 1688980957
transform 1 0 29256 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1447_
timestamp 1688980957
transform 1 0 32200 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1448_
timestamp 1688980957
transform 1 0 31832 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1449_
timestamp 1688980957
transform -1 0 6348 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1450_
timestamp 1688980957
transform -1 0 4876 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1451_
timestamp 1688980957
transform 1 0 21252 0 1 25568
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1452_
timestamp 1688980957
transform -1 0 14996 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1453_
timestamp 1688980957
transform 1 0 31188 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1454_
timestamp 1688980957
transform 1 0 6072 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1455_
timestamp 1688980957
transform -1 0 7268 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1456_
timestamp 1688980957
transform 1 0 21896 0 1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1457_
timestamp 1688980957
transform -1 0 6348 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1458_
timestamp 1688980957
transform 1 0 11500 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1459_
timestamp 1688980957
transform 1 0 16008 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1460_
timestamp 1688980957
transform 1 0 28612 0 -1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1461_
timestamp 1688980957
transform 1 0 26496 0 1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1462_
timestamp 1688980957
transform -1 0 25576 0 -1 28832
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1463_
timestamp 1688980957
transform 1 0 8004 0 -1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1464_
timestamp 1688980957
transform -1 0 25300 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1465_
timestamp 1688980957
transform -1 0 6256 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1466_
timestamp 1688980957
transform 1 0 27692 0 1 3808
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1467_
timestamp 1688980957
transform 1 0 24104 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1468_
timestamp 1688980957
transform 1 0 13340 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1469_
timestamp 1688980957
transform 1 0 17572 0 1 32096
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1470_
timestamp 1688980957
transform 1 0 3036 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1471_
timestamp 1688980957
transform 1 0 3036 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1472_
timestamp 1688980957
transform -1 0 22264 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1473_
timestamp 1688980957
transform 1 0 4876 0 -1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1474_
timestamp 1688980957
transform 1 0 16560 0 1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1475_
timestamp 1688980957
transform -1 0 4876 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1476_
timestamp 1688980957
transform -1 0 10488 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1477_
timestamp 1688980957
transform -1 0 9844 0 -1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1478_
timestamp 1688980957
transform 1 0 24012 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1479_
timestamp 1688980957
transform 1 0 23460 0 -1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1480_
timestamp 1688980957
transform 1 0 14720 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1481_
timestamp 1688980957
transform 1 0 18308 0 -1 27744
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1482_
timestamp 1688980957
transform 1 0 18308 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1483_
timestamp 1688980957
transform 1 0 3036 0 1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1484_
timestamp 1688980957
transform 1 0 8280 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1485_
timestamp 1688980957
transform 1 0 7360 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1486_
timestamp 1688980957
transform 1 0 16928 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1487_
timestamp 1688980957
transform 1 0 18308 0 -1 21216
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1488_
timestamp 1688980957
transform 1 0 20884 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1489_
timestamp 1688980957
transform 1 0 18952 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1490_
timestamp 1688980957
transform 1 0 23368 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1491_
timestamp 1688980957
transform 1 0 21252 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1492_
timestamp 1688980957
transform -1 0 27876 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1493_
timestamp 1688980957
transform 1 0 20424 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1494_
timestamp 1688980957
transform 1 0 23828 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1495_
timestamp 1688980957
transform 1 0 21528 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1496_
timestamp 1688980957
transform 1 0 26956 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1497_
timestamp 1688980957
transform 1 0 16376 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1498_
timestamp 1688980957
transform 1 0 15732 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1499_
timestamp 1688980957
transform 1 0 15732 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1500_
timestamp 1688980957
transform 1 0 13156 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1501_
timestamp 1688980957
transform 1 0 11960 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1502_
timestamp 1688980957
transform 1 0 11408 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1503_
timestamp 1688980957
transform 1 0 10212 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1504_
timestamp 1688980957
transform 1 0 10396 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1505_
timestamp 1688980957
transform 1 0 4232 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1506_
timestamp 1688980957
transform -1 0 4876 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1507_
timestamp 1688980957
transform 1 0 26036 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1508_
timestamp 1688980957
transform -1 0 7912 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1509_
timestamp 1688980957
transform 1 0 29164 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1510_
timestamp 1688980957
transform 1 0 27692 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1511_
timestamp 1688980957
transform 1 0 29624 0 -1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1512_
timestamp 1688980957
transform 1 0 21160 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1513_
timestamp 1688980957
transform -1 0 31648 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1514_
timestamp 1688980957
transform 1 0 8372 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1515_
timestamp 1688980957
transform 1 0 21252 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1516_
timestamp 1688980957
transform -1 0 18216 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1517_
timestamp 1688980957
transform -1 0 10672 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1518_
timestamp 1688980957
transform 1 0 25576 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1519_
timestamp 1688980957
transform -1 0 6808 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1520_
timestamp 1688980957
transform -1 0 6440 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1521_
timestamp 1688980957
transform 1 0 19688 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1522_
timestamp 1688980957
transform 1 0 4232 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1523_
timestamp 1688980957
transform 1 0 18952 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1524_
timestamp 1688980957
transform 1 0 4048 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1525_
timestamp 1688980957
transform 1 0 27600 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1526_
timestamp 1688980957
transform 1 0 28612 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1527_
timestamp 1688980957
transform 1 0 28612 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1528_
timestamp 1688980957
transform 1 0 21068 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1529_
timestamp 1688980957
transform 1 0 19964 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1530_
timestamp 1688980957
transform 1 0 5704 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1531_
timestamp 1688980957
transform -1 0 20148 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1532_
timestamp 1688980957
transform 1 0 19688 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1533_
timestamp 1688980957
transform 1 0 11224 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1534_
timestamp 1688980957
transform 1 0 18952 0 -1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1535_
timestamp 1688980957
transform 1 0 6900 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1536_
timestamp 1688980957
transform -1 0 8096 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1537_
timestamp 1688980957
transform -1 0 21804 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1538_
timestamp 1688980957
transform 1 0 5060 0 -1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1539_
timestamp 1688980957
transform 1 0 13156 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1540_
timestamp 1688980957
transform 1 0 10580 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1541_
timestamp 1688980957
transform 1 0 27324 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1542_
timestamp 1688980957
transform 1 0 25852 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1543_
timestamp 1688980957
transform 1 0 22540 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1544_
timestamp 1688980957
transform -1 0 22080 0 -1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1545_
timestamp 1688980957
transform 1 0 22540 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1546_
timestamp 1688980957
transform -1 0 8556 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1547_
timestamp 1688980957
transform -1 0 28520 0 1 4896
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1548_
timestamp 1688980957
transform 1 0 23460 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1549_
timestamp 1688980957
transform 1 0 11868 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1550_
timestamp 1688980957
transform 1 0 17664 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1551_
timestamp 1688980957
transform -1 0 7268 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1552_
timestamp 1688980957
transform -1 0 7268 0 1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1553_
timestamp 1688980957
transform 1 0 19044 0 -1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1554_
timestamp 1688980957
transform 1 0 4232 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1555_
timestamp 1688980957
transform 1 0 16376 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1556_
timestamp 1688980957
transform 1 0 4416 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1557_
timestamp 1688980957
transform 1 0 9200 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1558_
timestamp 1688980957
transform 1 0 7544 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1559_
timestamp 1688980957
transform 1 0 23460 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1560_
timestamp 1688980957
transform 1 0 20976 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1561_
timestamp 1688980957
transform 1 0 14260 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1562_
timestamp 1688980957
transform 1 0 14720 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1563_
timestamp 1688980957
transform 1 0 18308 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1564_
timestamp 1688980957
transform 1 0 17020 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1565_
timestamp 1688980957
transform 1 0 31188 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1566_
timestamp 1688980957
transform 1 0 13156 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1567_
timestamp 1688980957
transform 1 0 7912 0 1 29920
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1568_
timestamp 1688980957
transform 1 0 7452 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1569_
timestamp 1688980957
transform 1 0 7268 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1570_
timestamp 1688980957
transform 1 0 8556 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1571_
timestamp 1688980957
transform -1 0 17664 0 1 26656
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1572_
timestamp 1688980957
transform 1 0 13800 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1573_
timestamp 1688980957
transform 1 0 11684 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1574_
timestamp 1688980957
transform 1 0 15732 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1575_
timestamp 1688980957
transform 1 0 14812 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1576_
timestamp 1688980957
transform 1 0 15824 0 1 28832
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1577_
timestamp 1688980957
transform -1 0 17572 0 1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1578_
timestamp 1688980957
transform 1 0 13524 0 1 33184
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1579_
timestamp 1688980957
transform 1 0 8648 0 1 33184
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1580_
timestamp 1688980957
transform -1 0 13064 0 1 33184
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1581_
timestamp 1688980957
transform 1 0 9200 0 -1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1582_
timestamp 1688980957
transform 1 0 11960 0 1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1583_
timestamp 1688980957
transform 1 0 8004 0 -1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1584_
timestamp 1688980957
transform 1 0 8004 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1585_
timestamp 1688980957
transform 1 0 6716 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1586_
timestamp 1688980957
transform 1 0 5980 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1587_
timestamp 1688980957
transform 1 0 14260 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1588_
timestamp 1688980957
transform -1 0 15640 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1589_
timestamp 1688980957
transform 1 0 14904 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1590_
timestamp 1688980957
transform 1 0 14444 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1591_
timestamp 1688980957
transform -1 0 12788 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1592_
timestamp 1688980957
transform 1 0 8004 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1593_
timestamp 1688980957
transform -1 0 10488 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1594_
timestamp 1688980957
transform -1 0 7544 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1595_
timestamp 1688980957
transform 1 0 13156 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1596_
timestamp 1688980957
transform 1 0 22724 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1597_
timestamp 1688980957
transform 1 0 22908 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1598_
timestamp 1688980957
transform 1 0 23460 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1599_
timestamp 1688980957
transform -1 0 27876 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1600_
timestamp 1688980957
transform 1 0 21344 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1601_
timestamp 1688980957
transform 1 0 23828 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1602_
timestamp 1688980957
transform 1 0 23184 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1603_
timestamp 1688980957
transform -1 0 30452 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1604_
timestamp 1688980957
transform 1 0 29072 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _1605_
timestamp 1688980957
transform -1 0 12328 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1606_
timestamp 1688980957
transform 1 0 27048 0 1 14688
box -38 -48 2154 592
use sky130_fd_sc_hd__dfstp_1  _1607_
timestamp 1688980957
transform -1 0 26036 0 -1 16864
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1608_
timestamp 1688980957
transform 1 0 26036 0 1 24480
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1609_
timestamp 1688980957
transform 1 0 24012 0 1 23392
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1610_
timestamp 1688980957
transform 1 0 24012 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1611_
timestamp 1688980957
transform -1 0 28520 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1612_
timestamp 1688980957
transform 1 0 28980 0 1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1613_
timestamp 1688980957
transform -1 0 33120 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1614_
timestamp 1688980957
transform 1 0 29256 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1615_
timestamp 1688980957
transform 1 0 30544 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1616_
timestamp 1688980957
transform -1 0 33028 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1617_
timestamp 1688980957
transform -1 0 33028 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1618_
timestamp 1688980957
transform 1 0 27692 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1619_
timestamp 1688980957
transform 1 0 29992 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1620_
timestamp 1688980957
transform 1 0 24288 0 -1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1621_
timestamp 1688980957
transform 1 0 25944 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1622_
timestamp 1688980957
transform 1 0 24104 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1623_
timestamp 1688980957
transform -1 0 25300 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1624_
timestamp 1688980957
transform 1 0 26772 0 1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1625_
timestamp 1688980957
transform 1 0 27140 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1626_
timestamp 1688980957
transform -1 0 32108 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1627_
timestamp 1688980957
transform -1 0 32660 0 -1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1628_
timestamp 1688980957
transform 1 0 11776 0 1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1629_
timestamp 1688980957
transform 1 0 11684 0 1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1630_
timestamp 1688980957
transform 1 0 12696 0 1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1631_
timestamp 1688980957
transform 1 0 12236 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1632_
timestamp 1688980957
transform 1 0 10580 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1633_
timestamp 1688980957
transform 1 0 6716 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1634_
timestamp 1688980957
transform 1 0 6900 0 1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1635_
timestamp 1688980957
transform 1 0 6072 0 -1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  _1636_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13432 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15364 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A0
timestamp 1688980957
transform 1 0 12236 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A
timestamp 1688980957
transform 1 0 12880 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__B
timestamp 1688980957
transform 1 0 14260 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__C
timestamp 1688980957
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A_N
timestamp 1688980957
transform 1 0 16652 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A1
timestamp 1688980957
transform 1 0 17388 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A_N
timestamp 1688980957
transform 1 0 18492 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__C
timestamp 1688980957
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__D
timestamp 1688980957
transform 1 0 17664 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1688980957
transform 1 0 16468 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A2
timestamp 1688980957
transform 1 0 17756 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1688980957
transform 1 0 15364 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__B
timestamp 1688980957
transform -1 0 15640 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A0
timestamp 1688980957
transform 1 0 16928 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1688980957
transform 1 0 15916 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A0
timestamp 1688980957
transform 1 0 15916 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__C
timestamp 1688980957
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__C
timestamp 1688980957
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A2_N
timestamp 1688980957
transform 1 0 22632 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1688980957
transform 1 0 19688 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 1688980957
transform 1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__C_N
timestamp 1688980957
transform 1 0 17664 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1_N
timestamp 1688980957
transform -1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A2_N
timestamp 1688980957
transform -1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__B2
timestamp 1688980957
transform 1 0 22356 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A
timestamp 1688980957
transform 1 0 9936 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B
timestamp 1688980957
transform 1 0 10120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__C_N
timestamp 1688980957
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1_N
timestamp 1688980957
transform -1 0 7912 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A2_N
timestamp 1688980957
transform -1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B2
timestamp 1688980957
transform 1 0 8924 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1688980957
transform 1 0 9568 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__B
timestamp 1688980957
transform 1 0 12328 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A1_N
timestamp 1688980957
transform 1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B2
timestamp 1688980957
transform 1 0 10948 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1688980957
transform 1 0 6348 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B
timestamp 1688980957
transform 1 0 6532 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__C_N
timestamp 1688980957
transform 1 0 6716 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1_N
timestamp 1688980957
transform 1 0 8556 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B2
timestamp 1688980957
transform 1 0 8464 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__B
timestamp 1688980957
transform 1 0 17664 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A1_N
timestamp 1688980957
transform 1 0 16468 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1688980957
transform 1 0 9936 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__B
timestamp 1688980957
transform 1 0 9016 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__C_N
timestamp 1688980957
transform 1 0 9476 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1_N
timestamp 1688980957
transform 1 0 6532 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__B2
timestamp 1688980957
transform 1 0 6992 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1688980957
transform -1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B
timestamp 1688980957
transform 1 0 18032 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A1_N
timestamp 1688980957
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B2
timestamp 1688980957
transform 1 0 20516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A_N
timestamp 1688980957
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B
timestamp 1688980957
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A
timestamp 1688980957
transform 1 0 10304 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A2
timestamp 1688980957
transform -1 0 3496 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B1
timestamp 1688980957
transform 1 0 5060 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A_N
timestamp 1688980957
transform 1 0 6716 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B
timestamp 1688980957
transform 1 0 7360 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__C
timestamp 1688980957
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A
timestamp 1688980957
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A2
timestamp 1688980957
transform 1 0 6716 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B1
timestamp 1688980957
transform 1 0 4784 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B
timestamp 1688980957
transform 1 0 17388 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__C
timestamp 1688980957
transform 1 0 17204 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A
timestamp 1688980957
transform 1 0 18492 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B1
timestamp 1688980957
transform 1 0 18032 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A_N
timestamp 1688980957
transform 1 0 11132 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B
timestamp 1688980957
transform 1 0 11500 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1688980957
transform 1 0 12328 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A2
timestamp 1688980957
transform 1 0 12420 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B1
timestamp 1688980957
transform 1 0 12236 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A_N
timestamp 1688980957
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__B
timestamp 1688980957
transform 1 0 17020 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__C
timestamp 1688980957
transform -1 0 19044 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A
timestamp 1688980957
transform 1 0 17848 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__B1
timestamp 1688980957
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B
timestamp 1688980957
transform 1 0 18032 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A
timestamp 1688980957
transform 1 0 18860 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A2
timestamp 1688980957
transform 1 0 27968 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__B1
timestamp 1688980957
transform 1 0 25760 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__B2
timestamp 1688980957
transform -1 0 30176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A_N
timestamp 1688980957
transform 1 0 7360 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__B
timestamp 1688980957
transform 1 0 7452 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__C
timestamp 1688980957
transform 1 0 7452 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1688980957
transform 1 0 8648 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1688980957
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B1
timestamp 1688980957
transform 1 0 5152 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A_N
timestamp 1688980957
transform 1 0 20332 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1688980957
transform 1 0 19504 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A2
timestamp 1688980957
transform -1 0 23276 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B1
timestamp 1688980957
transform 1 0 23276 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B
timestamp 1688980957
transform 1 0 22264 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B1
timestamp 1688980957
transform -1 0 20792 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1688980957
transform 1 0 24288 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B
timestamp 1688980957
transform 1 0 23644 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B1
timestamp 1688980957
transform 1 0 22816 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B2
timestamp 1688980957
transform -1 0 22540 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1688980957
transform 1 0 26496 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1688980957
transform -1 0 27140 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A2
timestamp 1688980957
transform -1 0 26588 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__B1
timestamp 1688980957
transform -1 0 27508 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B
timestamp 1688980957
transform -1 0 28520 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A2
timestamp 1688980957
transform -1 0 27692 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__B1
timestamp 1688980957
transform -1 0 28428 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B
timestamp 1688980957
transform 1 0 7360 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A2
timestamp 1688980957
transform 1 0 12236 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__B1
timestamp 1688980957
transform -1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B
timestamp 1688980957
transform 1 0 19780 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A2
timestamp 1688980957
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B1
timestamp 1688980957
transform -1 0 13064 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B2
timestamp 1688980957
transform -1 0 13340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__B
timestamp 1688980957
transform 1 0 6624 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A2
timestamp 1688980957
transform 1 0 7544 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B1
timestamp 1688980957
transform 1 0 7452 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B
timestamp 1688980957
transform -1 0 18952 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B1
timestamp 1688980957
transform 1 0 19780 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B2
timestamp 1688980957
transform 1 0 19780 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B
timestamp 1688980957
transform 1 0 18400 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__C
timestamp 1688980957
transform 1 0 18768 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1688980957
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C
timestamp 1688980957
transform 1 0 20240 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A2
timestamp 1688980957
transform 1 0 8924 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__B2
timestamp 1688980957
transform -1 0 9476 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A2
timestamp 1688980957
transform 1 0 6348 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B2
timestamp 1688980957
transform -1 0 5888 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B2
timestamp 1688980957
transform -1 0 19688 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A2
timestamp 1688980957
transform 1 0 11592 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__B2
timestamp 1688980957
transform -1 0 11224 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B2
timestamp 1688980957
transform -1 0 19872 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B2
timestamp 1688980957
transform 1 0 19136 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1688980957
transform 1 0 7636 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B2
timestamp 1688980957
transform 1 0 5888 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B2
timestamp 1688980957
transform 1 0 19412 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A2_N
timestamp 1688980957
transform 1 0 22264 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1_N
timestamp 1688980957
transform -1 0 28244 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A2_N
timestamp 1688980957
transform 1 0 28704 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B2
timestamp 1688980957
transform 1 0 26680 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A1_N
timestamp 1688980957
transform -1 0 30636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A2_N
timestamp 1688980957
transform -1 0 30084 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B2
timestamp 1688980957
transform -1 0 30544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A2_N
timestamp 1688980957
transform -1 0 29256 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B2
timestamp 1688980957
transform 1 0 28152 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A2_N
timestamp 1688980957
transform 1 0 7820 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__B2
timestamp 1688980957
transform 1 0 6808 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A2_N
timestamp 1688980957
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A2_N
timestamp 1688980957
transform 1 0 7268 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B2
timestamp 1688980957
transform 1 0 7728 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A2_N
timestamp 1688980957
transform 1 0 21620 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B2
timestamp 1688980957
transform -1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A2
timestamp 1688980957
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__B2
timestamp 1688980957
transform 1 0 9568 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A2
timestamp 1688980957
transform 1 0 8188 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B2
timestamp 1688980957
transform 1 0 9936 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A2
timestamp 1688980957
transform 1 0 25668 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__B2
timestamp 1688980957
transform 1 0 27140 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A2
timestamp 1688980957
transform 1 0 10304 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__B2
timestamp 1688980957
transform 1 0 9844 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A2
timestamp 1688980957
transform 1 0 16928 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B2
timestamp 1688980957
transform 1 0 17296 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B1
timestamp 1688980957
transform 1 0 22264 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B2
timestamp 1688980957
transform 1 0 21896 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1
timestamp 1688980957
transform -1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A2
timestamp 1688980957
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B2
timestamp 1688980957
transform 1 0 9200 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A2
timestamp 1688980957
transform 1 0 29808 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B2
timestamp 1688980957
transform 1 0 29440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A2
timestamp 1688980957
transform 1 0 19596 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B2
timestamp 1688980957
transform 1 0 23000 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A2
timestamp 1688980957
transform 1 0 29808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__B1
timestamp 1688980957
transform -1 0 30728 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__B2
timestamp 1688980957
transform -1 0 30360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B2
timestamp 1688980957
transform -1 0 27876 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A2
timestamp 1688980957
transform 1 0 29624 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B2
timestamp 1688980957
transform -1 0 29256 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A2
timestamp 1688980957
transform 1 0 6992 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B2
timestamp 1688980957
transform 1 0 7360 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B1
timestamp 1688980957
transform -1 0 27692 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B2
timestamp 1688980957
transform 1 0 27324 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B2
timestamp 1688980957
transform -1 0 5336 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A2
timestamp 1688980957
transform -1 0 6624 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B1
timestamp 1688980957
transform -1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B2
timestamp 1688980957
transform -1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__S
timestamp 1688980957
transform 1 0 11500 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A0
timestamp 1688980957
transform 1 0 11868 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__S
timestamp 1688980957
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A0
timestamp 1688980957
transform 1 0 12696 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__S
timestamp 1688980957
transform 1 0 12880 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__S
timestamp 1688980957
transform 1 0 12236 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A0
timestamp 1688980957
transform 1 0 13616 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__S
timestamp 1688980957
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A0
timestamp 1688980957
transform 1 0 16192 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__S
timestamp 1688980957
transform 1 0 16928 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__S
timestamp 1688980957
transform 1 0 16560 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1688980957
transform -1 0 22724 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A1
timestamp 1688980957
transform -1 0 26404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__S0
timestamp 1688980957
transform 1 0 25208 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__S1
timestamp 1688980957
transform 1 0 25576 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A0
timestamp 1688980957
transform -1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__S0
timestamp 1688980957
transform 1 0 22264 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__S1
timestamp 1688980957
transform 1 0 18860 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A1
timestamp 1688980957
transform -1 0 25668 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__S0
timestamp 1688980957
transform 1 0 22724 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__S1
timestamp 1688980957
transform -1 0 23092 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A2
timestamp 1688980957
transform -1 0 20700 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__S0
timestamp 1688980957
transform 1 0 18492 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__S1
timestamp 1688980957
transform 1 0 18400 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A0
timestamp 1688980957
transform -1 0 26404 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A1
timestamp 1688980957
transform -1 0 26128 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A2
timestamp 1688980957
transform -1 0 28244 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__S0
timestamp 1688980957
transform 1 0 25484 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__S1
timestamp 1688980957
transform -1 0 26404 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A0
timestamp 1688980957
transform -1 0 15640 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__S0
timestamp 1688980957
transform 1 0 18308 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__S1
timestamp 1688980957
transform 1 0 19228 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A2
timestamp 1688980957
transform -1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__S0
timestamp 1688980957
transform 1 0 19872 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__S1
timestamp 1688980957
transform 1 0 23184 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A0
timestamp 1688980957
transform -1 0 5336 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__S0
timestamp 1688980957
transform 1 0 7820 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__S1
timestamp 1688980957
transform 1 0 7636 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A
timestamp 1688980957
transform 1 0 20056 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__B
timestamp 1688980957
transform 1 0 21344 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__C
timestamp 1688980957
transform 1 0 20608 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__B
timestamp 1688980957
transform 1 0 15456 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__S
timestamp 1688980957
transform 1 0 18032 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A0
timestamp 1688980957
transform -1 0 18584 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__S
timestamp 1688980957
transform 1 0 18584 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A0
timestamp 1688980957
transform 1 0 9108 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__S
timestamp 1688980957
transform 1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__S
timestamp 1688980957
transform 1 0 10764 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A0
timestamp 1688980957
transform -1 0 5152 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__S
timestamp 1688980957
transform -1 0 3772 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__S
timestamp 1688980957
transform 1 0 18216 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A0
timestamp 1688980957
transform -1 0 17940 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__S
timestamp 1688980957
transform 1 0 17204 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__S
timestamp 1688980957
transform 1 0 16468 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__S
timestamp 1688980957
transform 1 0 23000 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__S
timestamp 1688980957
transform 1 0 24380 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__S
timestamp 1688980957
transform -1 0 9108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__S
timestamp 1688980957
transform 1 0 10304 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__S
timestamp 1688980957
transform 1 0 7176 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__S
timestamp 1688980957
transform 1 0 17112 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__S
timestamp 1688980957
transform 1 0 6532 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__S
timestamp 1688980957
transform 1 0 20608 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__S
timestamp 1688980957
transform -1 0 3772 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__S
timestamp 1688980957
transform 1 0 4692 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__S
timestamp 1688980957
transform 1 0 19320 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__S
timestamp 1688980957
transform -1 0 14720 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__S
timestamp 1688980957
transform 1 0 23184 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__S
timestamp 1688980957
transform -1 0 28980 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__S
timestamp 1688980957
transform 1 0 5888 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__S
timestamp 1688980957
transform 1 0 23184 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__S
timestamp 1688980957
transform 1 0 10028 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__S
timestamp 1688980957
transform 1 0 22908 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__S
timestamp 1688980957
transform 1 0 26956 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__S
timestamp 1688980957
transform 1 0 28244 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__S
timestamp 1688980957
transform -1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__S
timestamp 1688980957
transform 1 0 14720 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__S
timestamp 1688980957
transform 1 0 6256 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__S
timestamp 1688980957
transform 1 0 21988 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__S
timestamp 1688980957
transform 1 0 7176 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__S
timestamp 1688980957
transform 1 0 8832 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__S
timestamp 1688980957
transform 1 0 32476 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__S
timestamp 1688980957
transform 1 0 12972 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__S
timestamp 1688980957
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__S
timestamp 1688980957
transform 1 0 6900 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__S
timestamp 1688980957
transform 1 0 5152 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__S
timestamp 1688980957
transform -1 0 34040 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__S
timestamp 1688980957
transform 1 0 32384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__S
timestamp 1688980957
transform 1 0 31464 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__S
timestamp 1688980957
transform 1 0 31464 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__S
timestamp 1688980957
transform 1 0 30360 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__S
timestamp 1688980957
transform 1 0 6440 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__S
timestamp 1688980957
transform 1 0 31740 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__S
timestamp 1688980957
transform 1 0 5152 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__S
timestamp 1688980957
transform 1 0 33304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__S
timestamp 1688980957
transform 1 0 3680 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__S
timestamp 1688980957
transform 1 0 3772 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__S
timestamp 1688980957
transform 1 0 32016 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__S
timestamp 1688980957
transform -1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__S
timestamp 1688980957
transform 1 0 4968 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__S
timestamp 1688980957
transform 1 0 24012 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A0
timestamp 1688980957
transform 1 0 31924 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__S
timestamp 1688980957
transform 1 0 33396 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__S
timestamp 1688980957
transform 1 0 33396 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__S
timestamp 1688980957
transform -1 0 26128 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__S
timestamp 1688980957
transform 1 0 32016 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__S
timestamp 1688980957
transform -1 0 30820 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__S
timestamp 1688980957
transform -1 0 31832 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__S
timestamp 1688980957
transform 1 0 8188 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__S
timestamp 1688980957
transform -1 0 33672 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__S
timestamp 1688980957
transform 1 0 3496 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__S
timestamp 1688980957
transform -1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__B1_N
timestamp 1688980957
transform 1 0 19228 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A0
timestamp 1688980957
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__B1_N
timestamp 1688980957
transform 1 0 14168 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B
timestamp 1688980957
transform 1 0 16744 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A2
timestamp 1688980957
transform -1 0 20056 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A1
timestamp 1688980957
transform 1 0 14904 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A2
timestamp 1688980957
transform -1 0 14168 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__A
timestamp 1688980957
transform 1 0 9844 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__A
timestamp 1688980957
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_0_clk_A
timestamp 1688980957
transform 1 0 8188 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_1_clk_A
timestamp 1688980957
transform 1 0 9936 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_2_clk_A
timestamp 1688980957
transform 1 0 11500 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_3_clk_A
timestamp 1688980957
transform 1 0 13432 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_4_clk_A
timestamp 1688980957
transform 1 0 9384 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_5_clk_A
timestamp 1688980957
transform 1 0 5980 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_6_clk_A
timestamp 1688980957
transform 1 0 7820 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_7_clk_A
timestamp 1688980957
transform 1 0 10028 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_8_clk_A
timestamp 1688980957
transform 1 0 15180 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_9_clk_A
timestamp 1688980957
transform -1 0 16008 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_10_clk_A
timestamp 1688980957
transform 1 0 22448 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_11_clk_A
timestamp 1688980957
transform 1 0 22724 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_12_clk_A
timestamp 1688980957
transform -1 0 28980 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_13_clk_A
timestamp 1688980957
transform 1 0 29348 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_14_clk_A
timestamp 1688980957
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_15_clk_A
timestamp 1688980957
transform 1 0 23184 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_16_clk_A
timestamp 1688980957
transform 1 0 27140 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_17_clk_A
timestamp 1688980957
transform -1 0 32568 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_18_clk_A
timestamp 1688980957
transform 1 0 31372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_19_clk_A
timestamp 1688980957
transform -1 0 30912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_20_clk_A
timestamp 1688980957
transform 1 0 23644 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_21_clk_A
timestamp 1688980957
transform 1 0 22632 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_22_clk_A
timestamp 1688980957
transform 1 0 24012 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_23_clk_A
timestamp 1688980957
transform -1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_24_clk_A
timestamp 1688980957
transform 1 0 12972 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_25_clk_A
timestamp 1688980957
transform 1 0 13616 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_26_clk_A
timestamp 1688980957
transform 1 0 10764 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_leaf_27_clk_A
timestamp 1688980957
transform 1 0 5612 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1688980957
transform -1 0 33212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1688980957
transform 1 0 14536 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 1688980957
transform 1 0 17296 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout108_A
timestamp 1688980957
transform -1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout109_A
timestamp 1688980957
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout110_A
timestamp 1688980957
transform 1 0 16468 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout111_A
timestamp 1688980957
transform 1 0 15364 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout113_A
timestamp 1688980957
transform 1 0 20884 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout117_A
timestamp 1688980957
transform 1 0 16836 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout119_A
timestamp 1688980957
transform 1 0 7544 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout120_A
timestamp 1688980957
transform 1 0 4692 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout121_A
timestamp 1688980957
transform 1 0 15456 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout122_A
timestamp 1688980957
transform 1 0 12880 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout126_A
timestamp 1688980957
transform 1 0 7176 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout127_A
timestamp 1688980957
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout128_A
timestamp 1688980957
transform 1 0 20424 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout130_A
timestamp 1688980957
transform 1 0 26956 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout134_A
timestamp 1688980957
transform 1 0 18032 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold115_A
timestamp 1688980957
transform 1 0 9476 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold165_A
timestamp 1688980957
transform -1 0 12788 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold173_A
timestamp 1688980957
transform 1 0 18676 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold204_A
timestamp 1688980957
transform 1 0 23644 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output99_A
timestamp 1688980957
transform -1 0 5152 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 1 19040
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1688980957
transform -1 0 12236 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1688980957
transform 1 0 20884 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_0_clk
timestamp 1688980957
transform 1 0 6072 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_1_clk
timestamp 1688980957
transform 1 0 5704 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_2_clk
timestamp 1688980957
transform 1 0 11316 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_3_clk
timestamp 1688980957
transform 1 0 14168 0 -1 20128
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_4_clk
timestamp 1688980957
transform -1 0 9200 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_5_clk
timestamp 1688980957
transform 1 0 4140 0 -1 23392
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_6_clk
timestamp 1688980957
transform 1 0 5612 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_7_clk
timestamp 1688980957
transform 1 0 7728 0 1 31008
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_8_clk
timestamp 1688980957
transform 1 0 15364 0 -1 32096
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_9_clk
timestamp 1688980957
transform 1 0 15732 0 1 25568
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_10_clk
timestamp 1688980957
transform 1 0 20608 0 -1 24480
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_11_clk
timestamp 1688980957
transform 1 0 22908 0 1 27744
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_12_clk
timestamp 1688980957
transform 1 0 29256 0 -1 29920
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_13_clk
timestamp 1688980957
transform 1 0 30360 0 -1 22304
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_14_clk
timestamp 1688980957
transform 1 0 23552 0 1 21216
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_15_clk
timestamp 1688980957
transform 1 0 21344 0 -1 17952
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_16_clk
timestamp 1688980957
transform 1 0 27324 0 1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_17_clk
timestamp 1688980957
transform 1 0 31832 0 -1 15776
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_18_clk
timestamp 1688980957
transform 1 0 30452 0 -1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_19_clk
timestamp 1688980957
transform 1 0 28612 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_20_clk
timestamp 1688980957
transform 1 0 23460 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_21_clk
timestamp 1688980957
transform 1 0 19872 0 -1 8160
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_22_clk
timestamp 1688980957
transform 1 0 21528 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_23_clk
timestamp 1688980957
transform -1 0 20240 0 -1 16864
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_24_clk
timestamp 1688980957
transform 1 0 13248 0 1 10336
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_25_clk
timestamp 1688980957
transform 1 0 13800 0 -1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_26_clk
timestamp 1688980957
transform 1 0 8648 0 1 7072
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_leaf_27_clk
timestamp 1688980957
transform -1 0 5336 0 1 5984
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32936 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout106
timestamp 1688980957
transform -1 0 14352 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout107
timestamp 1688980957
transform 1 0 15916 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout108
timestamp 1688980957
transform 1 0 15916 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout109
timestamp 1688980957
transform 1 0 14904 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout110 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout111 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout112 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16008 0 -1 17952
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout113
timestamp 1688980957
transform 1 0 20148 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout114
timestamp 1688980957
transform 1 0 20148 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout115
timestamp 1688980957
transform 1 0 19780 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout116
timestamp 1688980957
transform -1 0 16744 0 1 8160
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout117
timestamp 1688980957
transform 1 0 17020 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout118
timestamp 1688980957
transform -1 0 16652 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout119
timestamp 1688980957
transform -1 0 5612 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout120
timestamp 1688980957
transform -1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout121
timestamp 1688980957
transform 1 0 15732 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout122
timestamp 1688980957
transform 1 0 13156 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout123
timestamp 1688980957
transform -1 0 4508 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout124
timestamp 1688980957
transform -1 0 4784 0 -1 31008
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout125
timestamp 1688980957
transform 1 0 18400 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  fanout126
timestamp 1688980957
transform -1 0 6992 0 -1 33184
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout127
timestamp 1688980957
transform 1 0 18860 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout128
timestamp 1688980957
transform 1 0 20608 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout129
timestamp 1688980957
transform -1 0 27324 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout130
timestamp 1688980957
transform 1 0 27048 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout131
timestamp 1688980957
transform 1 0 20884 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  fanout132
timestamp 1688980957
transform 1 0 19504 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout133
timestamp 1688980957
transform 1 0 28336 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  fanout134
timestamp 1688980957
transform 1 0 19044 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  fanout135
timestamp 1688980957
transform 1 0 5428 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_76 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9752 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1688980957
transform 1 0 10948 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_93 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_113
timestamp 1688980957
transform 1 0 13156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1688980957
transform 1 0 13524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_121
timestamp 1688980957
transform 1 0 13892 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1688980957
transform 1 0 15732 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_149
timestamp 1688980957
transform 1 0 16468 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_169
timestamp 1688980957
transform 1 0 18308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_173
timestamp 1688980957
transform 1 0 18676 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_190
timestamp 1688980957
transform 1 0 20240 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1688980957
transform 1 0 20884 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_205
timestamp 1688980957
transform 1 0 21620 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_228
timestamp 1688980957
transform 1 0 23736 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_256
timestamp 1688980957
transform 1 0 26312 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_284
timestamp 1688980957
transform 1 0 28888 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_309
timestamp 1688980957
transform 1 0 31188 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_313
timestamp 1688980957
transform 1 0 31556 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_317
timestamp 1688980957
transform 1 0 31924 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_19
timestamp 1688980957
transform 1 0 4508 0 -1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_43 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 7820 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_57
timestamp 1688980957
transform 1 0 8004 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_65 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8740 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 10212 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 11316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 12420 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 12972 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_125
timestamp 1688980957
transform 1 0 14260 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_130
timestamp 1688980957
transform 1 0 14720 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_142
timestamp 1688980957
transform 1 0 15824 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_162
timestamp 1688980957
transform 1 0 17664 0 -1 3808
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 18308 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 19412 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_193
timestamp 1688980957
transform 1 0 20516 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_211
timestamp 1688980957
transform 1 0 22172 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 23276 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 23460 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 24564 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_249
timestamp 1688980957
transform 1 0 25668 0 -1 3808
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_254
timestamp 1688980957
transform 1 0 26128 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_266
timestamp 1688980957
transform 1 0 27232 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_278
timestamp 1688980957
transform 1 0 28336 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_281
timestamp 1688980957
transform 1 0 28612 0 -1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_285
timestamp 1688980957
transform 1 0 28980 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_297
timestamp 1688980957
transform 1 0 30084 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_309
timestamp 1688980957
transform 1 0 31188 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_317
timestamp 1688980957
transform 1 0 31924 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 5244 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_29
timestamp 1688980957
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_33
timestamp 1688980957
transform 1 0 5796 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_38
timestamp 1688980957
transform 1 0 6256 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_42
timestamp 1688980957
transform 1 0 6624 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_46
timestamp 1688980957
transform 1 0 6992 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_75
timestamp 1688980957
transform 1 0 9660 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 10396 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_109
timestamp 1688980957
transform 1 0 12788 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_115
timestamp 1688980957
transform 1 0 13340 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_128
timestamp 1688980957
transform 1 0 14536 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_132
timestamp 1688980957
transform 1 0 14904 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 1688980957
transform 1 0 15456 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_141
timestamp 1688980957
transform 1 0 15732 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_147
timestamp 1688980957
transform 1 0 16284 0 1 3808
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_151
timestamp 1688980957
transform 1 0 16652 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_163
timestamp 1688980957
transform 1 0 17756 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_167
timestamp 1688980957
transform 1 0 18124 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_179
timestamp 1688980957
transform 1 0 19228 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_190
timestamp 1688980957
transform 1 0 20240 0 1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_206
timestamp 1688980957
transform 1 0 21712 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_218
timestamp 1688980957
transform 1 0 22816 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_241
timestamp 1688980957
transform 1 0 24932 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1688980957
transform 1 0 25668 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_264
timestamp 1688980957
transform 1 0 27048 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_270
timestamp 1688980957
transform 1 0 27600 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_291
timestamp 1688980957
transform 1 0 29532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_303
timestamp 1688980957
transform 1 0 30636 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 31004 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 31188 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 32292 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_333
timestamp 1688980957
transform 1 0 33396 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_36
timestamp 1688980957
transform 1 0 6072 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_46
timestamp 1688980957
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_50
timestamp 1688980957
transform 1 0 7360 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_77
timestamp 1688980957
transform 1 0 9844 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_88
timestamp 1688980957
transform 1 0 10856 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_96
timestamp 1688980957
transform 1 0 11592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_101
timestamp 1688980957
transform 1 0 12052 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_105
timestamp 1688980957
transform 1 0 12420 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_109
timestamp 1688980957
transform 1 0 12788 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1688980957
transform 1 0 13156 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_143
timestamp 1688980957
transform 1 0 15916 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 18124 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_190
timestamp 1688980957
transform 1 0 20240 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 23276 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_273
timestamp 1688980957
transform 1 0 27876 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_277
timestamp 1688980957
transform 1 0 28244 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_293
timestamp 1688980957
transform 1 0 29716 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_317
timestamp 1688980957
transform 1 0 31924 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_337
timestamp 1688980957
transform 1 0 33764 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_49
timestamp 1688980957
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 1688980957
transform 1 0 11316 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_115
timestamp 1688980957
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_130
timestamp 1688980957
transform 1 0 14720 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1688980957
transform 1 0 15732 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_145
timestamp 1688980957
transform 1 0 16100 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_156
timestamp 1688980957
transform 1 0 17112 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_166
timestamp 1688980957
transform 1 0 18032 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_172
timestamp 1688980957
transform 1 0 18584 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_176
timestamp 1688980957
transform 1 0 18952 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_180
timestamp 1688980957
transform 1 0 19320 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_190
timestamp 1688980957
transform 1 0 20240 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 20608 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_197
timestamp 1688980957
transform 1 0 20884 0 1 4896
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_207
timestamp 1688980957
transform 1 0 21804 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_221
timestamp 1688980957
transform 1 0 23092 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_225
timestamp 1688980957
transform 1 0 23460 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_230
timestamp 1688980957
transform 1 0 23920 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_240
timestamp 1688980957
transform 1 0 24840 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_253
timestamp 1688980957
transform 1 0 26036 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_257
timestamp 1688980957
transform 1 0 26404 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_299
timestamp 1688980957
transform 1 0 30268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_303
timestamp 1688980957
transform 1 0 30636 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 31004 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_320
timestamp 1688980957
transform 1 0 32200 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_23
timestamp 1688980957
transform 1 0 4876 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_41
timestamp 1688980957
transform 1 0 6532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_65
timestamp 1688980957
transform 1 0 8740 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_161
timestamp 1688980957
transform 1 0 17572 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 18124 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_169
timestamp 1688980957
transform 1 0 18308 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_174
timestamp 1688980957
transform 1 0 18768 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_200
timestamp 1688980957
transform 1 0 21160 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_204
timestamp 1688980957
transform 1 0 21528 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_207
timestamp 1688980957
transform 1 0 21804 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_215
timestamp 1688980957
transform 1 0 22540 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_219
timestamp 1688980957
transform 1 0 22908 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 23276 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_225
timestamp 1688980957
transform 1 0 23460 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 28428 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_310
timestamp 1688980957
transform 1 0 31280 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_314
timestamp 1688980957
transform 1 0 31648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 33580 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_6
timestamp 1688980957
transform 1 0 3312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_29
timestamp 1688980957
transform 1 0 5428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_33
timestamp 1688980957
transform 1 0 5796 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_42
timestamp 1688980957
transform 1 0 6624 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_75
timestamp 1688980957
transform 1 0 9660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_79
timestamp 1688980957
transform 1 0 10028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_105
timestamp 1688980957
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_133
timestamp 1688980957
transform 1 0 14996 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_137
timestamp 1688980957
transform 1 0 15364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1688980957
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_152
timestamp 1688980957
transform 1 0 16744 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_191
timestamp 1688980957
transform 1 0 20332 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 20700 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_197
timestamp 1688980957
transform 1 0 20884 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_223
timestamp 1688980957
transform 1 0 23276 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_232
timestamp 1688980957
transform 1 0 24104 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_245
timestamp 1688980957
transform 1 0 25300 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 1688980957
transform 1 0 25668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_253
timestamp 1688980957
transform 1 0 26036 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_272
timestamp 1688980957
transform 1 0 27784 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_276
timestamp 1688980957
transform 1 0 28152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_294
timestamp 1688980957
transform 1 0 29808 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_298
timestamp 1688980957
transform 1 0 30176 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_302
timestamp 1688980957
transform 1 0 30544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 1688980957
transform 1 0 30912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_317
timestamp 1688980957
transform 1 0 31924 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_338
timestamp 1688980957
transform 1 0 33856 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_3
timestamp 1688980957
transform 1 0 3036 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_57
timestamp 1688980957
transform 1 0 8004 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_61
timestamp 1688980957
transform 1 0 8372 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_69
timestamp 1688980957
transform 1 0 9108 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_98
timestamp 1688980957
transform 1 0 11776 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_107
timestamp 1688980957
transform 1 0 12604 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_113
timestamp 1688980957
transform 1 0 13156 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_117
timestamp 1688980957
transform 1 0 13524 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_140
timestamp 1688980957
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_152
timestamp 1688980957
transform 1 0 16744 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_156
timestamp 1688980957
transform 1 0 17112 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_160
timestamp 1688980957
transform 1 0 17480 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 1688980957
transform 1 0 18308 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_173
timestamp 1688980957
transform 1 0 18676 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_212
timestamp 1688980957
transform 1 0 22264 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1688980957
transform 1 0 23184 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_250
timestamp 1688980957
transform 1 0 25760 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_254
timestamp 1688980957
transform 1 0 26128 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_277
timestamp 1688980957
transform 1 0 28244 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_310
timestamp 1688980957
transform 1 0 31280 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_314
timestamp 1688980957
transform 1 0 31648 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_337
timestamp 1688980957
transform 1 0 33764 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_19
timestamp 1688980957
transform 1 0 4508 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_44
timestamp 1688980957
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_48
timestamp 1688980957
transform 1 0 7176 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_52
timestamp 1688980957
transform 1 0 7544 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_60
timestamp 1688980957
transform 1 0 8280 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_96
timestamp 1688980957
transform 1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_130
timestamp 1688980957
transform 1 0 14720 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1688980957
transform 1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_153
timestamp 1688980957
transform 1 0 16836 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_175
timestamp 1688980957
transform 1 0 18860 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_181
timestamp 1688980957
transform 1 0 19412 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_212
timestamp 1688980957
transform 1 0 22264 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_235
timestamp 1688980957
transform 1 0 24380 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_248
timestamp 1688980957
transform 1 0 25576 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_273
timestamp 1688980957
transform 1 0 27876 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_286
timestamp 1688980957
transform 1 0 29072 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_335
timestamp 1688980957
transform 1 0 33580 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_339
timestamp 1688980957
transform 1 0 33948 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_6
timestamp 1688980957
transform 1 0 3312 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_28
timestamp 1688980957
transform 1 0 5336 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_48
timestamp 1688980957
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_52
timestamp 1688980957
transform 1 0 7544 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_57
timestamp 1688980957
transform 1 0 8004 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_71
timestamp 1688980957
transform 1 0 9292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_75
timestamp 1688980957
transform 1 0 9660 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_87
timestamp 1688980957
transform 1 0 10764 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_91
timestamp 1688980957
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_95
timestamp 1688980957
transform 1 0 11500 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_103
timestamp 1688980957
transform 1 0 12236 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_107
timestamp 1688980957
transform 1 0 12604 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_121
timestamp 1688980957
transform 1 0 13892 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_150
timestamp 1688980957
transform 1 0 16560 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_160
timestamp 1688980957
transform 1 0 17480 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_164
timestamp 1688980957
transform 1 0 17848 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_172
timestamp 1688980957
transform 1 0 18584 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_185
timestamp 1688980957
transform 1 0 19780 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_206
timestamp 1688980957
transform 1 0 21712 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_210
timestamp 1688980957
transform 1 0 22080 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_214
timestamp 1688980957
transform 1 0 22448 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_218
timestamp 1688980957
transform 1 0 22816 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1688980957
transform 1 0 23184 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_225
timestamp 1688980957
transform 1 0 23460 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_273
timestamp 1688980957
transform 1 0 27876 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_277
timestamp 1688980957
transform 1 0 28244 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_317
timestamp 1688980957
transform 1 0 31924 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 33580 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_337
timestamp 1688980957
transform 1 0 33764 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_23
timestamp 1688980957
transform 1 0 4876 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 5244 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_49
timestamp 1688980957
transform 1 0 7268 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_78
timestamp 1688980957
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 10304 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_85
timestamp 1688980957
transform 1 0 10580 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_89
timestamp 1688980957
transform 1 0 10948 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_93
timestamp 1688980957
transform 1 0 11316 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_97
timestamp 1688980957
transform 1 0 11684 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_105
timestamp 1688980957
transform 1 0 12420 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_133
timestamp 1688980957
transform 1 0 14996 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_166
timestamp 1688980957
transform 1 0 18032 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_172
timestamp 1688980957
transform 1 0 18584 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_184
timestamp 1688980957
transform 1 0 19688 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_191
timestamp 1688980957
transform 1 0 20332 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 20700 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_197
timestamp 1688980957
transform 1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_228
timestamp 1688980957
transform 1 0 23736 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_242
timestamp 1688980957
transform 1 0 25024 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_246
timestamp 1688980957
transform 1 0 25392 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 25760 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_253
timestamp 1688980957
transform 1 0 26036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_257
timestamp 1688980957
transform 1 0 26404 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_265
timestamp 1688980957
transform 1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_280
timestamp 1688980957
transform 1 0 28520 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_284
timestamp 1688980957
transform 1 0 28888 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_292
timestamp 1688980957
transform 1 0 29624 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_296
timestamp 1688980957
transform 1 0 29992 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_300
timestamp 1688980957
transform 1 0 30360 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_304
timestamp 1688980957
transform 1 0 30728 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_330
timestamp 1688980957
transform 1 0 33120 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_334
timestamp 1688980957
transform 1 0 33488 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_3
timestamp 1688980957
transform 1 0 3036 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_60
timestamp 1688980957
transform 1 0 8280 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_64
timestamp 1688980957
transform 1 0 8648 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_68
timestamp 1688980957
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_78
timestamp 1688980957
transform 1 0 9936 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_104
timestamp 1688980957
transform 1 0 12328 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_133
timestamp 1688980957
transform 1 0 14996 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_139
timestamp 1688980957
transform 1 0 15548 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_153
timestamp 1688980957
transform 1 0 16836 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_157
timestamp 1688980957
transform 1 0 17204 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_169
timestamp 1688980957
transform 1 0 18308 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_193
timestamp 1688980957
transform 1 0 20516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_233
timestamp 1688980957
transform 1 0 24196 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_248
timestamp 1688980957
transform 1 0 25576 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_270
timestamp 1688980957
transform 1 0 27600 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_315
timestamp 1688980957
transform 1 0 31740 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_326
timestamp 1688980957
transform 1 0 32752 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_334
timestamp 1688980957
transform 1 0 33488 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_337
timestamp 1688980957
transform 1 0 33764 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_19
timestamp 1688980957
transform 1 0 4508 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_37
timestamp 1688980957
transform 1 0 6164 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_64
timestamp 1688980957
transform 1 0 8648 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_68
timestamp 1688980957
transform 1 0 9016 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_76
timestamp 1688980957
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_80
timestamp 1688980957
transform 1 0 10120 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 10580 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_93
timestamp 1688980957
transform 1 0 11316 0 1 9248
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_98
timestamp 1688980957
transform 1 0 11776 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_110
timestamp 1688980957
transform 1 0 12880 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_116
timestamp 1688980957
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_126
timestamp 1688980957
transform 1 0 14352 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_130
timestamp 1688980957
transform 1 0 14720 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 15732 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_145
timestamp 1688980957
transform 1 0 16100 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_151
timestamp 1688980957
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_161
timestamp 1688980957
transform 1 0 17572 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_169
timestamp 1688980957
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_176
timestamp 1688980957
transform 1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_180
timestamp 1688980957
transform 1 0 19320 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_186
timestamp 1688980957
transform 1 0 19872 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_194
timestamp 1688980957
transform 1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_206
timestamp 1688980957
transform 1 0 21712 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_224
timestamp 1688980957
transform 1 0 23368 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_228
timestamp 1688980957
transform 1 0 23736 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_249
timestamp 1688980957
transform 1 0 25668 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_261
timestamp 1688980957
transform 1 0 26772 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_309
timestamp 1688980957
transform 1 0 31188 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_313
timestamp 1688980957
transform 1 0 31556 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_325
timestamp 1688980957
transform 1 0 32660 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_337
timestamp 1688980957
transform 1 0 33764 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 1688980957
transform 1 0 3036 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_46
timestamp 1688980957
transform 1 0 6992 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_50
timestamp 1688980957
transform 1 0 7360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1688980957
transform 1 0 7728 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_57
timestamp 1688980957
transform 1 0 8004 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_61
timestamp 1688980957
transform 1 0 8372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_65
timestamp 1688980957
transform 1 0 8740 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_69
timestamp 1688980957
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_73
timestamp 1688980957
transform 1 0 9476 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_79
timestamp 1688980957
transform 1 0 10028 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_87
timestamp 1688980957
transform 1 0 10764 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 13156 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_123
timestamp 1688980957
transform 1 0 14076 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_189
timestamp 1688980957
transform 1 0 20148 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 23276 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 1688980957
transform 1 0 23460 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_263
timestamp 1688980957
transform 1 0 26956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 27876 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 28428 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_321
timestamp 1688980957
transform 1 0 32292 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_333
timestamp 1688980957
transform 1 0 33396 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_23
timestamp 1688980957
transform 1 0 4876 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_68
timestamp 1688980957
transform 1 0 9016 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_80
timestamp 1688980957
transform 1 0 10120 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_85
timestamp 1688980957
transform 1 0 10580 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_134
timestamp 1688980957
transform 1 0 15088 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 15548 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_144
timestamp 1688980957
transform 1 0 16008 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_161
timestamp 1688980957
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_165
timestamp 1688980957
transform 1 0 17940 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_169
timestamp 1688980957
transform 1 0 18308 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_172
timestamp 1688980957
transform 1 0 18584 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_186
timestamp 1688980957
transform 1 0 19872 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_192
timestamp 1688980957
transform 1 0 20424 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_201
timestamp 1688980957
transform 1 0 21252 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_250
timestamp 1688980957
transform 1 0 25760 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_273
timestamp 1688980957
transform 1 0 27876 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_277
timestamp 1688980957
transform 1 0 28244 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_306
timestamp 1688980957
transform 1 0 30912 0 1 10336
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 31188 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_321
timestamp 1688980957
transform 1 0 32292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_31
timestamp 1688980957
transform 1 0 5612 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1688980957
transform 1 0 8740 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_86
timestamp 1688980957
transform 1 0 10672 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_94
timestamp 1688980957
transform 1 0 11408 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_108
timestamp 1688980957
transform 1 0 12696 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_125
timestamp 1688980957
transform 1 0 14260 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_136
timestamp 1688980957
transform 1 0 15272 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_140
timestamp 1688980957
transform 1 0 15640 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 18308 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_173
timestamp 1688980957
transform 1 0 18676 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_177
timestamp 1688980957
transform 1 0 19044 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_181
timestamp 1688980957
transform 1 0 19412 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_199
timestamp 1688980957
transform 1 0 21068 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_218
timestamp 1688980957
transform 1 0 22816 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_241
timestamp 1688980957
transform 1 0 24932 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_254
timestamp 1688980957
transform 1 0 26128 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1688980957
transform 1 0 28336 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_309
timestamp 1688980957
transform 1 0 31188 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_315
timestamp 1688980957
transform 1 0 31740 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_23
timestamp 1688980957
transform 1 0 4876 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_41
timestamp 1688980957
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_63
timestamp 1688980957
transform 1 0 8556 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_67
timestamp 1688980957
transform 1 0 8924 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_76
timestamp 1688980957
transform 1 0 9752 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1688980957
transform 1 0 10580 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_93
timestamp 1688980957
transform 1 0 11316 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_97
timestamp 1688980957
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_101
timestamp 1688980957
transform 1 0 12052 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_106
timestamp 1688980957
transform 1 0 12512 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_124
timestamp 1688980957
transform 1 0 14168 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_147
timestamp 1688980957
transform 1 0 16284 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_151
timestamp 1688980957
transform 1 0 16652 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_160
timestamp 1688980957
transform 1 0 17480 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_164
timestamp 1688980957
transform 1 0 17848 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_170
timestamp 1688980957
transform 1 0 18400 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_176
timestamp 1688980957
transform 1 0 18952 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_213
timestamp 1688980957
transform 1 0 22356 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_217
timestamp 1688980957
transform 1 0 22724 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_242
timestamp 1688980957
transform 1 0 25024 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_248
timestamp 1688980957
transform 1 0 25576 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_253
timestamp 1688980957
transform 1 0 26036 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_281
timestamp 1688980957
transform 1 0 28612 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_303
timestamp 1688980957
transform 1 0 30636 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 31004 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_312
timestamp 1688980957
transform 1 0 31464 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_316
timestamp 1688980957
transform 1 0 31832 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_337
timestamp 1688980957
transform 1 0 33764 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_3
timestamp 1688980957
transform 1 0 3036 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_53
timestamp 1688980957
transform 1 0 7636 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_60
timestamp 1688980957
transform 1 0 8280 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_101
timestamp 1688980957
transform 1 0 12052 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_105
timestamp 1688980957
transform 1 0 12420 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_122
timestamp 1688980957
transform 1 0 13984 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_128
timestamp 1688980957
transform 1 0 14536 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_156
timestamp 1688980957
transform 1 0 17112 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_183
timestamp 1688980957
transform 1 0 19596 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_187
timestamp 1688980957
transform 1 0 19964 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_192
timestamp 1688980957
transform 1 0 20424 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_222
timestamp 1688980957
transform 1 0 23184 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_232
timestamp 1688980957
transform 1 0 24104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_256
timestamp 1688980957
transform 1 0 26312 0 -1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_266
timestamp 1688980957
transform 1 0 27232 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_278
timestamp 1688980957
transform 1 0 28336 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_298
timestamp 1688980957
transform 1 0 30176 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_327
timestamp 1688980957
transform 1 0 32844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_331
timestamp 1688980957
transform 1 0 33212 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 33580 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_337
timestamp 1688980957
transform 1 0 33764 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_3
timestamp 1688980957
transform 1 0 3036 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_8
timestamp 1688980957
transform 1 0 3496 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_29
timestamp 1688980957
transform 1 0 5428 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_53
timestamp 1688980957
transform 1 0 7636 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_70
timestamp 1688980957
transform 1 0 9200 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_76
timestamp 1688980957
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_80
timestamp 1688980957
transform 1 0 10120 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1688980957
transform 1 0 10580 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_128
timestamp 1688980957
transform 1 0 14536 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 15548 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_169
timestamp 1688980957
transform 1 0 18308 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_173
timestamp 1688980957
transform 1 0 18676 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_189
timestamp 1688980957
transform 1 0 20148 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_193
timestamp 1688980957
transform 1 0 20516 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_197
timestamp 1688980957
transform 1 0 20884 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_201
timestamp 1688980957
transform 1 0 21252 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_261
timestamp 1688980957
transform 1 0 26772 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_276
timestamp 1688980957
transform 1 0 28152 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_288
timestamp 1688980957
transform 1 0 29256 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_299
timestamp 1688980957
transform 1 0 30268 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_317
timestamp 1688980957
transform 1 0 31924 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_329
timestamp 1688980957
transform 1 0 33028 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_19
timestamp 1688980957
transform 1 0 4508 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_40
timestamp 1688980957
transform 1 0 6440 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_52
timestamp 1688980957
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_62
timestamp 1688980957
transform 1 0 8464 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_66
timestamp 1688980957
transform 1 0 8832 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_72
timestamp 1688980957
transform 1 0 9384 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_76
timestamp 1688980957
transform 1 0 9752 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_86
timestamp 1688980957
transform 1 0 10672 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_90
timestamp 1688980957
transform 1 0 11040 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_93
timestamp 1688980957
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_105
timestamp 1688980957
transform 1 0 12420 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_109
timestamp 1688980957
transform 1 0 12788 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_121
timestamp 1688980957
transform 1 0 13892 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_148
timestamp 1688980957
transform 1 0 16376 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 18032 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_169
timestamp 1688980957
transform 1 0 18308 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_182
timestamp 1688980957
transform 1 0 19504 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_196
timestamp 1688980957
transform 1 0 20792 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_214
timestamp 1688980957
transform 1 0 22448 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_259
timestamp 1688980957
transform 1 0 26588 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 28428 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_288
timestamp 1688980957
transform 1 0 29256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_292
timestamp 1688980957
transform 1 0 29624 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_303
timestamp 1688980957
transform 1 0 30636 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_328
timestamp 1688980957
transform 1 0 32936 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_19
timestamp 1688980957
transform 1 0 4508 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1688980957
transform 1 0 5152 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_32
timestamp 1688980957
transform 1 0 5704 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_41
timestamp 1688980957
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_65
timestamp 1688980957
transform 1 0 8740 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1688980957
transform 1 0 10212 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1688980957
transform 1 0 10580 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp 1688980957
transform 1 0 10948 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_107
timestamp 1688980957
transform 1 0 12604 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_119
timestamp 1688980957
transform 1 0 13708 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_145
timestamp 1688980957
transform 1 0 16100 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_161
timestamp 1688980957
transform 1 0 17572 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_170
timestamp 1688980957
transform 1 0 18400 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_176
timestamp 1688980957
transform 1 0 18952 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_184
timestamp 1688980957
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_202
timestamp 1688980957
transform 1 0 21344 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_211
timestamp 1688980957
transform 1 0 22172 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_238
timestamp 1688980957
transform 1 0 24656 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_285
timestamp 1688980957
transform 1 0 28980 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_292
timestamp 1688980957
transform 1 0 29624 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 31004 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_314
timestamp 1688980957
transform 1 0 31648 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_320
timestamp 1688980957
transform 1 0 32200 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_329
timestamp 1688980957
transform 1 0 33028 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_339
timestamp 1688980957
transform 1 0 33948 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_45
timestamp 1688980957
transform 1 0 6900 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_49
timestamp 1688980957
transform 1 0 7268 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_52
timestamp 1688980957
transform 1 0 7544 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_80
timestamp 1688980957
transform 1 0 10120 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 12972 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_129
timestamp 1688980957
transform 1 0 14628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_134
timestamp 1688980957
transform 1 0 15088 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1688980957
transform 1 0 17940 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_169
timestamp 1688980957
transform 1 0 18308 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_220
timestamp 1688980957
transform 1 0 23000 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1688980957
transform 1 0 23460 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_229
timestamp 1688980957
transform 1 0 23828 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_233
timestamp 1688980957
transform 1 0 24196 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_237
timestamp 1688980957
transform 1 0 24564 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_241
timestamp 1688980957
transform 1 0 24932 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_247
timestamp 1688980957
transform 1 0 25484 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_261
timestamp 1688980957
transform 1 0 26772 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_281
timestamp 1688980957
transform 1 0 28612 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_314
timestamp 1688980957
transform 1 0 31648 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_331
timestamp 1688980957
transform 1 0 33212 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 33580 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_337
timestamp 1688980957
transform 1 0 33764 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_20
timestamp 1688980957
transform 1 0 4600 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_24
timestamp 1688980957
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1688980957
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_37
timestamp 1688980957
transform 1 0 6164 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_41
timestamp 1688980957
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_52
timestamp 1688980957
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_56
timestamp 1688980957
transform 1 0 7912 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_65
timestamp 1688980957
transform 1 0 8740 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_69
timestamp 1688980957
transform 1 0 9108 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_73
timestamp 1688980957
transform 1 0 9476 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_92
timestamp 1688980957
transform 1 0 11224 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_97
timestamp 1688980957
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_122
timestamp 1688980957
transform 1 0 13984 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_126
timestamp 1688980957
transform 1 0 14352 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_176
timestamp 1688980957
transform 1 0 18952 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 20608 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_224
timestamp 1688980957
transform 1 0 23368 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 25668 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_261
timestamp 1688980957
transform 1 0 26772 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_287
timestamp 1688980957
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_304
timestamp 1688980957
transform 1 0 30728 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_315
timestamp 1688980957
transform 1 0 31740 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_336
timestamp 1688980957
transform 1 0 33672 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_19
timestamp 1688980957
transform 1 0 4508 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_38
timestamp 1688980957
transform 1 0 6256 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 7728 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_62
timestamp 1688980957
transform 1 0 8464 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_82
timestamp 1688980957
transform 1 0 10304 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_88
timestamp 1688980957
transform 1 0 10856 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_93
timestamp 1688980957
transform 1 0 11316 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_97
timestamp 1688980957
transform 1 0 11684 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_102
timestamp 1688980957
transform 1 0 12144 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_106
timestamp 1688980957
transform 1 0 12512 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_116
timestamp 1688980957
transform 1 0 13432 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_144
timestamp 1688980957
transform 1 0 16008 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_162
timestamp 1688980957
transform 1 0 17664 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1688980957
transform 1 0 18308 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_195
timestamp 1688980957
transform 1 0 20700 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_205
timestamp 1688980957
transform 1 0 21620 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_215
timestamp 1688980957
transform 1 0 22540 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_219
timestamp 1688980957
transform 1 0 22908 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 23276 0 -1 15776
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_231
timestamp 1688980957
transform 1 0 24012 0 -1 15776
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_243
timestamp 1688980957
transform 1 0 25116 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_255
timestamp 1688980957
transform 1 0 26220 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_263
timestamp 1688980957
transform 1 0 26956 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_273
timestamp 1688980957
transform 1 0 27876 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1688980957
transform 1 0 28336 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_294
timestamp 1688980957
transform 1 0 29808 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1688980957
transform 1 0 5152 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_57
timestamp 1688980957
transform 1 0 8004 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_61
timestamp 1688980957
transform 1 0 8372 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_124
timestamp 1688980957
transform 1 0 14168 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_130
timestamp 1688980957
transform 1 0 14720 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1688980957
transform 1 0 15364 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_141
timestamp 1688980957
transform 1 0 15732 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_160
timestamp 1688980957
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_182
timestamp 1688980957
transform 1 0 19504 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_237
timestamp 1688980957
transform 1 0 24564 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_241
timestamp 1688980957
transform 1 0 24932 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1688980957
transform 1 0 25300 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 25852 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_287
timestamp 1688980957
transform 1 0 29164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_297
timestamp 1688980957
transform 1 0 30084 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1688980957
transform 1 0 30912 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_309
timestamp 1688980957
transform 1 0 31188 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_313
timestamp 1688980957
transform 1 0 31556 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_320
timestamp 1688980957
transform 1 0 32200 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_3
timestamp 1688980957
transform 1 0 3036 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_52
timestamp 1688980957
transform 1 0 7544 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_57
timestamp 1688980957
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_76
timestamp 1688980957
transform 1 0 9752 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_80
timestamp 1688980957
transform 1 0 10120 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1688980957
transform 1 0 12788 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_133
timestamp 1688980957
transform 1 0 14996 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_148
timestamp 1688980957
transform 1 0 16376 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_162
timestamp 1688980957
transform 1 0 17664 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_169
timestamp 1688980957
transform 1 0 18308 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_193
timestamp 1688980957
transform 1 0 20516 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_225
timestamp 1688980957
transform 1 0 23460 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_260
timestamp 1688980957
transform 1 0 26680 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_267
timestamp 1688980957
transform 1 0 27324 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_285
timestamp 1688980957
transform 1 0 28980 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_318
timestamp 1688980957
transform 1 0 32016 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_337
timestamp 1688980957
transform 1 0 33764 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1688980957
transform 1 0 5428 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_76
timestamp 1688980957
transform 1 0 9752 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_80
timestamp 1688980957
transform 1 0 10120 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_114
timestamp 1688980957
transform 1 0 13248 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_129
timestamp 1688980957
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_161
timestamp 1688980957
transform 1 0 17572 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_174
timestamp 1688980957
transform 1 0 18768 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_200
timestamp 1688980957
transform 1 0 21160 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_261
timestamp 1688980957
transform 1 0 26772 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_265
timestamp 1688980957
transform 1 0 27140 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_294
timestamp 1688980957
transform 1 0 29808 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_303
timestamp 1688980957
transform 1 0 30636 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 31004 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_337
timestamp 1688980957
transform 1 0 33764 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_23
timestamp 1688980957
transform 1 0 4876 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_48
timestamp 1688980957
transform 1 0 7176 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_52
timestamp 1688980957
transform 1 0 7544 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 7820 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_77
timestamp 1688980957
transform 1 0 9844 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 12972 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1688980957
transform 1 0 17940 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_177
timestamp 1688980957
transform 1 0 19044 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_200
timestamp 1688980957
transform 1 0 21160 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_222
timestamp 1688980957
transform 1 0 23184 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_245
timestamp 1688980957
transform 1 0 25300 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_251
timestamp 1688980957
transform 1 0 25852 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_272
timestamp 1688980957
transform 1 0 27784 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_292
timestamp 1688980957
transform 1 0 29624 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_296
timestamp 1688980957
transform 1 0 29992 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_3
timestamp 1688980957
transform 1 0 3036 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_21
timestamp 1688980957
transform 1 0 4692 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_25
timestamp 1688980957
transform 1 0 5060 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1688980957
transform 1 0 5428 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_51
timestamp 1688980957
transform 1 0 7452 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_57
timestamp 1688980957
transform 1 0 8004 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_77
timestamp 1688980957
transform 1 0 9844 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_85
timestamp 1688980957
transform 1 0 10580 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_96
timestamp 1688980957
transform 1 0 11592 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_118
timestamp 1688980957
transform 1 0 13616 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1688980957
transform 1 0 15364 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_149
timestamp 1688980957
transform 1 0 16468 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_179
timestamp 1688980957
transform 1 0 19228 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_184
timestamp 1688980957
transform 1 0 19688 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_188
timestamp 1688980957
transform 1 0 20056 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1688980957
transform 1 0 20608 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1688980957
transform 1 0 20884 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_298
timestamp 1688980957
transform 1 0 30176 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_306
timestamp 1688980957
transform 1 0 30912 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_338
timestamp 1688980957
transform 1 0 33856 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_6
timestamp 1688980957
transform 1 0 3312 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_47
timestamp 1688980957
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_51
timestamp 1688980957
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_57
timestamp 1688980957
transform 1 0 8004 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_76
timestamp 1688980957
transform 1 0 9752 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_80
timestamp 1688980957
transform 1 0 10120 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_84
timestamp 1688980957
transform 1 0 10488 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_108
timestamp 1688980957
transform 1 0 12696 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_122
timestamp 1688980957
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_145
timestamp 1688980957
transform 1 0 16100 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_189
timestamp 1688980957
transform 1 0 20148 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_193
timestamp 1688980957
transform 1 0 20516 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_197
timestamp 1688980957
transform 1 0 20884 0 -1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_203
timestamp 1688980957
transform 1 0 21436 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_215
timestamp 1688980957
transform 1 0 22540 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_221
timestamp 1688980957
transform 1 0 23092 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_233
timestamp 1688980957
transform 1 0 24196 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_254
timestamp 1688980957
transform 1 0 26128 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_276
timestamp 1688980957
transform 1 0 28152 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_313
timestamp 1688980957
transform 1 0 31556 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_337
timestamp 1688980957
transform 1 0 33764 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_19
timestamp 1688980957
transform 1 0 4508 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_32
timestamp 1688980957
transform 1 0 5704 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_71
timestamp 1688980957
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_75
timestamp 1688980957
transform 1 0 9660 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 10396 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_88
timestamp 1688980957
transform 1 0 10856 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_99
timestamp 1688980957
transform 1 0 11868 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_116
timestamp 1688980957
transform 1 0 13432 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_126
timestamp 1688980957
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 15548 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_144
timestamp 1688980957
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_148
timestamp 1688980957
transform 1 0 16376 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_152
timestamp 1688980957
transform 1 0 16744 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_200
timestamp 1688980957
transform 1 0 21160 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_208
timestamp 1688980957
transform 1 0 21896 0 1 19040
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_212
timestamp 1688980957
transform 1 0 22264 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_224
timestamp 1688980957
transform 1 0 23368 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_246
timestamp 1688980957
transform 1 0 25392 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_276
timestamp 1688980957
transform 1 0 28152 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_285
timestamp 1688980957
transform 1 0 28980 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_298
timestamp 1688980957
transform 1 0 30176 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_306
timestamp 1688980957
transform 1 0 30912 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_317
timestamp 1688980957
transform 1 0 31924 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_321
timestamp 1688980957
transform 1 0 32292 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_23
timestamp 1688980957
transform 1 0 4876 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_45
timestamp 1688980957
transform 1 0 6900 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 7820 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_65
timestamp 1688980957
transform 1 0 8740 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_84
timestamp 1688980957
transform 1 0 10488 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1688980957
transform 1 0 12604 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 13156 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_144
timestamp 1688980957
transform 1 0 16008 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_156
timestamp 1688980957
transform 1 0 17112 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_162
timestamp 1688980957
transform 1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_195
timestamp 1688980957
transform 1 0 20700 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_219
timestamp 1688980957
transform 1 0 22908 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_256
timestamp 1688980957
transform 1 0 26312 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_272
timestamp 1688980957
transform 1 0 27784 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_281
timestamp 1688980957
transform 1 0 28612 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_292
timestamp 1688980957
transform 1 0 29624 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_300
timestamp 1688980957
transform 1 0 30360 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_334
timestamp 1688980957
transform 1 0 33488 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_337
timestamp 1688980957
transform 1 0 33764 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1688980957
transform 1 0 3036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_7
timestamp 1688980957
transform 1 0 3404 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 5244 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_29
timestamp 1688980957
transform 1 0 5428 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_52
timestamp 1688980957
transform 1 0 7544 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_56
timestamp 1688980957
transform 1 0 7912 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_66
timestamp 1688980957
transform 1 0 8832 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_70
timestamp 1688980957
transform 1 0 9200 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_85
timestamp 1688980957
transform 1 0 10580 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_117
timestamp 1688980957
transform 1 0 13524 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_184
timestamp 1688980957
transform 1 0 19688 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 20700 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_200
timestamp 1688980957
transform 1 0 21160 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_210
timestamp 1688980957
transform 1 0 22080 0 1 20128
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_214
timestamp 1688980957
transform 1 0 22448 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_226
timestamp 1688980957
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_230
timestamp 1688980957
transform 1 0 23920 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_259
timestamp 1688980957
transform 1 0 26588 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_282
timestamp 1688980957
transform 1 0 28704 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_298
timestamp 1688980957
transform 1 0 30176 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_318
timestamp 1688980957
transform 1 0 32016 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_19
timestamp 1688980957
transform 1 0 4508 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_35
timestamp 1688980957
transform 1 0 5980 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_57
timestamp 1688980957
transform 1 0 8004 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_70
timestamp 1688980957
transform 1 0 9200 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_75
timestamp 1688980957
transform 1 0 9660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_86
timestamp 1688980957
transform 1 0 10672 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 12420 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 12972 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_113
timestamp 1688980957
transform 1 0 13156 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_134
timestamp 1688980957
transform 1 0 15088 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_146
timestamp 1688980957
transform 1 0 16192 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_155
timestamp 1688980957
transform 1 0 17020 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_161
timestamp 1688980957
transform 1 0 17572 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_164
timestamp 1688980957
transform 1 0 17848 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_201
timestamp 1688980957
transform 1 0 21252 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_210
timestamp 1688980957
transform 1 0 22080 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_214
timestamp 1688980957
transform 1 0 22448 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_218
timestamp 1688980957
transform 1 0 22816 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_225
timestamp 1688980957
transform 1 0 23460 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_232
timestamp 1688980957
transform 1 0 24104 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_236
timestamp 1688980957
transform 1 0 24472 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_259
timestamp 1688980957
transform 1 0 26588 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_277
timestamp 1688980957
transform 1 0 28244 0 -1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 28612 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_293
timestamp 1688980957
transform 1 0 29716 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_302
timestamp 1688980957
transform 1 0 30544 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_316
timestamp 1688980957
transform 1 0 31832 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1688980957
transform 1 0 33488 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_23
timestamp 1688980957
transform 1 0 4876 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_40
timestamp 1688980957
transform 1 0 6440 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_44
timestamp 1688980957
transform 1 0 6808 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_48
timestamp 1688980957
transform 1 0 7176 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_70
timestamp 1688980957
transform 1 0 9200 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_79
timestamp 1688980957
transform 1 0 10028 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 10396 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1688980957
transform 1 0 10580 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_91
timestamp 1688980957
transform 1 0 11132 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_99
timestamp 1688980957
transform 1 0 11868 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_123
timestamp 1688980957
transform 1 0 14076 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_135
timestamp 1688980957
transform 1 0 15180 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 15548 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_144
timestamp 1688980957
transform 1 0 16008 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_168
timestamp 1688980957
transform 1 0 18216 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_174
timestamp 1688980957
transform 1 0 18768 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_177
timestamp 1688980957
transform 1 0 19044 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_183
timestamp 1688980957
transform 1 0 19596 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_187
timestamp 1688980957
transform 1 0 19964 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 20700 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_197
timestamp 1688980957
transform 1 0 20884 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_218
timestamp 1688980957
transform 1 0 22816 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_222
timestamp 1688980957
transform 1 0 23184 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_246
timestamp 1688980957
transform 1 0 25392 0 1 21216
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_261
timestamp 1688980957
transform 1 0 26772 0 1 21216
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_273
timestamp 1688980957
transform 1 0 27876 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_285
timestamp 1688980957
transform 1 0 28980 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_289
timestamp 1688980957
transform 1 0 29348 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_317
timestamp 1688980957
transform 1 0 31924 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_323
timestamp 1688980957
transform 1 0 32476 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_3
timestamp 1688980957
transform 1 0 3036 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_39
timestamp 1688980957
transform 1 0 6348 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_43
timestamp 1688980957
transform 1 0 6716 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_47
timestamp 1688980957
transform 1 0 7084 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_63
timestamp 1688980957
transform 1 0 8556 0 -1 22304
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_83
timestamp 1688980957
transform 1 0 10396 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_106
timestamp 1688980957
transform 1 0 12512 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_124
timestamp 1688980957
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_147
timestamp 1688980957
transform 1 0 16284 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_159
timestamp 1688980957
transform 1 0 17388 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_176
timestamp 1688980957
transform 1 0 18952 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_182
timestamp 1688980957
transform 1 0 19504 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_207
timestamp 1688980957
transform 1 0 21804 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_211
timestamp 1688980957
transform 1 0 22172 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_215
timestamp 1688980957
transform 1 0 22540 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_245
timestamp 1688980957
transform 1 0 25300 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_249
timestamp 1688980957
transform 1 0 25668 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_257
timestamp 1688980957
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_268
timestamp 1688980957
transform 1 0 27416 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 28428 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_287
timestamp 1688980957
transform 1 0 29164 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_299
timestamp 1688980957
transform 1 0 30268 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_325
timestamp 1688980957
transform 1 0 32660 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1688980957
transform 1 0 33396 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_337
timestamp 1688980957
transform 1 0 33764 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1688980957
transform 1 0 5152 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_37
timestamp 1688980957
transform 1 0 6164 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_63
timestamp 1688980957
transform 1 0 8556 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_72
timestamp 1688980957
transform 1 0 9384 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_90
timestamp 1688980957
transform 1 0 11040 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_95
timestamp 1688980957
transform 1 0 11500 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_107
timestamp 1688980957
transform 1 0 12604 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_128
timestamp 1688980957
transform 1 0 14536 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_152
timestamp 1688980957
transform 1 0 16744 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_164
timestamp 1688980957
transform 1 0 17848 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_168
timestamp 1688980957
transform 1 0 18216 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_216
timestamp 1688980957
transform 1 0 22632 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_220
timestamp 1688980957
transform 1 0 23000 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 25852 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_253
timestamp 1688980957
transform 1 0 26036 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_272
timestamp 1688980957
transform 1 0 27784 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_281
timestamp 1688980957
transform 1 0 28612 0 1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_287
timestamp 1688980957
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_309
timestamp 1688980957
transform 1 0 31188 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_333
timestamp 1688980957
transform 1 0 33396 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_3
timestamp 1688980957
transform 1 0 3036 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 7820 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_74
timestamp 1688980957
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_81
timestamp 1688980957
transform 1 0 10212 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_91
timestamp 1688980957
transform 1 0 11132 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_95
timestamp 1688980957
transform 1 0 11500 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_109
timestamp 1688980957
transform 1 0 12788 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_121
timestamp 1688980957
transform 1 0 13892 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_152
timestamp 1688980957
transform 1 0 16744 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 1688980957
transform 1 0 17848 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_176
timestamp 1688980957
transform 1 0 18952 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_180
timestamp 1688980957
transform 1 0 19320 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_184
timestamp 1688980957
transform 1 0 19688 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_207
timestamp 1688980957
transform 1 0 21804 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_220
timestamp 1688980957
transform 1 0 23000 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_233
timestamp 1688980957
transform 1 0 24196 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_252
timestamp 1688980957
transform 1 0 25944 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_270
timestamp 1688980957
transform 1 0 27600 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 28428 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 1688980957
transform 1 0 28612 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_287
timestamp 1688980957
transform 1 0 29164 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_295
timestamp 1688980957
transform 1 0 29900 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_301
timestamp 1688980957
transform 1 0 30452 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_305
timestamp 1688980957
transform 1 0 30820 0 -1 23392
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 31924 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 33028 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 33580 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_337
timestamp 1688980957
transform 1 0 33764 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_19
timestamp 1688980957
transform 1 0 4508 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_29
timestamp 1688980957
transform 1 0 5428 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_39
timestamp 1688980957
transform 1 0 6348 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_48
timestamp 1688980957
transform 1 0 7176 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_71
timestamp 1688980957
transform 1 0 9292 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_80
timestamp 1688980957
transform 1 0 10120 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_85
timestamp 1688980957
transform 1 0 10580 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_90
timestamp 1688980957
transform 1 0 11040 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_105
timestamp 1688980957
transform 1 0 12420 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_111
timestamp 1688980957
transform 1 0 12972 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_117
timestamp 1688980957
transform 1 0 13524 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_149
timestamp 1688980957
transform 1 0 16468 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_159
timestamp 1688980957
transform 1 0 17388 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_167
timestamp 1688980957
transform 1 0 18124 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_171
timestamp 1688980957
transform 1 0 18492 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_178
timestamp 1688980957
transform 1 0 19136 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_190
timestamp 1688980957
transform 1 0 20240 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_197
timestamp 1688980957
transform 1 0 20884 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_201
timestamp 1688980957
transform 1 0 21252 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_207
timestamp 1688980957
transform 1 0 21804 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_228
timestamp 1688980957
transform 1 0 23736 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_261
timestamp 1688980957
transform 1 0 26772 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_265
timestamp 1688980957
transform 1 0 27140 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_269
timestamp 1688980957
transform 1 0 27508 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_281
timestamp 1688980957
transform 1 0 28612 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_289
timestamp 1688980957
transform 1 0 29348 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_300
timestamp 1688980957
transform 1 0 30360 0 1 23392
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 31188 0 1 23392
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 32292 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_333
timestamp 1688980957
transform 1 0 33396 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_339
timestamp 1688980957
transform 1 0 33948 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_3
timestamp 1688980957
transform 1 0 3036 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_11
timestamp 1688980957
transform 1 0 3772 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_49
timestamp 1688980957
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_77
timestamp 1688980957
transform 1 0 9844 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_81
timestamp 1688980957
transform 1 0 10212 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_100
timestamp 1688980957
transform 1 0 11960 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_104
timestamp 1688980957
transform 1 0 12328 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 12972 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_133
timestamp 1688980957
transform 1 0 14996 0 -1 24480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_139
timestamp 1688980957
transform 1 0 15548 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_151
timestamp 1688980957
transform 1 0 16652 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_157
timestamp 1688980957
transform 1 0 17204 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_169
timestamp 1688980957
transform 1 0 18308 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_173
timestamp 1688980957
transform 1 0 18676 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_177
timestamp 1688980957
transform 1 0 19044 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 19412 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_193
timestamp 1688980957
transform 1 0 20516 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_222
timestamp 1688980957
transform 1 0 23184 0 -1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_228
timestamp 1688980957
transform 1 0 23736 0 -1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_240
timestamp 1688980957
transform 1 0 24840 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_252
timestamp 1688980957
transform 1 0 25944 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_284
timestamp 1688980957
transform 1 0 28888 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_288
timestamp 1688980957
transform 1 0 29256 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_297
timestamp 1688980957
transform 1 0 30084 0 -1 24480
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_307
timestamp 1688980957
transform 1 0 31004 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_319
timestamp 1688980957
transform 1 0 32108 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_337
timestamp 1688980957
transform 1 0 33764 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_22
timestamp 1688980957
transform 1 0 4784 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_26
timestamp 1688980957
transform 1 0 5152 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_29
timestamp 1688980957
transform 1 0 5428 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_37
timestamp 1688980957
transform 1 0 6164 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_41
timestamp 1688980957
transform 1 0 6532 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_46
timestamp 1688980957
transform 1 0 6992 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_50
timestamp 1688980957
transform 1 0 7360 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_53
timestamp 1688980957
transform 1 0 7636 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_57
timestamp 1688980957
transform 1 0 8004 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_61
timestamp 1688980957
transform 1 0 8372 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_65
timestamp 1688980957
transform 1 0 8740 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_69
timestamp 1688980957
transform 1 0 9108 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_82
timestamp 1688980957
transform 1 0 10304 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_85
timestamp 1688980957
transform 1 0 10580 0 1 24480
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_99
timestamp 1688980957
transform 1 0 11868 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_111
timestamp 1688980957
transform 1 0 12972 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_123
timestamp 1688980957
transform 1 0 14076 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_135
timestamp 1688980957
transform 1 0 15180 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_162
timestamp 1688980957
transform 1 0 17664 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_178
timestamp 1688980957
transform 1 0 19136 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_182
timestamp 1688980957
transform 1 0 19504 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_194
timestamp 1688980957
transform 1 0 20608 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_206
timestamp 1688980957
transform 1 0 21712 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_216
timestamp 1688980957
transform 1 0 22632 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_220
timestamp 1688980957
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_224
timestamp 1688980957
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_237
timestamp 1688980957
transform 1 0 24564 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_248
timestamp 1688980957
transform 1 0 25576 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_274
timestamp 1688980957
transform 1 0 27968 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_305
timestamp 1688980957
transform 1 0 30820 0 1 24480
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 31188 0 1 24480
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 32292 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_333
timestamp 1688980957
transform 1 0 33396 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_339
timestamp 1688980957
transform 1 0 33948 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_31
timestamp 1688980957
transform 1 0 5612 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_51
timestamp 1688980957
transform 1 0 7452 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 7820 0 -1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_77
timestamp 1688980957
transform 1 0 9844 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_89
timestamp 1688980957
transform 1 0 10948 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_95
timestamp 1688980957
transform 1 0 11500 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_102
timestamp 1688980957
transform 1 0 12144 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1688980957
transform 1 0 12880 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 13156 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_143
timestamp 1688980957
transform 1 0 15916 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_147
timestamp 1688980957
transform 1 0 16284 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_169
timestamp 1688980957
transform 1 0 18308 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_216
timestamp 1688980957
transform 1 0 22632 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_253
timestamp 1688980957
transform 1 0 26036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_284
timestamp 1688980957
transform 1 0 28888 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_296
timestamp 1688980957
transform 1 0 29992 0 -1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_300
timestamp 1688980957
transform 1 0 30360 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_312
timestamp 1688980957
transform 1 0 31464 0 -1 25568
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_324
timestamp 1688980957
transform 1 0 32568 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_337
timestamp 1688980957
transform 1 0 33764 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_3
timestamp 1688980957
transform 1 0 3036 0 1 25568
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_14
timestamp 1688980957
transform 1 0 4048 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_26
timestamp 1688980957
transform 1 0 5152 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_29
timestamp 1688980957
transform 1 0 5428 0 1 25568
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_55
timestamp 1688980957
transform 1 0 7820 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_67
timestamp 1688980957
transform 1 0 8924 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_73
timestamp 1688980957
transform 1 0 9476 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 1688980957
transform 1 0 10212 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_90
timestamp 1688980957
transform 1 0 11040 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_96
timestamp 1688980957
transform 1 0 11592 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_171
timestamp 1688980957
transform 1 0 18492 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_180
timestamp 1688980957
transform 1 0 19320 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_184
timestamp 1688980957
transform 1 0 19688 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_200
timestamp 1688980957
transform 1 0 21160 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_230
timestamp 1688980957
transform 1 0 23920 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_260
timestamp 1688980957
transform 1 0 26680 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_265
timestamp 1688980957
transform 1 0 27140 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_269
timestamp 1688980957
transform 1 0 27508 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_290
timestamp 1688980957
transform 1 0 29440 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_294
timestamp 1688980957
transform 1 0 29808 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_302
timestamp 1688980957
transform 1 0 30544 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_309
timestamp 1688980957
transform 1 0 31188 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_317
timestamp 1688980957
transform 1 0 31924 0 1 25568
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_320
timestamp 1688980957
transform 1 0 32200 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_332
timestamp 1688980957
transform 1 0 33304 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 7820 0 -1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 8004 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_69
timestamp 1688980957
transform 1 0 9108 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_79
timestamp 1688980957
transform 1 0 10028 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_85
timestamp 1688980957
transform 1 0 10580 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_89
timestamp 1688980957
transform 1 0 10948 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_113
timestamp 1688980957
transform 1 0 13156 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_117
timestamp 1688980957
transform 1 0 13524 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_121
timestamp 1688980957
transform 1 0 13892 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_126
timestamp 1688980957
transform 1 0 14352 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_131
timestamp 1688980957
transform 1 0 14812 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_140
timestamp 1688980957
transform 1 0 15640 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_144
timestamp 1688980957
transform 1 0 16008 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_151
timestamp 1688980957
transform 1 0 16652 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_156
timestamp 1688980957
transform 1 0 17112 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_169
timestamp 1688980957
transform 1 0 18308 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_175
timestamp 1688980957
transform 1 0 18860 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_199
timestamp 1688980957
transform 1 0 21068 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_203
timestamp 1688980957
transform 1 0 21436 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_212
timestamp 1688980957
transform 1 0 22264 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_220
timestamp 1688980957
transform 1 0 23000 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_233
timestamp 1688980957
transform 1 0 24196 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_267
timestamp 1688980957
transform 1 0 27324 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_271
timestamp 1688980957
transform 1 0 27692 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_289
timestamp 1688980957
transform 1 0 29348 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_308
timestamp 1688980957
transform 1 0 31096 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_337
timestamp 1688980957
transform 1 0 33764 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_6
timestamp 1688980957
transform 1 0 3312 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_10
timestamp 1688980957
transform 1 0 3680 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_22
timestamp 1688980957
transform 1 0 4784 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_49
timestamp 1688980957
transform 1 0 7268 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_53
timestamp 1688980957
transform 1 0 7636 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_57
timestamp 1688980957
transform 1 0 8004 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 10396 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_93
timestamp 1688980957
transform 1 0 11316 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_116
timestamp 1688980957
transform 1 0 13432 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_123
timestamp 1688980957
transform 1 0 14076 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_141
timestamp 1688980957
transform 1 0 15732 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_162
timestamp 1688980957
transform 1 0 17664 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_170
timestamp 1688980957
transform 1 0 18400 0 1 26656
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_174
timestamp 1688980957
transform 1 0 18768 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_186
timestamp 1688980957
transform 1 0 19872 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_204
timestamp 1688980957
transform 1 0 21528 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_212
timestamp 1688980957
transform 1 0 22264 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_242
timestamp 1688980957
transform 1 0 25024 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 25852 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_276
timestamp 1688980957
transform 1 0 28152 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_280
timestamp 1688980957
transform 1 0 28520 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_284
timestamp 1688980957
transform 1 0 28888 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_332
timestamp 1688980957
transform 1 0 33304 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_336
timestamp 1688980957
transform 1 0 33672 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_34
timestamp 1688980957
transform 1 0 5888 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_50
timestamp 1688980957
transform 1 0 7360 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_54
timestamp 1688980957
transform 1 0 7728 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_57
timestamp 1688980957
transform 1 0 8004 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_63
timestamp 1688980957
transform 1 0 8556 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_71
timestamp 1688980957
transform 1 0 9292 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_76
timestamp 1688980957
transform 1 0 9752 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_84
timestamp 1688980957
transform 1 0 10488 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_91
timestamp 1688980957
transform 1 0 11132 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_107
timestamp 1688980957
transform 1 0 12604 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 12972 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_113
timestamp 1688980957
transform 1 0 13156 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_119
timestamp 1688980957
transform 1 0 13708 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_127
timestamp 1688980957
transform 1 0 14444 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_148
timestamp 1688980957
transform 1 0 16376 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_154
timestamp 1688980957
transform 1 0 16928 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_210
timestamp 1688980957
transform 1 0 22080 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_218
timestamp 1688980957
transform 1 0 22816 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_261
timestamp 1688980957
transform 1 0 26772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_265
timestamp 1688980957
transform 1 0 27140 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_274
timestamp 1688980957
transform 1 0 27968 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_278
timestamp 1688980957
transform 1 0 28336 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_299
timestamp 1688980957
transform 1 0 30268 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_321
timestamp 1688980957
transform 1 0 32292 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_334
timestamp 1688980957
transform 1 0 33488 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_3
timestamp 1688980957
transform 1 0 3036 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_11
timestamp 1688980957
transform 1 0 3772 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_29
timestamp 1688980957
transform 1 0 5428 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_71
timestamp 1688980957
transform 1 0 9292 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_75
timestamp 1688980957
transform 1 0 9660 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_79
timestamp 1688980957
transform 1 0 10028 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 10396 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_93
timestamp 1688980957
transform 1 0 11316 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_102
timestamp 1688980957
transform 1 0 12144 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_124
timestamp 1688980957
transform 1 0 14168 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_134
timestamp 1688980957
transform 1 0 15088 0 1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_161
timestamp 1688980957
transform 1 0 17572 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_165
timestamp 1688980957
transform 1 0 17940 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_173
timestamp 1688980957
transform 1 0 18676 0 1 27744
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_184
timestamp 1688980957
transform 1 0 19688 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_200
timestamp 1688980957
transform 1 0 21160 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_210
timestamp 1688980957
transform 1 0 22080 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_214
timestamp 1688980957
transform 1 0 22448 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_247
timestamp 1688980957
transform 1 0 25484 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 25852 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_263
timestamp 1688980957
transform 1 0 26956 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_306
timestamp 1688980957
transform 1 0 30912 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_318
timestamp 1688980957
transform 1 0 32016 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_19
timestamp 1688980957
transform 1 0 4508 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_57
timestamp 1688980957
transform 1 0 8004 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_90
timestamp 1688980957
transform 1 0 11040 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_102
timestamp 1688980957
transform 1 0 12144 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 1688980957
transform 1 0 12880 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_121
timestamp 1688980957
transform 1 0 13892 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_152
timestamp 1688980957
transform 1 0 16744 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_158
timestamp 1688980957
transform 1 0 17296 0 -1 28832
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_184
timestamp 1688980957
transform 1 0 19688 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_196
timestamp 1688980957
transform 1 0 20792 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 23184 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_275
timestamp 1688980957
transform 1 0 28060 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 28428 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_281
timestamp 1688980957
transform 1 0 28612 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_285
timestamp 1688980957
transform 1 0 28980 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 33580 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1688980957
transform 1 0 5152 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_38
timestamp 1688980957
transform 1 0 6256 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_42
timestamp 1688980957
transform 1 0 6624 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_48
timestamp 1688980957
transform 1 0 7176 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_69
timestamp 1688980957
transform 1 0 9108 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_76
timestamp 1688980957
transform 1 0 9752 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_93
timestamp 1688980957
transform 1 0 11316 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_104
timestamp 1688980957
transform 1 0 12328 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_115
timestamp 1688980957
transform 1 0 13340 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_126
timestamp 1688980957
transform 1 0 14352 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_135
timestamp 1688980957
transform 1 0 15180 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 15548 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_141
timestamp 1688980957
transform 1 0 15732 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_185
timestamp 1688980957
transform 1 0 19780 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_193
timestamp 1688980957
transform 1 0 20516 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_197
timestamp 1688980957
transform 1 0 20884 0 1 28832
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_240
timestamp 1688980957
transform 1 0 24840 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_253
timestamp 1688980957
transform 1 0 26036 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_267
timestamp 1688980957
transform 1 0 27324 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 31004 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_309
timestamp 1688980957
transform 1 0 31188 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_3
timestamp 1688980957
transform 1 0 3036 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_47
timestamp 1688980957
transform 1 0 7084 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 7820 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_57
timestamp 1688980957
transform 1 0 8004 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_68
timestamp 1688980957
transform 1 0 9016 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_87
timestamp 1688980957
transform 1 0 10764 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_95
timestamp 1688980957
transform 1 0 11500 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_128
timestamp 1688980957
transform 1 0 14536 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_132
timestamp 1688980957
transform 1 0 14904 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_136
timestamp 1688980957
transform 1 0 15272 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_140
timestamp 1688980957
transform 1 0 15640 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_150
timestamp 1688980957
transform 1 0 16560 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_158
timestamp 1688980957
transform 1 0 17296 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_162
timestamp 1688980957
transform 1 0 17664 0 -1 29920
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_177
timestamp 1688980957
transform 1 0 19044 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_189
timestamp 1688980957
transform 1 0 20148 0 -1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_201
timestamp 1688980957
transform 1 0 21252 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_213
timestamp 1688980957
transform 1 0 22356 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_221
timestamp 1688980957
transform 1 0 23092 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_225
timestamp 1688980957
transform 1 0 23460 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_229
timestamp 1688980957
transform 1 0 23828 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_233
timestamp 1688980957
transform 1 0 24196 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_246
timestamp 1688980957
transform 1 0 25392 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_250
timestamp 1688980957
transform 1 0 25760 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 28428 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_334
timestamp 1688980957
transform 1 0 33488 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_337
timestamp 1688980957
transform 1 0 33764 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_7
timestamp 1688980957
transform 1 0 3404 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_49
timestamp 1688980957
transform 1 0 7268 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_55
timestamp 1688980957
transform 1 0 7820 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_77
timestamp 1688980957
transform 1 0 9844 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_81
timestamp 1688980957
transform 1 0 10212 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_93
timestamp 1688980957
transform 1 0 11316 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_99
timestamp 1688980957
transform 1 0 11868 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_120
timestamp 1688980957
transform 1 0 13800 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_155
timestamp 1688980957
transform 1 0 17020 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_167
timestamp 1688980957
transform 1 0 18124 0 1 29920
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_179
timestamp 1688980957
transform 1 0 19228 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_191
timestamp 1688980957
transform 1 0 20332 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 20700 0 1 29920
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 20884 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_209
timestamp 1688980957
transform 1 0 21988 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_217
timestamp 1688980957
transform 1 0 22724 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_230
timestamp 1688980957
transform 1 0 23920 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_256
timestamp 1688980957
transform 1 0 26312 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_265
timestamp 1688980957
transform 1 0 27140 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_269
timestamp 1688980957
transform 1 0 27508 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_281
timestamp 1688980957
transform 1 0 28612 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_299
timestamp 1688980957
transform 1 0 30268 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_329
timestamp 1688980957
transform 1 0 33028 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_3
timestamp 1688980957
transform 1 0 3036 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_22
timestamp 1688980957
transform 1 0 4784 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_34
timestamp 1688980957
transform 1 0 5888 0 -1 31008
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_40
timestamp 1688980957
transform 1 0 6440 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_52
timestamp 1688980957
transform 1 0 7544 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_57
timestamp 1688980957
transform 1 0 8004 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_99
timestamp 1688980957
transform 1 0 11868 0 -1 31008
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_116
timestamp 1688980957
transform 1 0 13432 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_128
timestamp 1688980957
transform 1 0 14536 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_154
timestamp 1688980957
transform 1 0 16928 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 18124 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_172
timestamp 1688980957
transform 1 0 18584 0 -1 31008
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_186
timestamp 1688980957
transform 1 0 19872 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_198
timestamp 1688980957
transform 1 0 20976 0 -1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_210
timestamp 1688980957
transform 1 0 22080 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_222
timestamp 1688980957
transform 1 0 23184 0 -1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 25668 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_261
timestamp 1688980957
transform 1 0 26772 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_274
timestamp 1688980957
transform 1 0 27968 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_281
timestamp 1688980957
transform 1 0 28612 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 5152 0 1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 6532 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_53
timestamp 1688980957
transform 1 0 7636 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_74
timestamp 1688980957
transform 1 0 9568 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_85
timestamp 1688980957
transform 1 0 10580 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_94
timestamp 1688980957
transform 1 0 11408 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_98
timestamp 1688980957
transform 1 0 11776 0 1 31008
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_106
timestamp 1688980957
transform 1 0 12512 0 1 31008
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_118
timestamp 1688980957
transform 1 0 13616 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_130
timestamp 1688980957
transform 1 0 14720 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_134
timestamp 1688980957
transform 1 0 15088 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_141
timestamp 1688980957
transform 1 0 15732 0 1 31008
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_182
timestamp 1688980957
transform 1 0 19504 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 1688980957
transform 1 0 20608 0 1 31008
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 20884 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_209
timestamp 1688980957
transform 1 0 21988 0 1 31008
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_232
timestamp 1688980957
transform 1 0 24104 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_244
timestamp 1688980957
transform 1 0 25208 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_253
timestamp 1688980957
transform 1 0 26036 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_257
timestamp 1688980957
transform 1 0 26404 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_306
timestamp 1688980957
transform 1 0 30912 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_312
timestamp 1688980957
transform 1 0 31464 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_19
timestamp 1688980957
transform 1 0 4508 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_46
timestamp 1688980957
transform 1 0 6992 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_54
timestamp 1688980957
transform 1 0 7728 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_77
timestamp 1688980957
transform 1 0 9844 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_81
timestamp 1688980957
transform 1 0 10212 0 -1 32096
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_97
timestamp 1688980957
transform 1 0 11684 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_109
timestamp 1688980957
transform 1 0 12788 0 -1 32096
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 13156 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_125
timestamp 1688980957
transform 1 0 14260 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_133
timestamp 1688980957
transform 1 0 14996 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_165
timestamp 1688980957
transform 1 0 17940 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_178
timestamp 1688980957
transform 1 0 19136 0 -1 32096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_182
timestamp 1688980957
transform 1 0 19504 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_194
timestamp 1688980957
transform 1 0 20608 0 -1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_206
timestamp 1688980957
transform 1 0 21712 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_218
timestamp 1688980957
transform 1 0 22816 0 -1 32096
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_245
timestamp 1688980957
transform 1 0 25300 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_257
timestamp 1688980957
transform 1 0 26404 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_274
timestamp 1688980957
transform 1 0 27968 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_301
timestamp 1688980957
transform 1 0 30452 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_305
timestamp 1688980957
transform 1 0 30820 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_309
timestamp 1688980957
transform 1 0 31188 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_337
timestamp 1688980957
transform 1 0 33764 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_19
timestamp 1688980957
transform 1 0 4508 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_29
timestamp 1688980957
transform 1 0 5428 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_39
timestamp 1688980957
transform 1 0 6348 0 1 32096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_43
timestamp 1688980957
transform 1 0 6716 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_55
timestamp 1688980957
transform 1 0 7820 0 1 32096
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_72
timestamp 1688980957
transform 1 0 9384 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_90
timestamp 1688980957
transform 1 0 11040 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_98
timestamp 1688980957
transform 1 0 11776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_107
timestamp 1688980957
transform 1 0 12604 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_118
timestamp 1688980957
transform 1 0 13616 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_132
timestamp 1688980957
transform 1 0 14904 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_136
timestamp 1688980957
transform 1 0 15272 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_191
timestamp 1688980957
transform 1 0 20332 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 20700 0 1 32096
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 20884 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_209
timestamp 1688980957
transform 1 0 21988 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_217
timestamp 1688980957
transform 1 0 22724 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_242
timestamp 1688980957
transform 1 0 25024 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_250
timestamp 1688980957
transform 1 0 25760 0 1 32096
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 26036 0 1 32096
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 27140 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_288
timestamp 1688980957
transform 1 0 29256 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_300
timestamp 1688980957
transform 1 0 30360 0 1 32096
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 31188 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_321
timestamp 1688980957
transform 1 0 32292 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_46
timestamp 1688980957
transform 1 0 6992 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_50
timestamp 1688980957
transform 1 0 7360 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_57
timestamp 1688980957
transform 1 0 8004 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_65
timestamp 1688980957
transform 1 0 8740 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_84
timestamp 1688980957
transform 1 0 10488 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_88
timestamp 1688980957
transform 1 0 10856 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_95
timestamp 1688980957
transform 1 0 11500 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_119
timestamp 1688980957
transform 1 0 13708 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_143
timestamp 1688980957
transform 1 0 15916 0 -1 33184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_153
timestamp 1688980957
transform 1 0 16836 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_165
timestamp 1688980957
transform 1 0 17940 0 -1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_183
timestamp 1688980957
transform 1 0 19596 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_195
timestamp 1688980957
transform 1 0 20700 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_207
timestamp 1688980957
transform 1 0 21804 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_219
timestamp 1688980957
transform 1 0 22908 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 23276 0 -1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 23460 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 24564 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 25668 0 -1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 26772 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 27876 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 28428 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_281
timestamp 1688980957
transform 1 0 28612 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_287
timestamp 1688980957
transform 1 0 29164 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_337
timestamp 1688980957
transform 1 0 33764 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_3
timestamp 1688980957
transform 1 0 3036 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_22
timestamp 1688980957
transform 1 0 4784 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_26
timestamp 1688980957
transform 1 0 5152 0 1 33184
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_45
timestamp 1688980957
transform 1 0 6900 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_57
timestamp 1688980957
transform 1 0 8004 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_63
timestamp 1688980957
transform 1 0 8556 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_88
timestamp 1688980957
transform 1 0 10856 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_116
timestamp 1688980957
transform 1 0 13432 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 15732 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 16836 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_165
timestamp 1688980957
transform 1 0 17940 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_171
timestamp 1688980957
transform 1 0 18492 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_178
timestamp 1688980957
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_190
timestamp 1688980957
transform 1 0 20240 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_197
timestamp 1688980957
transform 1 0 20884 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_201
timestamp 1688980957
transform 1 0 21252 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_205
timestamp 1688980957
transform 1 0 21620 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_217
timestamp 1688980957
transform 1 0 22724 0 1 33184
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_229
timestamp 1688980957
transform 1 0 23828 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_241
timestamp 1688980957
transform 1 0 24932 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_249
timestamp 1688980957
transform 1 0 25668 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_253
timestamp 1688980957
transform 1 0 26036 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_257
timestamp 1688980957
transform 1 0 26404 0 1 33184
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_274
timestamp 1688980957
transform 1 0 27968 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_286
timestamp 1688980957
transform 1 0 29072 0 1 33184
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_325
timestamp 1688980957
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_337
timestamp 1688980957
transform 1 0 33764 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_6
timestamp 1688980957
transform 1 0 3312 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_29
timestamp 1688980957
transform 1 0 5428 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_33
timestamp 1688980957
transform 1 0 5796 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_50
timestamp 1688980957
transform 1 0 7360 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_60
timestamp 1688980957
transform 1 0 8280 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_95
timestamp 1688980957
transform 1 0 11500 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_107
timestamp 1688980957
transform 1 0 12604 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 12972 0 -1 34272
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_144
timestamp 1688980957
transform 1 0 16008 0 -1 34272
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_156
timestamp 1688980957
transform 1 0 17112 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_185
timestamp 1688980957
transform 1 0 19780 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_193
timestamp 1688980957
transform 1 0 20516 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_213
timestamp 1688980957
transform 1 0 22356 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_219
timestamp 1688980957
transform 1 0 22908 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 23276 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_225
timestamp 1688980957
transform 1 0 23460 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_229
timestamp 1688980957
transform 1 0 23828 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_246
timestamp 1688980957
transform 1 0 25392 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_269
timestamp 1688980957
transform 1 0 27508 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_277
timestamp 1688980957
transform 1 0 28244 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_297
timestamp 1688980957
transform 1 0 30084 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_305
timestamp 1688980957
transform 1 0 30820 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_325
timestamp 1688980957
transform 1 0 32660 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_333
timestamp 1688980957
transform 1 0 33396 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_337
timestamp 1688980957
transform 1 0 33764 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24196 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 9752 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 9844 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 9016 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform 1 0 9568 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 25852 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform -1 0 26036 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 23736 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 24472 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform 1 0 21068 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 23000 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 30636 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform 1 0 29164 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 31096 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform 1 0 29900 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 14904 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform -1 0 16468 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 6256 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 5428 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform -1 0 25116 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 24932 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 6992 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 8740 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 12236 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 11592 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 7820 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform 1 0 5152 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 6256 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 7084 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold30
timestamp 1688980957
transform -1 0 10304 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 9292 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 28060 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform -1 0 29900 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 7176 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform 1 0 3864 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform -1 0 33580 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 33580 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform -1 0 11408 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform 1 0 9108 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform 1 0 13800 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 15272 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform -1 0 31924 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 31924 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform -1 0 26772 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 25668 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform 1 0 29532 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 32016 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 26772 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 25944 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform -1 0 31096 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 30268 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform -1 0 19872 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 19044 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold54
timestamp 1688980957
transform -1 0 9660 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform 1 0 9752 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10488 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 9476 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 20792 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform 1 0 19872 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 25852 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform 1 0 22632 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 26772 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 25852 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform -1 0 14720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 14444 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform -1 0 11316 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform 1 0 8924 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 30452 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 33580 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 31924 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 31188 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold72 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11868 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 3404 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform -1 0 6624 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 5336 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform -1 0 5612 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform -1 0 3864 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 23920 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 22264 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold80
timestamp 1688980957
transform 1 0 17940 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  hold81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14444 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 8004 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform 1 0 6348 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold84
timestamp 1688980957
transform 1 0 17756 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 23552 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold86
timestamp 1688980957
transform 1 0 20884 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 29808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 6164 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 6532 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 7636 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold91
timestamp 1688980957
transform 1 0 7820 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform 1 0 4508 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 5336 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold94
timestamp 1688980957
transform 1 0 16284 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform -1 0 5336 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold96
timestamp 1688980957
transform 1 0 4600 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform 1 0 5704 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 13340 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform 1 0 13984 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 5612 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 3772 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 5796 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform 1 0 4508 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform -1 0 26404 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold105
timestamp 1688980957
transform -1 0 25024 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold106
timestamp 1688980957
transform -1 0 23276 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 20792 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold108
timestamp 1688980957
transform 1 0 23460 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 22540 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 25760 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold111
timestamp 1688980957
transform -1 0 26496 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform 1 0 21160 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform -1 0 22632 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold114
timestamp 1688980957
transform -1 0 10672 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  hold115
timestamp 1688980957
transform 1 0 8924 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform -1 0 8740 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold117
timestamp 1688980957
transform 1 0 17664 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform 1 0 19780 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold119
timestamp 1688980957
transform -1 0 20240 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform 1 0 28888 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold121
timestamp 1688980957
transform -1 0 11868 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform 1 0 6716 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 7084 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform 1 0 23460 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 21988 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform 1 0 23092 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform -1 0 22264 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold128
timestamp 1688980957
transform 1 0 10948 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  hold129
timestamp 1688980957
transform 1 0 19412 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform -1 0 29348 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 29992 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform 1 0 29992 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform -1 0 24196 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 23184 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform -1 0 24932 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 25668 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform 1 0 11040 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform -1 0 11316 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform 1 0 8188 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform -1 0 8740 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 22264 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 21528 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold143
timestamp 1688980957
transform 1 0 6808 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 6808 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 23460 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform -1 0 5336 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform 1 0 5336 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 6900 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform 1 0 4600 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform -1 0 6900 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform 1 0 3496 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 22264 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 28428 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform -1 0 27324 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform 1 0 27692 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform 1 0 27048 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform -1 0 29440 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform -1 0 28612 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform -1 0 33948 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform -1 0 33028 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold162
timestamp 1688980957
transform 1 0 14168 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform 1 0 28336 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold164
timestamp 1688980957
transform -1 0 15088 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold165 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15548 0 1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform -1 0 30176 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform -1 0 27692 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform 1 0 13432 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform -1 0 13064 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform -1 0 24840 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform 1 0 24196 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold173
timestamp 1688980957
transform 1 0 19596 0 1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform -1 0 19044 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform 1 0 23460 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform -1 0 24748 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold177
timestamp 1688980957
transform -1 0 20056 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  hold178
timestamp 1688980957
transform 1 0 19412 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 12236 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform 1 0 24288 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 6992 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform 1 0 5152 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform 1 0 6072 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform -1 0 31556 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform -1 0 30912 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 29992 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 29256 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform -1 0 5336 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform -1 0 4324 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold190
timestamp 1688980957
transform 1 0 11132 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 13156 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform 1 0 11132 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 24932 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform -1 0 24196 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform -1 0 31004 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 30636 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold197
timestamp 1688980957
transform 1 0 9016 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform 1 0 11684 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform -1 0 13892 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform -1 0 23184 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform -1 0 22264 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform 1 0 5428 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform 1 0 3864 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform -1 0 24564 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform 1 0 24748 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform -1 0 32660 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform 1 0 30360 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform 1 0 14352 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform -1 0 15640 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold210
timestamp 1688980957
transform 1 0 13616 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform 1 0 13616 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform -1 0 18216 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform -1 0 17940 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform 1 0 26404 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform 1 0 27048 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform 1 0 27140 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform -1 0 32752 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform -1 0 27876 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 26772 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold220
timestamp 1688980957
transform -1 0 13892 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold221
timestamp 1688980957
transform -1 0 30360 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform 1 0 27048 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold223
timestamp 1688980957
transform -1 0 14536 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform -1 0 15916 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform 1 0 5980 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold226
timestamp 1688980957
transform -1 0 5336 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold227
timestamp 1688980957
transform -1 0 31924 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold228
timestamp 1688980957
transform 1 0 30176 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform -1 0 19044 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold230
timestamp 1688980957
transform -1 0 12604 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 29900 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold232
timestamp 1688980957
transform 1 0 27416 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform -1 0 33764 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform -1 0 7176 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform 1 0 6624 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold236
timestamp 1688980957
transform -1 0 8740 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 18032 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform 1 0 12236 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform 1 0 27968 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold240
timestamp 1688980957
transform -1 0 33488 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 30360 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform -1 0 17480 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform -1 0 16744 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold244
timestamp 1688980957
transform 1 0 13432 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold245
timestamp 1688980957
transform -1 0 15548 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold246
timestamp 1688980957
transform -1 0 15364 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold247
timestamp 1688980957
transform 1 0 12328 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold248
timestamp 1688980957
transform 1 0 11592 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold249
timestamp 1688980957
transform 1 0 17572 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold250
timestamp 1688980957
transform -1 0 8648 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold251
timestamp 1688980957
transform -1 0 7084 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold252
timestamp 1688980957
transform 1 0 11684 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold253
timestamp 1688980957
transform 1 0 26496 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold254
timestamp 1688980957
transform -1 0 32200 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold255
timestamp 1688980957
transform 1 0 18308 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold256
timestamp 1688980957
transform 1 0 22356 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold257
timestamp 1688980957
transform 1 0 20976 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold258
timestamp 1688980957
transform 1 0 14996 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold259
timestamp 1688980957
transform -1 0 15272 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold260
timestamp 1688980957
transform -1 0 9108 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  hold261 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold262
timestamp 1688980957
transform 1 0 8832 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold263
timestamp 1688980957
transform 1 0 27876 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold264
timestamp 1688980957
transform -1 0 32568 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold265
timestamp 1688980957
transform -1 0 11868 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold266
timestamp 1688980957
transform -1 0 5612 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold267
timestamp 1688980957
transform -1 0 15640 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold268
timestamp 1688980957
transform -1 0 14904 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold269
timestamp 1688980957
transform -1 0 20976 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold270
timestamp 1688980957
transform 1 0 28612 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold271
timestamp 1688980957
transform -1 0 28980 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold272
timestamp 1688980957
transform -1 0 22540 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold273
timestamp 1688980957
transform -1 0 21620 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold274
timestamp 1688980957
transform 1 0 29532 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold275
timestamp 1688980957
transform -1 0 29348 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold276
timestamp 1688980957
transform -1 0 18400 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold277
timestamp 1688980957
transform -1 0 16468 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold278
timestamp 1688980957
transform -1 0 30360 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold279
timestamp 1688980957
transform 1 0 27784 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold280
timestamp 1688980957
transform -1 0 26772 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold281
timestamp 1688980957
transform -1 0 16560 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold282
timestamp 1688980957
transform -1 0 15640 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold283
timestamp 1688980957
transform 1 0 16376 0 -1 14688
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold284
timestamp 1688980957
transform 1 0 26864 0 1 22304
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold285
timestamp 1688980957
transform -1 0 25944 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold286
timestamp 1688980957
transform 1 0 22264 0 -1 12512
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold287
timestamp 1688980957
transform -1 0 32844 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold288
timestamp 1688980957
transform -1 0 19688 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold289
timestamp 1688980957
transform -1 0 17664 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold290
timestamp 1688980957
transform -1 0 17020 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold291
timestamp 1688980957
transform 1 0 28888 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold292
timestamp 1688980957
transform 1 0 29532 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold293
timestamp 1688980957
transform 1 0 30360 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold294
timestamp 1688980957
transform 1 0 10672 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold295
timestamp 1688980957
transform -1 0 13892 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold296
timestamp 1688980957
transform 1 0 26496 0 -1 19040
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold297
timestamp 1688980957
transform -1 0 26772 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold298
timestamp 1688980957
transform -1 0 13064 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold299
timestamp 1688980957
transform 1 0 12604 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold300
timestamp 1688980957
transform 1 0 11224 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold301
timestamp 1688980957
transform -1 0 11224 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold302
timestamp 1688980957
transform -1 0 9752 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold303
timestamp 1688980957
transform 1 0 9476 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold304
timestamp 1688980957
transform -1 0 9200 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold305
timestamp 1688980957
transform -1 0 20240 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold306
timestamp 1688980957
transform -1 0 17296 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold307
timestamp 1688980957
transform -1 0 10948 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold308
timestamp 1688980957
transform -1 0 10028 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold309
timestamp 1688980957
transform -1 0 31188 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold310
timestamp 1688980957
transform -1 0 30268 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold311
timestamp 1688980957
transform 1 0 28244 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold312
timestamp 1688980957
transform -1 0 29348 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold313
timestamp 1688980957
transform 1 0 28888 0 -1 15776
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold314
timestamp 1688980957
transform 1 0 31188 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold315
timestamp 1688980957
transform 1 0 11132 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold316
timestamp 1688980957
transform -1 0 10488 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  hold317
timestamp 1688980957
transform -1 0 29256 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold318
timestamp 1688980957
transform -1 0 28152 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold319
timestamp 1688980957
transform -1 0 31004 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold320
timestamp 1688980957
transform -1 0 29992 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold321
timestamp 1688980957
transform -1 0 27508 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold322
timestamp 1688980957
transform -1 0 26772 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold323
timestamp 1688980957
transform 1 0 13616 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold324
timestamp 1688980957
transform -1 0 12696 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold325
timestamp 1688980957
transform 1 0 18952 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold326
timestamp 1688980957
transform -1 0 5336 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold327
timestamp 1688980957
transform -1 0 10488 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold328
timestamp 1688980957
transform 1 0 9752 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold329
timestamp 1688980957
transform -1 0 9936 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold330
timestamp 1688980957
transform -1 0 16376 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold331
timestamp 1688980957
transform 1 0 26036 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold332
timestamp 1688980957
transform -1 0 25944 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold333
timestamp 1688980957
transform -1 0 9936 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold334
timestamp 1688980957
transform -1 0 15640 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold335
timestamp 1688980957
transform 1 0 16100 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold336
timestamp 1688980957
transform 1 0 13156 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold337
timestamp 1688980957
transform 1 0 30360 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold338
timestamp 1688980957
transform -1 0 31740 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold339
timestamp 1688980957
transform 1 0 30360 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold340
timestamp 1688980957
transform -1 0 32752 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold341
timestamp 1688980957
transform -1 0 31832 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold342
timestamp 1688980957
transform -1 0 26036 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold343
timestamp 1688980957
transform 1 0 24380 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold344
timestamp 1688980957
transform -1 0 14720 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold345
timestamp 1688980957
transform -1 0 13432 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold346
timestamp 1688980957
transform 1 0 16836 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold347
timestamp 1688980957
transform -1 0 15364 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold348
timestamp 1688980957
transform 1 0 11408 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold349
timestamp 1688980957
transform -1 0 13892 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold350
timestamp 1688980957
transform 1 0 27784 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold351
timestamp 1688980957
transform -1 0 27784 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold352
timestamp 1688980957
transform -1 0 26588 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold353
timestamp 1688980957
transform -1 0 26772 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold354
timestamp 1688980957
transform -1 0 25392 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold355
timestamp 1688980957
transform -1 0 11316 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold356
timestamp 1688980957
transform -1 0 31924 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold357
timestamp 1688980957
transform -1 0 31556 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold358
timestamp 1688980957
transform 1 0 31096 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold359
timestamp 1688980957
transform 1 0 28612 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold360
timestamp 1688980957
transform -1 0 31096 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold361
timestamp 1688980957
transform -1 0 16100 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold362
timestamp 1688980957
transform -1 0 31924 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold363
timestamp 1688980957
transform -1 0 18584 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold364
timestamp 1688980957
transform -1 0 28520 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold365
timestamp 1688980957
transform -1 0 30360 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold366
timestamp 1688980957
transform -1 0 25760 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold367
timestamp 1688980957
transform 1 0 7084 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold368
timestamp 1688980957
transform -1 0 26772 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold369
timestamp 1688980957
transform -1 0 25208 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold370
timestamp 1688980957
transform -1 0 16468 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold371
timestamp 1688980957
transform -1 0 17020 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold372
timestamp 1688980957
transform -1 0 16468 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold373
timestamp 1688980957
transform -1 0 13892 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold374
timestamp 1688980957
transform 1 0 5980 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold375
timestamp 1688980957
transform 1 0 8280 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold376
timestamp 1688980957
transform -1 0 15640 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold377
timestamp 1688980957
transform -1 0 15640 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold378
timestamp 1688980957
transform 1 0 17112 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold379
timestamp 1688980957
transform 1 0 16928 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold380
timestamp 1688980957
transform 1 0 10212 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold381
timestamp 1688980957
transform -1 0 19044 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold382
timestamp 1688980957
transform -1 0 11316 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold383
timestamp 1688980957
transform 1 0 24288 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold384
timestamp 1688980957
transform 1 0 8924 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold385
timestamp 1688980957
transform 1 0 25300 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold386
timestamp 1688980957
transform -1 0 20700 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold387
timestamp 1688980957
transform 1 0 17112 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold388
timestamp 1688980957
transform 1 0 11868 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold389
timestamp 1688980957
transform 1 0 20332 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold390
timestamp 1688980957
transform -1 0 16100 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1688980957
transform 1 0 3036 0 1 24480
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform 1 0 3036 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 34040 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform -1 0 15640 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform -1 0 34040 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 9476 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1688980957
transform -1 0 34040 0 1 29920
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform -1 0 34040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 21344 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 3312 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1688980957
transform 1 0 10580 0 -1 34272
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 16008 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1688980957
transform -1 0 32200 0 -1 32096
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform -1 0 34040 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 18860 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 13616 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 34040 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform -1 0 34040 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform -1 0 3312 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 22632 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 8004 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 28612 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 3036 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform -1 0 23736 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1688980957
transform 1 0 5428 0 1 2720
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 11040 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform -1 0 34040 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 3036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform -1 0 34040 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 26036 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1688980957
transform 1 0 3036 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform -1 0 33764 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 3036 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 33764 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output37 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22356 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 1688980957
transform -1 0 4508 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output39
timestamp 1688980957
transform 1 0 23920 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output40
timestamp 1688980957
transform -1 0 4508 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output41
timestamp 1688980957
transform -1 0 4508 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output42
timestamp 1688980957
transform 1 0 32568 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output43
timestamp 1688980957
transform -1 0 4508 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output44
timestamp 1688980957
transform -1 0 4508 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output45
timestamp 1688980957
transform 1 0 32200 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output46
timestamp 1688980957
transform -1 0 4508 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output47
timestamp 1688980957
transform -1 0 33672 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output48
timestamp 1688980957
transform -1 0 4508 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output49
timestamp 1688980957
transform -1 0 4508 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output50
timestamp 1688980957
transform 1 0 32200 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output51
timestamp 1688980957
transform 1 0 32200 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output52
timestamp 1688980957
transform 1 0 32568 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output53
timestamp 1688980957
transform 1 0 32568 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output54
timestamp 1688980957
transform 1 0 32568 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output55
timestamp 1688980957
transform -1 0 5336 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output56
timestamp 1688980957
transform 1 0 3036 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output57
timestamp 1688980957
transform 1 0 26496 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output58
timestamp 1688980957
transform 1 0 14168 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output59
timestamp 1688980957
transform -1 0 32200 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output60
timestamp 1688980957
transform -1 0 31096 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output61
timestamp 1688980957
transform 1 0 8004 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output62
timestamp 1688980957
transform -1 0 5336 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output63
timestamp 1688980957
transform 1 0 3036 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1688980957
transform 1 0 32568 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1688980957
transform 1 0 31188 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1688980957
transform 1 0 32200 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1688980957
transform 1 0 27048 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1688980957
transform 1 0 32568 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1688980957
transform 1 0 32568 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1688980957
transform 1 0 13156 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1688980957
transform 1 0 32200 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1688980957
transform 1 0 29624 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1688980957
transform 1 0 32200 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1688980957
transform 1 0 16744 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1688980957
transform -1 0 4508 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1688980957
transform -1 0 4508 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1688980957
transform -1 0 4508 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1688980957
transform 1 0 21896 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1688980957
transform 1 0 5888 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1688980957
transform 1 0 18308 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1688980957
transform -1 0 4508 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1688980957
transform -1 0 5980 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1688980957
transform -1 0 6716 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1688980957
transform -1 0 4508 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1688980957
transform 1 0 32200 0 -1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1688980957
transform 1 0 26036 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1688980957
transform 1 0 16192 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1688980957
transform 1 0 29256 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1688980957
transform 1 0 32200 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1688980957
transform 1 0 5428 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1688980957
transform -1 0 4508 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1688980957
transform -1 0 7912 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1688980957
transform -1 0 13064 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1688980957
transform 1 0 18768 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1688980957
transform 1 0 32568 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1688980957
transform 1 0 20700 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1688980957
transform 1 0 31188 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1688980957
transform -1 0 30084 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1688980957
transform -1 0 4784 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1688980957
transform 1 0 9016 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1688980957
transform 1 0 24472 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1688980957
transform -1 0 4508 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1688980957
transform -1 0 4508 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1688980957
transform 1 0 32200 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 2760 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 34316 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 2760 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 34316 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 2760 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 34316 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 2760 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 34316 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 2760 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 34316 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 2760 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 34316 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 2760 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 34316 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 2760 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 34316 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 2760 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 34316 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 2760 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 34316 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 2760 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 34316 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 2760 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 34316 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 2760 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 34316 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 2760 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 34316 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 2760 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 34316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 2760 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 34316 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 2760 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 34316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 2760 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 34316 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 2760 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 34316 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 2760 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 34316 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 2760 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 34316 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 2760 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 34316 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 2760 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 34316 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 2760 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 34316 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 2760 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 34316 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 2760 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 34316 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 2760 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 34316 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 2760 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 34316 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 2760 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 34316 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 2760 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 34316 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 2760 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 34316 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 2760 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 34316 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 2760 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 34316 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 2760 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 34316 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 2760 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 34316 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 2760 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 34316 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 2760 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 34316 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 2760 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 34316 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 2760 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 34316 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 2760 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 34316 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 2760 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 34316 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 2760 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 34316 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 2760 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 34316 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 2760 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 34316 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 2760 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 34316 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 2760 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 34316 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 2760 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 34316 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 2760 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 34316 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 2760 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 34316 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 2760 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 34316 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 2760 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 34316 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 2760 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 34316 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 2760 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 34316 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 2760 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 34316 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 2760 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 34316 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 2760 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 34316 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 2760 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 34316 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 2760 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 34316 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 7912 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 10488 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 13064 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 15640 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 18216 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 20792 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 23368 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 25944 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 28520 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 31096 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 33672 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 7912 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 13064 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 18216 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 23368 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 28520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 33672 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 5336 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 10488 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 15640 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 20792 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 25944 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 31096 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 7912 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 13064 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 18216 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 23368 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 28520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 33672 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 5336 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 10488 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 15640 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 20792 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 25944 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 31096 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 7912 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 13064 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 18216 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 23368 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 28520 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 33672 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 5336 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 10488 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 15640 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 20792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 25944 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 31096 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 7912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 13064 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 18216 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 23368 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 28520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 33672 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 5336 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 10488 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 15640 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 20792 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 25944 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 31096 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 7912 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 13064 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 18216 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 23368 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 28520 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 33672 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 5336 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 10488 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 15640 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 20792 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 25944 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 31096 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 7912 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13064 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 18216 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 23368 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 28520 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 33672 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 5336 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 10488 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 15640 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 20792 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 25944 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 31096 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 7912 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13064 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 18216 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 23368 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 28520 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 33672 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 5336 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 10488 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 15640 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 20792 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 25944 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 31096 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 7912 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 13064 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 18216 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 23368 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 28520 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 33672 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 5336 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 10488 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 15640 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 20792 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 25944 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 31096 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 7912 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13064 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 18216 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 23368 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 28520 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 33672 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 5336 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 10488 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 15640 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 20792 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 25944 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 31096 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 7912 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 13064 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 18216 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 23368 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 28520 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 33672 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 5336 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 10488 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 15640 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 20792 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 25944 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 31096 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 7912 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 13064 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 18216 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 23368 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 28520 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 33672 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 5336 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 10488 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 15640 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 25944 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 31096 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 7912 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13064 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 18216 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 23368 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 28520 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 33672 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 5336 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 10488 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 15640 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 20792 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 25944 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 31096 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 7912 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 13064 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 18216 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 23368 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 28520 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 33672 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 5336 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 10488 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 15640 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 20792 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 25944 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 31096 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 7912 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13064 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 18216 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 23368 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 28520 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 33672 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 5336 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 10488 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 15640 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 20792 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 25944 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 31096 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 7912 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 13064 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 18216 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 23368 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 28520 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 33672 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 5336 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 10488 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 15640 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 20792 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 25944 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 31096 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 7912 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 13064 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 18216 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 23368 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 28520 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 33672 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 5336 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 10488 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 15640 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 20792 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 25944 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 31096 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 7912 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13064 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 18216 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 23368 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 28520 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 33672 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 5336 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 10488 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 15640 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 20792 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 25944 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 31096 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 7912 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13064 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 18216 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 23368 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 28520 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 33672 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 5336 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 10488 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 15640 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 20792 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 25944 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 31096 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 7912 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 13064 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 18216 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 23368 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 28520 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 33672 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 5336 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 10488 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 15640 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 20792 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 25944 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 31096 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 7912 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 13064 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 18216 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 23368 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 28520 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 33672 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 5336 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 10488 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 15640 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 20792 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 25944 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 31096 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 7912 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13064 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 18216 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 23368 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 28520 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 33672 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 5336 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 10488 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 15640 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 20792 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 25944 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 31096 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 7912 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 13064 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 18216 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 23368 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 28520 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 33672 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 5336 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 10488 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 15640 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 20792 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 25944 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 31096 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 7912 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 13064 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 18216 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 23368 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 28520 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 33672 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 5336 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 10488 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 15640 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 20792 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 25944 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 31096 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 7912 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 13064 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 18216 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 23368 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 28520 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 33672 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 5336 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 10488 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 15640 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 20792 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 25944 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 31096 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 7912 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 13064 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 18216 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 23368 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 28520 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 33672 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 5336 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 10488 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 15640 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 20792 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 25944 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 31096 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 7912 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 13064 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 18216 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 23368 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 28520 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 33672 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 5336 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 10488 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 15640 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 20792 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 25944 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 31096 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 7912 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 13064 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 18216 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 23368 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 28520 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 33672 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 5336 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 10488 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 15640 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 20792 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 25944 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 31096 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 7912 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 13064 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 18216 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 23368 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 28520 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 33672 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 5336 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 10488 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 15640 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 20792 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 25944 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 31096 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 5336 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 7912 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 10488 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 13064 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 15640 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 18216 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 23368 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 25944 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 28520 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 31096 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 33672 0 -1 34272
box -38 -48 130 592
<< labels >>
flabel metal2 s 11610 35678 11666 36478 0 FreeSans 224 90 0 0 clk
port 0 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 i_start_rx
port 1 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 i_uart_rx
port 2 nsew signal input
flabel metal2 s 19982 35678 20038 36478 0 FreeSans 224 90 0 0 o_uart_tx
port 3 nsew signal tristate
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 rst
port 4 nsew signal input
flabel metal4 s 6544 2672 6864 34320 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 14433 2672 14753 34320 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 22322 2672 22642 34320 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 30211 2672 30531 34320 0 FreeSans 1920 90 0 0 vccd1
port 5 nsew power bidirectional
flabel metal4 s 7204 2672 7524 34320 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 15093 2672 15413 34320 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 22982 2672 23302 34320 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal4 s 30871 2672 31191 34320 0 FreeSans 1920 90 0 0 vssd1
port 6 nsew ground bidirectional
flabel metal3 s 36302 12248 37102 12368 0 FreeSans 480 0 0 0 wb_ack_i
port 7 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 wb_adr_o[0]
port 8 nsew signal tristate
flabel metal2 s 23846 35678 23902 36478 0 FreeSans 224 90 0 0 wb_adr_o[10]
port 9 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 wb_adr_o[11]
port 10 nsew signal tristate
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 wb_adr_o[12]
port 11 nsew signal tristate
flabel metal3 s 36302 28568 37102 28688 0 FreeSans 480 0 0 0 wb_adr_o[13]
port 12 nsew signal tristate
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 wb_adr_o[14]
port 13 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 wb_adr_o[15]
port 14 nsew signal tristate
flabel metal3 s 36302 6808 37102 6928 0 FreeSans 480 0 0 0 wb_adr_o[16]
port 15 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 wb_adr_o[17]
port 16 nsew signal tristate
flabel metal3 s 36302 18368 37102 18488 0 FreeSans 480 0 0 0 wb_adr_o[18]
port 17 nsew signal tristate
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 wb_adr_o[19]
port 18 nsew signal tristate
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 wb_adr_o[1]
port 19 nsew signal tristate
flabel metal2 s 32218 35678 32274 36478 0 FreeSans 224 90 0 0 wb_adr_o[20]
port 20 nsew signal tristate
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 wb_adr_o[21]
port 21 nsew signal tristate
flabel metal3 s 36302 5448 37102 5568 0 FreeSans 480 0 0 0 wb_adr_o[22]
port 22 nsew signal tristate
flabel metal3 s 36302 19728 37102 19848 0 FreeSans 480 0 0 0 wb_adr_o[23]
port 23 nsew signal tristate
flabel metal3 s 36302 32648 37102 32768 0 FreeSans 480 0 0 0 wb_adr_o[24]
port 24 nsew signal tristate
flabel metal2 s 4526 35678 4582 36478 0 FreeSans 224 90 0 0 wb_adr_o[25]
port 25 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 wb_adr_o[26]
port 26 nsew signal tristate
flabel metal2 s 26422 35678 26478 36478 0 FreeSans 224 90 0 0 wb_adr_o[27]
port 27 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wb_adr_o[28]
port 28 nsew signal tristate
flabel metal2 s 34794 35678 34850 36478 0 FreeSans 224 90 0 0 wb_adr_o[29]
port 29 nsew signal tristate
flabel metal3 s 36302 34008 37102 34128 0 FreeSans 480 0 0 0 wb_adr_o[2]
port 30 nsew signal tristate
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 wb_adr_o[30]
port 31 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 wb_adr_o[31]
port 32 nsew signal tristate
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 wb_adr_o[3]
port 33 nsew signal tristate
flabel metal3 s 36302 35368 37102 35488 0 FreeSans 480 0 0 0 wb_adr_o[4]
port 34 nsew signal tristate
flabel metal2 s 30930 35678 30986 36478 0 FreeSans 224 90 0 0 wb_adr_o[5]
port 35 nsew signal tristate
flabel metal3 s 36302 688 37102 808 0 FreeSans 480 0 0 0 wb_adr_o[6]
port 36 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 wb_adr_o[7]
port 37 nsew signal tristate
flabel metal3 s 36302 15648 37102 15768 0 FreeSans 480 0 0 0 wb_adr_o[8]
port 38 nsew signal tristate
flabel metal3 s 36302 10888 37102 11008 0 FreeSans 480 0 0 0 wb_adr_o[9]
port 39 nsew signal tristate
flabel metal2 s 12898 35678 12954 36478 0 FreeSans 224 90 0 0 wb_cyc_o
port 40 nsew signal tristate
flabel metal2 s 14186 35678 14242 36478 0 FreeSans 224 90 0 0 wb_dat_i[0]
port 41 nsew signal input
flabel metal3 s 36302 27208 37102 27328 0 FreeSans 480 0 0 0 wb_dat_i[10]
port 42 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 wb_dat_i[11]
port 43 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 wb_dat_i[12]
port 44 nsew signal input
flabel metal3 s 36302 29928 37102 30048 0 FreeSans 480 0 0 0 wb_dat_i[13]
port 45 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 wb_dat_i[14]
port 46 nsew signal input
flabel metal2 s 21270 35678 21326 36478 0 FreeSans 224 90 0 0 wb_dat_i[15]
port 47 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 wb_dat_i[16]
port 48 nsew signal input
flabel metal2 s 10322 35678 10378 36478 0 FreeSans 224 90 0 0 wb_dat_i[17]
port 49 nsew signal input
flabel metal2 s 15474 35678 15530 36478 0 FreeSans 224 90 0 0 wb_dat_i[18]
port 50 nsew signal input
flabel metal3 s 36302 31288 37102 31408 0 FreeSans 480 0 0 0 wb_dat_i[19]
port 51 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 wb_dat_i[1]
port 52 nsew signal input
flabel metal2 s 18694 35678 18750 36478 0 FreeSans 224 90 0 0 wb_dat_i[20]
port 53 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 wb_dat_i[21]
port 54 nsew signal input
flabel metal3 s 36302 8168 37102 8288 0 FreeSans 480 0 0 0 wb_dat_i[22]
port 55 nsew signal input
flabel metal3 s 36302 22448 37102 22568 0 FreeSans 480 0 0 0 wb_dat_i[23]
port 56 nsew signal input
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 wb_dat_i[24]
port 57 nsew signal input
flabel metal2 s 22558 35678 22614 36478 0 FreeSans 224 90 0 0 wb_dat_i[25]
port 58 nsew signal input
flabel metal2 s 7746 35678 7802 36478 0 FreeSans 224 90 0 0 wb_dat_i[26]
port 59 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 wb_dat_i[27]
port 60 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 wb_dat_i[28]
port 61 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 wb_dat_i[29]
port 62 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 wb_dat_i[2]
port 63 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 wb_dat_i[30]
port 64 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 wb_dat_i[31]
port 65 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 wb_dat_i[3]
port 66 nsew signal input
flabel metal3 s 36302 9528 37102 9648 0 FreeSans 480 0 0 0 wb_dat_i[4]
port 67 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 wb_dat_i[5]
port 68 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 wb_dat_i[6]
port 69 nsew signal input
flabel metal3 s 36302 2048 37102 2168 0 FreeSans 480 0 0 0 wb_dat_i[7]
port 70 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 wb_dat_i[8]
port 71 nsew signal input
flabel metal3 s 36302 13608 37102 13728 0 FreeSans 480 0 0 0 wb_dat_i[9]
port 72 nsew signal input
flabel metal3 s 36302 23808 37102 23928 0 FreeSans 480 0 0 0 wb_dat_o[0]
port 73 nsew signal tristate
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 wb_dat_o[10]
port 74 nsew signal tristate
flabel metal3 s 36302 25848 37102 25968 0 FreeSans 480 0 0 0 wb_dat_o[11]
port 75 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 wb_dat_o[12]
port 76 nsew signal tristate
flabel metal2 s 662 35678 718 36478 0 FreeSans 224 90 0 0 wb_dat_o[13]
port 77 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 wb_dat_o[14]
port 78 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 wb_dat_o[15]
port 79 nsew signal tristate
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 wb_dat_o[16]
port 80 nsew signal tristate
flabel metal2 s 5814 35678 5870 36478 0 FreeSans 224 90 0 0 wb_dat_o[17]
port 81 nsew signal tristate
flabel metal2 s 17406 35678 17462 36478 0 FreeSans 224 90 0 0 wb_dat_o[18]
port 82 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 wb_dat_o[19]
port 83 nsew signal tristate
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 wb_dat_o[1]
port 84 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 wb_dat_o[20]
port 85 nsew signal tristate
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 wb_dat_o[21]
port 86 nsew signal tristate
flabel metal2 s 33506 35678 33562 36478 0 FreeSans 224 90 0 0 wb_dat_o[22]
port 87 nsew signal tristate
flabel metal2 s 25134 35678 25190 36478 0 FreeSans 224 90 0 0 wb_dat_o[23]
port 88 nsew signal tristate
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 wb_dat_o[24]
port 89 nsew signal tristate
flabel metal2 s 36082 35678 36138 36478 0 FreeSans 224 90 0 0 wb_dat_o[25]
port 90 nsew signal tristate
flabel metal3 s 36302 4088 37102 4208 0 FreeSans 480 0 0 0 wb_dat_o[26]
port 91 nsew signal tristate
flabel metal2 s 1950 35678 2006 36478 0 FreeSans 224 90 0 0 wb_dat_o[27]
port 92 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 wb_dat_o[28]
port 93 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 wb_dat_o[29]
port 94 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 wb_dat_o[2]
port 95 nsew signal tristate
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 wb_dat_o[30]
port 96 nsew signal tristate
flabel metal3 s 36302 21088 37102 21208 0 FreeSans 480 0 0 0 wb_dat_o[31]
port 97 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 wb_dat_o[3]
port 98 nsew signal tristate
flabel metal2 s 29642 35678 29698 36478 0 FreeSans 224 90 0 0 wb_dat_o[4]
port 99 nsew signal tristate
flabel metal2 s 28354 35678 28410 36478 0 FreeSans 224 90 0 0 wb_dat_o[5]
port 100 nsew signal tristate
flabel metal2 s 3238 35678 3294 36478 0 FreeSans 224 90 0 0 wb_dat_o[6]
port 101 nsew signal tristate
flabel metal2 s 9034 35678 9090 36478 0 FreeSans 224 90 0 0 wb_dat_o[7]
port 102 nsew signal tristate
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 wb_dat_o[8]
port 103 nsew signal tristate
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 wb_dat_o[9]
port 104 nsew signal tristate
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 wb_stb_o
port 105 nsew signal tristate
flabel metal3 s 36302 17008 37102 17128 0 FreeSans 480 0 0 0 wb_we_o
port 106 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 37102 36478
<< end >>
