// This is the unpowered netlist.
module mem (clk,
    rst,
    wb_ack_o,
    wb_cyc_i,
    wb_stb_i,
    wb_we_i,
    wb_adr_i,
    wb_dat_i,
    wb_dat_o);
 input clk;
 input rst;
 output wb_ack_o;
 input wb_cyc_i;
 input wb_stb_i;
 input wb_we_i;
 input [4:0] wb_adr_i;
 input [31:0] wb_dat_i;
 output [31:0] wb_dat_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_9_clk;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][16] ;
 wire \mem[0][17] ;
 wire \mem[0][18] ;
 wire \mem[0][19] ;
 wire \mem[0][1] ;
 wire \mem[0][20] ;
 wire \mem[0][21] ;
 wire \mem[0][22] ;
 wire \mem[0][23] ;
 wire \mem[0][24] ;
 wire \mem[0][25] ;
 wire \mem[0][26] ;
 wire \mem[0][27] ;
 wire \mem[0][28] ;
 wire \mem[0][29] ;
 wire \mem[0][2] ;
 wire \mem[0][30] ;
 wire \mem[0][31] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][16] ;
 wire \mem[10][17] ;
 wire \mem[10][18] ;
 wire \mem[10][19] ;
 wire \mem[10][1] ;
 wire \mem[10][20] ;
 wire \mem[10][21] ;
 wire \mem[10][22] ;
 wire \mem[10][23] ;
 wire \mem[10][24] ;
 wire \mem[10][25] ;
 wire \mem[10][26] ;
 wire \mem[10][27] ;
 wire \mem[10][28] ;
 wire \mem[10][29] ;
 wire \mem[10][2] ;
 wire \mem[10][30] ;
 wire \mem[10][31] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][16] ;
 wire \mem[11][17] ;
 wire \mem[11][18] ;
 wire \mem[11][19] ;
 wire \mem[11][1] ;
 wire \mem[11][20] ;
 wire \mem[11][21] ;
 wire \mem[11][22] ;
 wire \mem[11][23] ;
 wire \mem[11][24] ;
 wire \mem[11][25] ;
 wire \mem[11][26] ;
 wire \mem[11][27] ;
 wire \mem[11][28] ;
 wire \mem[11][29] ;
 wire \mem[11][2] ;
 wire \mem[11][30] ;
 wire \mem[11][31] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][16] ;
 wire \mem[12][17] ;
 wire \mem[12][18] ;
 wire \mem[12][19] ;
 wire \mem[12][1] ;
 wire \mem[12][20] ;
 wire \mem[12][21] ;
 wire \mem[12][22] ;
 wire \mem[12][23] ;
 wire \mem[12][24] ;
 wire \mem[12][25] ;
 wire \mem[12][26] ;
 wire \mem[12][27] ;
 wire \mem[12][28] ;
 wire \mem[12][29] ;
 wire \mem[12][2] ;
 wire \mem[12][30] ;
 wire \mem[12][31] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][16] ;
 wire \mem[13][17] ;
 wire \mem[13][18] ;
 wire \mem[13][19] ;
 wire \mem[13][1] ;
 wire \mem[13][20] ;
 wire \mem[13][21] ;
 wire \mem[13][22] ;
 wire \mem[13][23] ;
 wire \mem[13][24] ;
 wire \mem[13][25] ;
 wire \mem[13][26] ;
 wire \mem[13][27] ;
 wire \mem[13][28] ;
 wire \mem[13][29] ;
 wire \mem[13][2] ;
 wire \mem[13][30] ;
 wire \mem[13][31] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][16] ;
 wire \mem[14][17] ;
 wire \mem[14][18] ;
 wire \mem[14][19] ;
 wire \mem[14][1] ;
 wire \mem[14][20] ;
 wire \mem[14][21] ;
 wire \mem[14][22] ;
 wire \mem[14][23] ;
 wire \mem[14][24] ;
 wire \mem[14][25] ;
 wire \mem[14][26] ;
 wire \mem[14][27] ;
 wire \mem[14][28] ;
 wire \mem[14][29] ;
 wire \mem[14][2] ;
 wire \mem[14][30] ;
 wire \mem[14][31] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][16] ;
 wire \mem[15][17] ;
 wire \mem[15][18] ;
 wire \mem[15][19] ;
 wire \mem[15][1] ;
 wire \mem[15][20] ;
 wire \mem[15][21] ;
 wire \mem[15][22] ;
 wire \mem[15][23] ;
 wire \mem[15][24] ;
 wire \mem[15][25] ;
 wire \mem[15][26] ;
 wire \mem[15][27] ;
 wire \mem[15][28] ;
 wire \mem[15][29] ;
 wire \mem[15][2] ;
 wire \mem[15][30] ;
 wire \mem[15][31] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[16][0] ;
 wire \mem[16][10] ;
 wire \mem[16][11] ;
 wire \mem[16][12] ;
 wire \mem[16][13] ;
 wire \mem[16][14] ;
 wire \mem[16][15] ;
 wire \mem[16][16] ;
 wire \mem[16][17] ;
 wire \mem[16][18] ;
 wire \mem[16][19] ;
 wire \mem[16][1] ;
 wire \mem[16][20] ;
 wire \mem[16][21] ;
 wire \mem[16][22] ;
 wire \mem[16][23] ;
 wire \mem[16][24] ;
 wire \mem[16][25] ;
 wire \mem[16][26] ;
 wire \mem[16][27] ;
 wire \mem[16][28] ;
 wire \mem[16][29] ;
 wire \mem[16][2] ;
 wire \mem[16][30] ;
 wire \mem[16][31] ;
 wire \mem[16][3] ;
 wire \mem[16][4] ;
 wire \mem[16][5] ;
 wire \mem[16][6] ;
 wire \mem[16][7] ;
 wire \mem[16][8] ;
 wire \mem[16][9] ;
 wire \mem[17][0] ;
 wire \mem[17][10] ;
 wire \mem[17][11] ;
 wire \mem[17][12] ;
 wire \mem[17][13] ;
 wire \mem[17][14] ;
 wire \mem[17][15] ;
 wire \mem[17][16] ;
 wire \mem[17][17] ;
 wire \mem[17][18] ;
 wire \mem[17][19] ;
 wire \mem[17][1] ;
 wire \mem[17][20] ;
 wire \mem[17][21] ;
 wire \mem[17][22] ;
 wire \mem[17][23] ;
 wire \mem[17][24] ;
 wire \mem[17][25] ;
 wire \mem[17][26] ;
 wire \mem[17][27] ;
 wire \mem[17][28] ;
 wire \mem[17][29] ;
 wire \mem[17][2] ;
 wire \mem[17][30] ;
 wire \mem[17][31] ;
 wire \mem[17][3] ;
 wire \mem[17][4] ;
 wire \mem[17][5] ;
 wire \mem[17][6] ;
 wire \mem[17][7] ;
 wire \mem[17][8] ;
 wire \mem[17][9] ;
 wire \mem[18][0] ;
 wire \mem[18][10] ;
 wire \mem[18][11] ;
 wire \mem[18][12] ;
 wire \mem[18][13] ;
 wire \mem[18][14] ;
 wire \mem[18][15] ;
 wire \mem[18][16] ;
 wire \mem[18][17] ;
 wire \mem[18][18] ;
 wire \mem[18][19] ;
 wire \mem[18][1] ;
 wire \mem[18][20] ;
 wire \mem[18][21] ;
 wire \mem[18][22] ;
 wire \mem[18][23] ;
 wire \mem[18][24] ;
 wire \mem[18][25] ;
 wire \mem[18][26] ;
 wire \mem[18][27] ;
 wire \mem[18][28] ;
 wire \mem[18][29] ;
 wire \mem[18][2] ;
 wire \mem[18][30] ;
 wire \mem[18][31] ;
 wire \mem[18][3] ;
 wire \mem[18][4] ;
 wire \mem[18][5] ;
 wire \mem[18][6] ;
 wire \mem[18][7] ;
 wire \mem[18][8] ;
 wire \mem[18][9] ;
 wire \mem[19][0] ;
 wire \mem[19][10] ;
 wire \mem[19][11] ;
 wire \mem[19][12] ;
 wire \mem[19][13] ;
 wire \mem[19][14] ;
 wire \mem[19][15] ;
 wire \mem[19][16] ;
 wire \mem[19][17] ;
 wire \mem[19][18] ;
 wire \mem[19][19] ;
 wire \mem[19][1] ;
 wire \mem[19][20] ;
 wire \mem[19][21] ;
 wire \mem[19][22] ;
 wire \mem[19][23] ;
 wire \mem[19][24] ;
 wire \mem[19][25] ;
 wire \mem[19][26] ;
 wire \mem[19][27] ;
 wire \mem[19][28] ;
 wire \mem[19][29] ;
 wire \mem[19][2] ;
 wire \mem[19][30] ;
 wire \mem[19][31] ;
 wire \mem[19][3] ;
 wire \mem[19][4] ;
 wire \mem[19][5] ;
 wire \mem[19][6] ;
 wire \mem[19][7] ;
 wire \mem[19][8] ;
 wire \mem[19][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][16] ;
 wire \mem[1][17] ;
 wire \mem[1][18] ;
 wire \mem[1][19] ;
 wire \mem[1][1] ;
 wire \mem[1][20] ;
 wire \mem[1][21] ;
 wire \mem[1][22] ;
 wire \mem[1][23] ;
 wire \mem[1][24] ;
 wire \mem[1][25] ;
 wire \mem[1][26] ;
 wire \mem[1][27] ;
 wire \mem[1][28] ;
 wire \mem[1][29] ;
 wire \mem[1][2] ;
 wire \mem[1][30] ;
 wire \mem[1][31] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[20][0] ;
 wire \mem[20][10] ;
 wire \mem[20][11] ;
 wire \mem[20][12] ;
 wire \mem[20][13] ;
 wire \mem[20][14] ;
 wire \mem[20][15] ;
 wire \mem[20][16] ;
 wire \mem[20][17] ;
 wire \mem[20][18] ;
 wire \mem[20][19] ;
 wire \mem[20][1] ;
 wire \mem[20][20] ;
 wire \mem[20][21] ;
 wire \mem[20][22] ;
 wire \mem[20][23] ;
 wire \mem[20][24] ;
 wire \mem[20][25] ;
 wire \mem[20][26] ;
 wire \mem[20][27] ;
 wire \mem[20][28] ;
 wire \mem[20][29] ;
 wire \mem[20][2] ;
 wire \mem[20][30] ;
 wire \mem[20][31] ;
 wire \mem[20][3] ;
 wire \mem[20][4] ;
 wire \mem[20][5] ;
 wire \mem[20][6] ;
 wire \mem[20][7] ;
 wire \mem[20][8] ;
 wire \mem[20][9] ;
 wire \mem[21][0] ;
 wire \mem[21][10] ;
 wire \mem[21][11] ;
 wire \mem[21][12] ;
 wire \mem[21][13] ;
 wire \mem[21][14] ;
 wire \mem[21][15] ;
 wire \mem[21][16] ;
 wire \mem[21][17] ;
 wire \mem[21][18] ;
 wire \mem[21][19] ;
 wire \mem[21][1] ;
 wire \mem[21][20] ;
 wire \mem[21][21] ;
 wire \mem[21][22] ;
 wire \mem[21][23] ;
 wire \mem[21][24] ;
 wire \mem[21][25] ;
 wire \mem[21][26] ;
 wire \mem[21][27] ;
 wire \mem[21][28] ;
 wire \mem[21][29] ;
 wire \mem[21][2] ;
 wire \mem[21][30] ;
 wire \mem[21][31] ;
 wire \mem[21][3] ;
 wire \mem[21][4] ;
 wire \mem[21][5] ;
 wire \mem[21][6] ;
 wire \mem[21][7] ;
 wire \mem[21][8] ;
 wire \mem[21][9] ;
 wire \mem[22][0] ;
 wire \mem[22][10] ;
 wire \mem[22][11] ;
 wire \mem[22][12] ;
 wire \mem[22][13] ;
 wire \mem[22][14] ;
 wire \mem[22][15] ;
 wire \mem[22][16] ;
 wire \mem[22][17] ;
 wire \mem[22][18] ;
 wire \mem[22][19] ;
 wire \mem[22][1] ;
 wire \mem[22][20] ;
 wire \mem[22][21] ;
 wire \mem[22][22] ;
 wire \mem[22][23] ;
 wire \mem[22][24] ;
 wire \mem[22][25] ;
 wire \mem[22][26] ;
 wire \mem[22][27] ;
 wire \mem[22][28] ;
 wire \mem[22][29] ;
 wire \mem[22][2] ;
 wire \mem[22][30] ;
 wire \mem[22][31] ;
 wire \mem[22][3] ;
 wire \mem[22][4] ;
 wire \mem[22][5] ;
 wire \mem[22][6] ;
 wire \mem[22][7] ;
 wire \mem[22][8] ;
 wire \mem[22][9] ;
 wire \mem[23][0] ;
 wire \mem[23][10] ;
 wire \mem[23][11] ;
 wire \mem[23][12] ;
 wire \mem[23][13] ;
 wire \mem[23][14] ;
 wire \mem[23][15] ;
 wire \mem[23][16] ;
 wire \mem[23][17] ;
 wire \mem[23][18] ;
 wire \mem[23][19] ;
 wire \mem[23][1] ;
 wire \mem[23][20] ;
 wire \mem[23][21] ;
 wire \mem[23][22] ;
 wire \mem[23][23] ;
 wire \mem[23][24] ;
 wire \mem[23][25] ;
 wire \mem[23][26] ;
 wire \mem[23][27] ;
 wire \mem[23][28] ;
 wire \mem[23][29] ;
 wire \mem[23][2] ;
 wire \mem[23][30] ;
 wire \mem[23][31] ;
 wire \mem[23][3] ;
 wire \mem[23][4] ;
 wire \mem[23][5] ;
 wire \mem[23][6] ;
 wire \mem[23][7] ;
 wire \mem[23][8] ;
 wire \mem[23][9] ;
 wire \mem[24][0] ;
 wire \mem[24][10] ;
 wire \mem[24][11] ;
 wire \mem[24][12] ;
 wire \mem[24][13] ;
 wire \mem[24][14] ;
 wire \mem[24][15] ;
 wire \mem[24][16] ;
 wire \mem[24][17] ;
 wire \mem[24][18] ;
 wire \mem[24][19] ;
 wire \mem[24][1] ;
 wire \mem[24][20] ;
 wire \mem[24][21] ;
 wire \mem[24][22] ;
 wire \mem[24][23] ;
 wire \mem[24][24] ;
 wire \mem[24][25] ;
 wire \mem[24][26] ;
 wire \mem[24][27] ;
 wire \mem[24][28] ;
 wire \mem[24][29] ;
 wire \mem[24][2] ;
 wire \mem[24][30] ;
 wire \mem[24][31] ;
 wire \mem[24][3] ;
 wire \mem[24][4] ;
 wire \mem[24][5] ;
 wire \mem[24][6] ;
 wire \mem[24][7] ;
 wire \mem[24][8] ;
 wire \mem[24][9] ;
 wire \mem[25][0] ;
 wire \mem[25][10] ;
 wire \mem[25][11] ;
 wire \mem[25][12] ;
 wire \mem[25][13] ;
 wire \mem[25][14] ;
 wire \mem[25][15] ;
 wire \mem[25][16] ;
 wire \mem[25][17] ;
 wire \mem[25][18] ;
 wire \mem[25][19] ;
 wire \mem[25][1] ;
 wire \mem[25][20] ;
 wire \mem[25][21] ;
 wire \mem[25][22] ;
 wire \mem[25][23] ;
 wire \mem[25][24] ;
 wire \mem[25][25] ;
 wire \mem[25][26] ;
 wire \mem[25][27] ;
 wire \mem[25][28] ;
 wire \mem[25][29] ;
 wire \mem[25][2] ;
 wire \mem[25][30] ;
 wire \mem[25][31] ;
 wire \mem[25][3] ;
 wire \mem[25][4] ;
 wire \mem[25][5] ;
 wire \mem[25][6] ;
 wire \mem[25][7] ;
 wire \mem[25][8] ;
 wire \mem[25][9] ;
 wire \mem[26][0] ;
 wire \mem[26][10] ;
 wire \mem[26][11] ;
 wire \mem[26][12] ;
 wire \mem[26][13] ;
 wire \mem[26][14] ;
 wire \mem[26][15] ;
 wire \mem[26][16] ;
 wire \mem[26][17] ;
 wire \mem[26][18] ;
 wire \mem[26][19] ;
 wire \mem[26][1] ;
 wire \mem[26][20] ;
 wire \mem[26][21] ;
 wire \mem[26][22] ;
 wire \mem[26][23] ;
 wire \mem[26][24] ;
 wire \mem[26][25] ;
 wire \mem[26][26] ;
 wire \mem[26][27] ;
 wire \mem[26][28] ;
 wire \mem[26][29] ;
 wire \mem[26][2] ;
 wire \mem[26][30] ;
 wire \mem[26][31] ;
 wire \mem[26][3] ;
 wire \mem[26][4] ;
 wire \mem[26][5] ;
 wire \mem[26][6] ;
 wire \mem[26][7] ;
 wire \mem[26][8] ;
 wire \mem[26][9] ;
 wire \mem[27][0] ;
 wire \mem[27][10] ;
 wire \mem[27][11] ;
 wire \mem[27][12] ;
 wire \mem[27][13] ;
 wire \mem[27][14] ;
 wire \mem[27][15] ;
 wire \mem[27][16] ;
 wire \mem[27][17] ;
 wire \mem[27][18] ;
 wire \mem[27][19] ;
 wire \mem[27][1] ;
 wire \mem[27][20] ;
 wire \mem[27][21] ;
 wire \mem[27][22] ;
 wire \mem[27][23] ;
 wire \mem[27][24] ;
 wire \mem[27][25] ;
 wire \mem[27][26] ;
 wire \mem[27][27] ;
 wire \mem[27][28] ;
 wire \mem[27][29] ;
 wire \mem[27][2] ;
 wire \mem[27][30] ;
 wire \mem[27][31] ;
 wire \mem[27][3] ;
 wire \mem[27][4] ;
 wire \mem[27][5] ;
 wire \mem[27][6] ;
 wire \mem[27][7] ;
 wire \mem[27][8] ;
 wire \mem[27][9] ;
 wire \mem[28][0] ;
 wire \mem[28][10] ;
 wire \mem[28][11] ;
 wire \mem[28][12] ;
 wire \mem[28][13] ;
 wire \mem[28][14] ;
 wire \mem[28][15] ;
 wire \mem[28][16] ;
 wire \mem[28][17] ;
 wire \mem[28][18] ;
 wire \mem[28][19] ;
 wire \mem[28][1] ;
 wire \mem[28][20] ;
 wire \mem[28][21] ;
 wire \mem[28][22] ;
 wire \mem[28][23] ;
 wire \mem[28][24] ;
 wire \mem[28][25] ;
 wire \mem[28][26] ;
 wire \mem[28][27] ;
 wire \mem[28][28] ;
 wire \mem[28][29] ;
 wire \mem[28][2] ;
 wire \mem[28][30] ;
 wire \mem[28][31] ;
 wire \mem[28][3] ;
 wire \mem[28][4] ;
 wire \mem[28][5] ;
 wire \mem[28][6] ;
 wire \mem[28][7] ;
 wire \mem[28][8] ;
 wire \mem[28][9] ;
 wire \mem[29][0] ;
 wire \mem[29][10] ;
 wire \mem[29][11] ;
 wire \mem[29][12] ;
 wire \mem[29][13] ;
 wire \mem[29][14] ;
 wire \mem[29][15] ;
 wire \mem[29][16] ;
 wire \mem[29][17] ;
 wire \mem[29][18] ;
 wire \mem[29][19] ;
 wire \mem[29][1] ;
 wire \mem[29][20] ;
 wire \mem[29][21] ;
 wire \mem[29][22] ;
 wire \mem[29][23] ;
 wire \mem[29][24] ;
 wire \mem[29][25] ;
 wire \mem[29][26] ;
 wire \mem[29][27] ;
 wire \mem[29][28] ;
 wire \mem[29][29] ;
 wire \mem[29][2] ;
 wire \mem[29][30] ;
 wire \mem[29][31] ;
 wire \mem[29][3] ;
 wire \mem[29][4] ;
 wire \mem[29][5] ;
 wire \mem[29][6] ;
 wire \mem[29][7] ;
 wire \mem[29][8] ;
 wire \mem[29][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][16] ;
 wire \mem[2][17] ;
 wire \mem[2][18] ;
 wire \mem[2][19] ;
 wire \mem[2][1] ;
 wire \mem[2][20] ;
 wire \mem[2][21] ;
 wire \mem[2][22] ;
 wire \mem[2][23] ;
 wire \mem[2][24] ;
 wire \mem[2][25] ;
 wire \mem[2][26] ;
 wire \mem[2][27] ;
 wire \mem[2][28] ;
 wire \mem[2][29] ;
 wire \mem[2][2] ;
 wire \mem[2][30] ;
 wire \mem[2][31] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[30][0] ;
 wire \mem[30][10] ;
 wire \mem[30][11] ;
 wire \mem[30][12] ;
 wire \mem[30][13] ;
 wire \mem[30][14] ;
 wire \mem[30][15] ;
 wire \mem[30][16] ;
 wire \mem[30][17] ;
 wire \mem[30][18] ;
 wire \mem[30][19] ;
 wire \mem[30][1] ;
 wire \mem[30][20] ;
 wire \mem[30][21] ;
 wire \mem[30][22] ;
 wire \mem[30][23] ;
 wire \mem[30][24] ;
 wire \mem[30][25] ;
 wire \mem[30][26] ;
 wire \mem[30][27] ;
 wire \mem[30][28] ;
 wire \mem[30][29] ;
 wire \mem[30][2] ;
 wire \mem[30][30] ;
 wire \mem[30][31] ;
 wire \mem[30][3] ;
 wire \mem[30][4] ;
 wire \mem[30][5] ;
 wire \mem[30][6] ;
 wire \mem[30][7] ;
 wire \mem[30][8] ;
 wire \mem[30][9] ;
 wire \mem[31][0] ;
 wire \mem[31][10] ;
 wire \mem[31][11] ;
 wire \mem[31][12] ;
 wire \mem[31][13] ;
 wire \mem[31][14] ;
 wire \mem[31][15] ;
 wire \mem[31][16] ;
 wire \mem[31][17] ;
 wire \mem[31][18] ;
 wire \mem[31][19] ;
 wire \mem[31][1] ;
 wire \mem[31][20] ;
 wire \mem[31][21] ;
 wire \mem[31][22] ;
 wire \mem[31][23] ;
 wire \mem[31][24] ;
 wire \mem[31][25] ;
 wire \mem[31][26] ;
 wire \mem[31][27] ;
 wire \mem[31][28] ;
 wire \mem[31][29] ;
 wire \mem[31][2] ;
 wire \mem[31][30] ;
 wire \mem[31][31] ;
 wire \mem[31][3] ;
 wire \mem[31][4] ;
 wire \mem[31][5] ;
 wire \mem[31][6] ;
 wire \mem[31][7] ;
 wire \mem[31][8] ;
 wire \mem[31][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][16] ;
 wire \mem[3][17] ;
 wire \mem[3][18] ;
 wire \mem[3][19] ;
 wire \mem[3][1] ;
 wire \mem[3][20] ;
 wire \mem[3][21] ;
 wire \mem[3][22] ;
 wire \mem[3][23] ;
 wire \mem[3][24] ;
 wire \mem[3][25] ;
 wire \mem[3][26] ;
 wire \mem[3][27] ;
 wire \mem[3][28] ;
 wire \mem[3][29] ;
 wire \mem[3][2] ;
 wire \mem[3][30] ;
 wire \mem[3][31] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][16] ;
 wire \mem[4][17] ;
 wire \mem[4][18] ;
 wire \mem[4][19] ;
 wire \mem[4][1] ;
 wire \mem[4][20] ;
 wire \mem[4][21] ;
 wire \mem[4][22] ;
 wire \mem[4][23] ;
 wire \mem[4][24] ;
 wire \mem[4][25] ;
 wire \mem[4][26] ;
 wire \mem[4][27] ;
 wire \mem[4][28] ;
 wire \mem[4][29] ;
 wire \mem[4][2] ;
 wire \mem[4][30] ;
 wire \mem[4][31] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][16] ;
 wire \mem[5][17] ;
 wire \mem[5][18] ;
 wire \mem[5][19] ;
 wire \mem[5][1] ;
 wire \mem[5][20] ;
 wire \mem[5][21] ;
 wire \mem[5][22] ;
 wire \mem[5][23] ;
 wire \mem[5][24] ;
 wire \mem[5][25] ;
 wire \mem[5][26] ;
 wire \mem[5][27] ;
 wire \mem[5][28] ;
 wire \mem[5][29] ;
 wire \mem[5][2] ;
 wire \mem[5][30] ;
 wire \mem[5][31] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][16] ;
 wire \mem[6][17] ;
 wire \mem[6][18] ;
 wire \mem[6][19] ;
 wire \mem[6][1] ;
 wire \mem[6][20] ;
 wire \mem[6][21] ;
 wire \mem[6][22] ;
 wire \mem[6][23] ;
 wire \mem[6][24] ;
 wire \mem[6][25] ;
 wire \mem[6][26] ;
 wire \mem[6][27] ;
 wire \mem[6][28] ;
 wire \mem[6][29] ;
 wire \mem[6][2] ;
 wire \mem[6][30] ;
 wire \mem[6][31] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][16] ;
 wire \mem[7][17] ;
 wire \mem[7][18] ;
 wire \mem[7][19] ;
 wire \mem[7][1] ;
 wire \mem[7][20] ;
 wire \mem[7][21] ;
 wire \mem[7][22] ;
 wire \mem[7][23] ;
 wire \mem[7][24] ;
 wire \mem[7][25] ;
 wire \mem[7][26] ;
 wire \mem[7][27] ;
 wire \mem[7][28] ;
 wire \mem[7][29] ;
 wire \mem[7][2] ;
 wire \mem[7][30] ;
 wire \mem[7][31] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][16] ;
 wire \mem[8][17] ;
 wire \mem[8][18] ;
 wire \mem[8][19] ;
 wire \mem[8][1] ;
 wire \mem[8][20] ;
 wire \mem[8][21] ;
 wire \mem[8][22] ;
 wire \mem[8][23] ;
 wire \mem[8][24] ;
 wire \mem[8][25] ;
 wire \mem[8][26] ;
 wire \mem[8][27] ;
 wire \mem[8][28] ;
 wire \mem[8][29] ;
 wire \mem[8][2] ;
 wire \mem[8][30] ;
 wire \mem[8][31] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][16] ;
 wire \mem[9][17] ;
 wire \mem[9][18] ;
 wire \mem[9][19] ;
 wire \mem[9][1] ;
 wire \mem[9][20] ;
 wire \mem[9][21] ;
 wire \mem[9][22] ;
 wire \mem[9][23] ;
 wire \mem[9][24] ;
 wire \mem[9][25] ;
 wire \mem[9][26] ;
 wire \mem[9][27] ;
 wire \mem[9][28] ;
 wire \mem[9][29] ;
 wire \mem[9][2] ;
 wire \mem[9][30] ;
 wire \mem[9][31] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net166;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net167;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net168;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net2350;
 wire net2351;
 wire net2352;
 wire net2353;
 wire net2354;
 wire net2355;
 wire net2356;
 wire net2357;
 wire net2358;
 wire net2359;
 wire net236;
 wire net2360;
 wire net2361;
 wire net2362;
 wire net2363;
 wire net2364;
 wire net2365;
 wire net2366;
 wire net2367;
 wire net2368;
 wire net2369;
 wire net237;
 wire net2370;
 wire net2371;
 wire net2372;
 wire net2373;
 wire net2374;
 wire net2375;
 wire net2376;
 wire net2377;
 wire net2378;
 wire net2379;
 wire net238;
 wire net2380;
 wire net2381;
 wire net2382;
 wire net2383;
 wire net2384;
 wire net2385;
 wire net2386;
 wire net2387;
 wire net2388;
 wire net2389;
 wire net239;
 wire net2390;
 wire net2391;
 wire net2392;
 wire net2393;
 wire net2394;
 wire net2395;
 wire net2396;
 wire net2397;
 wire net2398;
 wire net2399;
 wire net24;
 wire net240;
 wire net2400;
 wire net2401;
 wire net2402;
 wire net2403;
 wire net2404;
 wire net2405;
 wire net2406;
 wire net2407;
 wire net2408;
 wire net2409;
 wire net241;
 wire net2410;
 wire net2411;
 wire net2412;
 wire net2413;
 wire net2414;
 wire net2415;
 wire net2416;
 wire net2417;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__1810__A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__A_N (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__1811__C (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1812__C_N (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__A_N (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__B (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1813__C (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__1814__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1815__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1816__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1817__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1818__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__1819__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1825__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1826__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1828__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__1833__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1834__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1835__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1836__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1837__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1838__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1839__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__1840__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1846__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1847__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1849__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__1854__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1855__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__1856__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__1857__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__1858__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__1859__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__1860__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__1861__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__S0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1862__S1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1863__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1864__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1865__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1866__A_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1867__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__1868__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__S0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1869__S1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1870__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__1871__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1872__A_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1873__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1874__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__1875__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__1876__C1 (.DIODE(_1074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__1877__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__1878__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__1879__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__1880__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1881__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__1882__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__1883__S1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1885__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1887__A_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1888__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1889__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1890__S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__1891__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__1892__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__1896__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__A3 (.DIODE(_1108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1897__B1 (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1900__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1901__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1902__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__1903__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1909__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1910__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1912__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__1917__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__1917__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1918__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1921__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1922__S1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1923__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__1924__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1930__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__1931__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1933__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__1938__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1939__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__1940__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__1941__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__1942__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__1943__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__1944__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__1945__B (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__1946__S1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__1948__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1950__A_N (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__1951__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__1952__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__1953__S1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1954__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__1955__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__1958__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__1959__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__1960__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__1961__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__1962__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__1963__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__1964__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__1965__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__1966__B (.DIODE(_1173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__S0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1967__S1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1968__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1969__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1970__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1971__A_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1972__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__1973__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__1974__S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__1975__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__1976__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__1977__A_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1979__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__1980__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__1981__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__1982__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__1983__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__1984__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__1985__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__1986__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__1987__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__1988__S1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1989__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__1990__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1991__S (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__1992__A_N (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__1993__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__1994__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__1995__S1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1996__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__1997__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__1998__A_N (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__1999__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2000__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2001__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2001__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2002__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2003__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2004__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2005__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2006__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2007__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2008__B (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2009__S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2010__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2012__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2014__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2015__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__S0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__2016__S1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__2017__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2018__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2020__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2022__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2023__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2024__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2025__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2026__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2027__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2028__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2029__B (.DIODE(_1233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2030__S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2032__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2035__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2036__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2037__S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2038__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2040__A_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2042__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2043__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2044__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2045__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2046__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2047__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2048__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2049__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2050__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2051__S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2052__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2054__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2056__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2057__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2058__S1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2059__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2062__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2064__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2065__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2066__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2067__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2068__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2069__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2070__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2071__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2073__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2077__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2078__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2079__S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2080__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2081__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2083__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2085__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2086__C1 (.DIODE(_1274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2087__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2088__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2089__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2090__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2091__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2092__B (.DIODE(_1293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2093__S1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2098__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2099__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2100__S1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2101__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__2103__A_N (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2104__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2105__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__A1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__2106__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2107__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2108__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2109__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2110__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2111__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__S0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2112__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__2113__B (.DIODE(_1313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__S0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2114__S1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2115__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2116__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2117__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2118__A_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2119__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__2120__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2121__S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2122__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2123__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2125__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2127__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__2128__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2129__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2130__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2131__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2132__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2133__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2134__B (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2136__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2138__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2140__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2141__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2142__S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2143__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2145__A_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2147__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2148__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2149__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2150__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2151__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2151__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2152__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2153__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__S0 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2154__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2155__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2161__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2162__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2163__S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2164__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2165__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2167__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2169__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2170__C1 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2171__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2172__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2173__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2174__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__S0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2175__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2176__B (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2177__S1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2182__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__2183__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__S0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2184__S1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2185__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__2187__A_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2188__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2189__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2190__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__A1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2191__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2192__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2193__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2194__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2195__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2196__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2197__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2203__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2204__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2205__S1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2206__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2208__A_N (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2209__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2210__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2211__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2212__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2213__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2214__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2215__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2216__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__S0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2217__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2218__B (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2224__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__2225__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__S0 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2226__S1 (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2227__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__2229__A_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2230__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2231__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__2232__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2233__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2234__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2235__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2236__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__S0 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__2237__S1 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__S0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2238__S1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2239__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2242__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2244__A_N (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2245__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2246__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2247__S1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2248__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2250__A_N (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2252__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2253__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2254__C1 (.DIODE(_1434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2255__S1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2256__S1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2257__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2258__S1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2259__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2260__B (.DIODE(_1453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2262__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2264__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2266__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2267__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2269__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2270__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2274__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2275__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2276__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2277__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2278__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2279__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2280__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2281__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2285__S (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2287__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2288__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2289__S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2290__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2291__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2293__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2295__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2296__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2297__S1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2298__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__S0 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__2299__S1 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__S0 (.DIODE(net336));
 sky130_fd_sc_hd__diode_2 ANTENNA__2300__S1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2301__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2302__B (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2308__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2309__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__S0 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2310__S1 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2311__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2314__S (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA__2315__A (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2316__C1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__A1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2317__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2318__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2319__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2320__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2321__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2322__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2323__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2324__S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2325__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2327__S (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2329__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2330__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__S0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__2331__S1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__2332__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2333__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__2334__A_N (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__2335__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__2336__A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2337__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2338__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2339__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2340__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2341__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2342__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__S0 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__2343__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2344__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2348__S (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2350__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2351__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2352__S0 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__2353__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__2358__C1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2359__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2360__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2361__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2362__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2363__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2364__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2365__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__2371__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2372__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2373__S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2374__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__2376__A_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2378__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2379__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__A3 (.DIODE(_1568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2380__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2381__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__S0 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2383__S1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__S0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2385__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2386__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2392__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2393__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2394__S0 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2395__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2396__S (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__2399__A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__2400__C1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__2401__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2402__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2403__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2404__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2405__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2406__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2407__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2413__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2414__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2415__S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2416__A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__2418__A_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2420__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2421__C1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2422__C1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2423__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2424__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2425__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2426__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2427__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2428__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__S0 (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__2429__S1 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA__2430__S (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA__2431__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2432__S (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__2433__A_N (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2434__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2435__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2437__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2438__S (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__2439__A_N (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2440__S (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__2441__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2442__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2443__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S0 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA__2444__S1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__S0 (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA__2445__S1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2446__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__S0 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__2447__S1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__S0 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__2448__S1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__2449__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__S0 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__2450__S1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2451__S (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__2452__A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2453__S (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__2454__A_N (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2455__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2456__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__2457__S1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2458__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2460__A_N (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2462__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__2463__C1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__2464__C1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2465__S1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S0 (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__2466__S1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__2467__S1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2468__S1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S0 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__2469__S1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__2470__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__2476__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__2477__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2479__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__2480__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2481__A_N (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2482__S (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2483__A (.DIODE(net281));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__2484__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2485__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__A_N (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__2486__C (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__A_N (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__B (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__C (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__2487__D (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__2488__A_N (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2490__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2491__B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2492__B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2493__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2494__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2495__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2496__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2497__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2498__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2499__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2500__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2501__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2502__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2503__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2504__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2505__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2506__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2507__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2508__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2509__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2510__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2511__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2512__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2513__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2514__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2515__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2516__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2517__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2518__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2519__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2520__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2521__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2522__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__2523__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__A2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__2524__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__2526__B (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2527__C (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2528__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__2529__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2530__B (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2531__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2532__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2533__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2534__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2535__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2536__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2537__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2538__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2539__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2540__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2541__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2542__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2543__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2544__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2545__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2546__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2547__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2548__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2549__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2550__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2551__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2552__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2553__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2554__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2555__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2556__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2557__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2558__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2559__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2560__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__2561__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__2562__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2563__C (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2564__B (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2565__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__2566__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__2567__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2568__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__2569__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2570__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2571__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2572__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2573__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2574__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2575__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2576__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2577__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2578__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2579__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2580__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2581__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2582__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2583__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2584__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2585__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2586__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2587__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2588__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2589__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2590__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2591__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2592__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2593__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2594__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2595__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2596__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2597__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__2598__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__A2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__2599__B1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__A_N (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2600__C (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2601__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__2602__B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__2603__B (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__2604__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__2605__B (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2606__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2608__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2609__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2610__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2611__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2612__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2613__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2614__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2615__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2616__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2617__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2618__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2619__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2620__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2621__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2622__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2623__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2624__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2625__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2626__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2627__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2628__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2629__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2630__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2631__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2632__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2633__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2634__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2635__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__2636__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__A2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__2637__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__A_N (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__B (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__2638__C (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__2640__B (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2641__C (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2642__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2643__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__2644__B (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2645__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2646__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2647__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2648__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2649__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2650__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2651__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2652__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2653__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2654__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2655__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2656__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2657__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2658__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2659__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2660__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2661__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2662__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2663__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2664__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2665__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2666__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2667__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2668__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2669__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2670__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2671__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2672__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2673__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2674__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__A2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__2675__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__A2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__2676__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__2678__B (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__2679__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__2680__B (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2681__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__2682__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2683__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2684__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2685__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2686__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2687__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2688__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2689__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2690__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2691__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2692__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2693__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2694__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2695__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2696__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2697__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2698__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2699__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2700__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2701__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2702__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2703__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2704__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2705__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2706__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2707__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2708__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2709__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2710__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__2711__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__2712__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__2714__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2715__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2716__B (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2717__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2718__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2719__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2720__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2721__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2722__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2723__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2724__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2725__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2726__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2727__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2728__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2729__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2730__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2731__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2732__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2733__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2734__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2735__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2736__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2737__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2738__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2739__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2740__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2741__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2742__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2743__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2744__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2745__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2746__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__A2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__2747__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__A2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__2748__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__2749__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__2750__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2751__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2752__B (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2753__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2754__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2755__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2756__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2757__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2758__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2759__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2760__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2761__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2762__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2763__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2764__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2765__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2766__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2767__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2768__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2769__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2770__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2771__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2772__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2773__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2774__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2775__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2776__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2777__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2778__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2779__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2780__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2781__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2782__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__A2 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__2783__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__2784__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2785__C (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2786__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__2787__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__2788__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__2789__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2790__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2792__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2793__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2794__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2795__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2796__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2797__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2798__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2799__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2800__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2801__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2802__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2803__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2804__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2805__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2806__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2807__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2808__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2809__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2810__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2811__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2811__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2812__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2813__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2814__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2815__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2816__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2817__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2818__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2819__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__A2 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__2820__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__2821__B1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__2822__C (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2823__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__2824__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2825__B (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2826__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2827__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2828__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2829__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2830__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2831__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2832__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2833__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2834__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2835__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2836__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2837__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2838__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2839__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2840__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2841__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2842__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2843__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2843__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2844__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2845__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2846__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2847__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2848__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2849__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2850__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2851__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2852__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2853__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2854__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2854__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2855__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__2856__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__2857__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__2858__B (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2859__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__2860__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2861__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__2861__B (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2862__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2864__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2865__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2866__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2867__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2868__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2869__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2870__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2871__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2872__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2872__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2873__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2874__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2875__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2876__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2877__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2878__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2879__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2880__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2881__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2882__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2883__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2883__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2884__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2885__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2886__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2887__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2888__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2889__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2889__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2890__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2891__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2891__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__A2 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__2892__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__2893__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__2895__B (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__2896__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2897__B (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2898__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2899__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2900__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2901__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2902__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2903__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2904__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2904__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2904__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2905__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2906__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2906__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2907__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2908__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2909__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2910__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2911__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2912__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2913__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2914__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2915__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2916__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2917__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2917__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2918__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2919__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2920__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2921__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2922__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2923__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2924__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2925__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2926__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2927__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__A2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__2928__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__A2 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__2929__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__2931__B (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2932__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__2932__B (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__2933__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2934__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__2935__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2936__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2937__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2938__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__2939__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2940__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2941__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2942__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2943__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2944__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2945__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2946__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2947__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2948__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2949__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2950__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2951__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2952__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2953__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2954__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2955__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2956__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2957__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2958__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2959__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2960__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2961__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2962__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2963__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__2964__B1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__A2 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__2965__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__B (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__2966__C_N (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__2967__B (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2968__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__2969__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__2970__B (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2971__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2973__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2974__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2975__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__2976__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2977__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2978__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2979__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2980__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2981__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2982__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2983__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2984__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2985__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2986__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2987__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2988__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2989__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2990__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2991__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2992__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2993__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2994__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2995__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2996__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2997__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__2998__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__2999__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3000__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3001__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3002__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__3004__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3005__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3006__B (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3007__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3008__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3009__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3010__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3011__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3012__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3013__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3014__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3015__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3016__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3017__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3018__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3019__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3019__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3019__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3020__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3021__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3022__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3023__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3024__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3025__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3026__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3027__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3028__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3029__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3030__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3031__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3032__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3033__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3034__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3035__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3036__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__A2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3037__B1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3038__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__B (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__3039__C_N (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__3040__B (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3041__A (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3042__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3043__B (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3044__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3046__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3046__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3047__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3048__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3049__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3050__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3051__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3052__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3053__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3054__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3055__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3056__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3057__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3058__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3059__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3060__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3061__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3062__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3063__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3064__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3065__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3066__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3067__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3068__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3069__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3070__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3071__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3072__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3073__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__A2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3074__B1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__A2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3075__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__3077__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3078__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3079__B (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3080__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3082__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3083__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3084__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3085__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3086__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3087__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3088__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3089__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3090__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3091__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3092__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3093__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3094__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3095__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3096__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3097__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3098__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3099__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3100__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3101__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3102__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3103__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3104__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3105__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3106__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3107__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3108__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3109__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3110__B1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__A2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3111__B1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__3112__B (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3113__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3114__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3115__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3116__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3117__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3118__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3119__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3120__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3121__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3122__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3123__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3124__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3125__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3126__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3127__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3128__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3129__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3130__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3131__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3132__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3133__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3134__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3135__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3136__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3137__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3138__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3139__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3140__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3141__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3142__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3143__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3144__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3145__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__A2 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3146__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__A2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3147__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__3148__A_N (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__3149__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3150__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3151__B (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3152__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3154__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3155__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3156__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3157__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3158__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3159__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3160__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3161__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3162__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3163__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3164__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3165__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3166__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3167__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3168__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3169__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3170__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3171__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3172__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3173__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3174__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3175__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3176__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3177__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3178__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3179__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3180__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3181__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__A2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3182__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__A2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3183__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__3184__C (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3185__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3186__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3187__B (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3188__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3190__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3191__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3192__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3193__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3194__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3195__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3196__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3197__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3198__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3199__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3200__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3201__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3202__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3203__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3204__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3205__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3206__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3207__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3208__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3209__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3210__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3211__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3212__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3213__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3214__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3215__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3216__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3217__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__3218__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__3219__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__3221__B (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3222__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__3223__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3224__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3225__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3226__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3227__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3228__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3229__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3230__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3231__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3232__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3233__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3234__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3235__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3236__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3237__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3238__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3239__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3240__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3241__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3242__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3243__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3244__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3245__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3246__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3247__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3248__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3249__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3250__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3251__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3252__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3253__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__3254__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__3255__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__3256__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__3257__A (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3258__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3259__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3260__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3262__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3263__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3264__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3265__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3266__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3267__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3268__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3269__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3270__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3271__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3272__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3273__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3274__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3275__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3276__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3277__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3278__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3279__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3280__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3281__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3282__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3283__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3284__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3285__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3286__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3287__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3288__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3289__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__3290__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__3291__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__3292__C (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3293__B (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3294__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3295__B (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3296__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3297__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3298__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3299__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3300__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3301__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3302__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3303__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3304__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3305__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3306__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3307__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3308__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3309__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3310__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3311__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3312__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3313__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3314__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3315__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3316__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3317__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3318__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3319__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3320__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3321__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3322__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3323__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3324__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3325__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__3326__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__3327__B1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3328__B (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3329__A (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3330__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3331__B (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3332__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3334__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3335__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3336__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3337__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3338__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3339__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3340__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3341__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3342__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3343__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3346__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3347__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3348__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3349__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3350__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3352__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3353__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3354__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3356__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3357__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3358__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A_N (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__C (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3365__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__B (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3370__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3372__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3373__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3374__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3376__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3380__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3383__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3384__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3394__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__B1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__3399__B1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3400__B (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3402__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__B (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3411__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3413__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3422__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3423__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3426__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3429__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3432__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3433__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__C (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3437__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__B (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3442__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3446__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3449__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3453__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3454__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__3470__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__3471__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__C (.DIODE(_1693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__B (.DIODE(_1694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__A1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A1 (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3482__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3485__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3486__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A1 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3488__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3492__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3494__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A1 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A1 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3499__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A1 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A1 (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A1 (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3505__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__B1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3508__B (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3510__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3511__B (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3514__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3515__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3517__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3518__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3519__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3523__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3524__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3525__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3526__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3527__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3530__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A2 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__B (.DIODE(_1675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A (.DIODE(_1676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__B (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3548__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3551__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3563__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3566__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3567__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3569__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3577__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__A2 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__A_N (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__B (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__3580__C (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3581__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__B (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3586__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3590__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3594__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3596__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3598__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3601__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3609__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3613__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__A2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3614__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__3615__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3616__C (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3617__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA__3618__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__A (.DIODE(net368));
 sky130_fd_sc_hd__diode_2 ANTENNA__3619__B (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3620__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3622__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__3625__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3627__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3628__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3630__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3631__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3632__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3633__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3634__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A1 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3635__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3636__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3637__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3639__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3640__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3641__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A1 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3643__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3644__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3645__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3646__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3649__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A1 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7__f_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_clk_A (.DIODE(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_clk_A (.DIODE(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(_1748_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(_1806_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(_1699_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(_1682_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(_1669_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(_1026_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(_1025_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout308_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout311_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout315_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout319_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout325_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout343_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout344_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout351_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout352_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout362_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout364_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output61_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire78_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire86_A (.DIODE(net54));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_137_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_157_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_159_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_161_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_163_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_165_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_167_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_171_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_173_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_173_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_173_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_899 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_938 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_964 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _1810_ (.A(net244),
    .Y(_1025_));
 sky130_fd_sc_hd__nand3b_4 _1811_ (.A_N(net41),
    .B(net7),
    .C(net40),
    .Y(_1026_));
 sky130_fd_sc_hd__nor3b_4 _1812_ (.A(net236),
    .B(net243),
    .C_N(net233),
    .Y(_1027_));
 sky130_fd_sc_hd__and3b_2 _1813_ (.A_N(net236),
    .B(net243),
    .C(net233),
    .X(_1028_));
 sky130_fd_sc_hd__mux4_1 _1814_ (.A0(\mem[0][0] ),
    .A1(\mem[1][0] ),
    .A2(\mem[2][0] ),
    .A3(\mem[3][0] ),
    .S0(net340),
    .S1(net292),
    .X(_1029_));
 sky130_fd_sc_hd__mux4_1 _1815_ (.A0(\mem[4][0] ),
    .A1(\mem[5][0] ),
    .A2(\mem[6][0] ),
    .A3(\mem[7][0] ),
    .S0(net341),
    .S1(net292),
    .X(_1030_));
 sky130_fd_sc_hd__mux4_1 _1816_ (.A0(\mem[12][0] ),
    .A1(\mem[13][0] ),
    .A2(\mem[14][0] ),
    .A3(\mem[15][0] ),
    .S0(net340),
    .S1(net292),
    .X(_1031_));
 sky130_fd_sc_hd__mux4_1 _1817_ (.A0(\mem[8][0] ),
    .A1(\mem[9][0] ),
    .A2(\mem[10][0] ),
    .A3(\mem[11][0] ),
    .S0(net340),
    .S1(net292),
    .X(_1032_));
 sky130_fd_sc_hd__mux4_1 _1818_ (.A0(_1029_),
    .A1(_1030_),
    .A2(_1032_),
    .A3(_1031_),
    .S0(net247),
    .S1(net239),
    .X(_1033_));
 sky130_fd_sc_hd__nor2_1 _1819_ (.A(net231),
    .B(_1033_),
    .Y(_1034_));
 sky130_fd_sc_hd__mux4_1 _1820_ (.A0(\mem[24][0] ),
    .A1(\mem[25][0] ),
    .A2(\mem[26][0] ),
    .A3(\mem[27][0] ),
    .S0(net332),
    .S1(net284),
    .X(_1035_));
 sky130_fd_sc_hd__mux2_1 _1821_ (.A0(\mem[30][0] ),
    .A1(\mem[31][0] ),
    .S(net340),
    .X(_1036_));
 sky130_fd_sc_hd__nand2_1 _1822_ (.A(net284),
    .B(_1036_),
    .Y(_1037_));
 sky130_fd_sc_hd__mux2_1 _1823_ (.A0(\mem[28][0] ),
    .A1(\mem[29][0] ),
    .S(net332),
    .X(_1038_));
 sky130_fd_sc_hd__nand2b_1 _1824_ (.A_N(net284),
    .B(_1038_),
    .Y(_1039_));
 sky130_fd_sc_hd__o21ai_1 _1825_ (.A1(net243),
    .A2(_1035_),
    .B1(net236),
    .Y(_1040_));
 sky130_fd_sc_hd__a31o_1 _1826_ (.A1(net247),
    .A2(_1037_),
    .A3(_1039_),
    .B1(_1040_),
    .X(_1041_));
 sky130_fd_sc_hd__mux4_1 _1827_ (.A0(\mem[20][0] ),
    .A1(\mem[21][0] ),
    .A2(\mem[22][0] ),
    .A3(\mem[23][0] ),
    .S0(net331),
    .S1(net283),
    .X(_1042_));
 sky130_fd_sc_hd__nor2_1 _1828_ (.A(net224),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__mux2_1 _1829_ (.A0(\mem[16][0] ),
    .A1(\mem[17][0] ),
    .S(net331),
    .X(_1044_));
 sky130_fd_sc_hd__nand2b_1 _1830_ (.A_N(net283),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__mux2_1 _1831_ (.A0(\mem[18][0] ),
    .A1(\mem[19][0] ),
    .S(net331),
    .X(_1046_));
 sky130_fd_sc_hd__nand2_1 _1832_ (.A(net283),
    .B(_1046_),
    .Y(_1047_));
 sky130_fd_sc_hd__a311o_1 _1833_ (.A1(net224),
    .A2(_1045_),
    .A3(_1047_),
    .B1(_1043_),
    .C1(net236),
    .X(_1048_));
 sky130_fd_sc_hd__a311oi_4 _1834_ (.A1(net231),
    .A2(_1041_),
    .A3(_1048_),
    .B1(net219),
    .C1(_1034_),
    .Y(net43));
 sky130_fd_sc_hd__mux4_1 _1835_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[2][1] ),
    .A3(\mem[3][1] ),
    .S0(net340),
    .S1(net292),
    .X(_1049_));
 sky130_fd_sc_hd__mux4_1 _1836_ (.A0(\mem[4][1] ),
    .A1(\mem[5][1] ),
    .A2(\mem[6][1] ),
    .A3(\mem[7][1] ),
    .S0(net341),
    .S1(net292),
    .X(_1050_));
 sky130_fd_sc_hd__mux4_1 _1837_ (.A0(\mem[12][1] ),
    .A1(\mem[13][1] ),
    .A2(\mem[14][1] ),
    .A3(\mem[15][1] ),
    .S0(net340),
    .S1(net292),
    .X(_1051_));
 sky130_fd_sc_hd__mux4_1 _1838_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[10][1] ),
    .A3(\mem[11][1] ),
    .S0(net340),
    .S1(net292),
    .X(_1052_));
 sky130_fd_sc_hd__mux4_1 _1839_ (.A0(_1049_),
    .A1(_1050_),
    .A2(_1052_),
    .A3(_1051_),
    .S0(net247),
    .S1(net239),
    .X(_1053_));
 sky130_fd_sc_hd__nor2_1 _1840_ (.A(net231),
    .B(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__mux4_1 _1841_ (.A0(\mem[24][1] ),
    .A1(\mem[25][1] ),
    .A2(\mem[26][1] ),
    .A3(\mem[27][1] ),
    .S0(net332),
    .S1(net284),
    .X(_1055_));
 sky130_fd_sc_hd__mux2_1 _1842_ (.A0(\mem[30][1] ),
    .A1(\mem[31][1] ),
    .S(net332),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_1 _1843_ (.A(net284),
    .B(_1056_),
    .Y(_1057_));
 sky130_fd_sc_hd__mux2_1 _1844_ (.A0(\mem[28][1] ),
    .A1(\mem[29][1] ),
    .S(net332),
    .X(_1058_));
 sky130_fd_sc_hd__nand2b_1 _1845_ (.A_N(net284),
    .B(_1058_),
    .Y(_1059_));
 sky130_fd_sc_hd__o21ai_1 _1846_ (.A1(net243),
    .A2(_1055_),
    .B1(net236),
    .Y(_1060_));
 sky130_fd_sc_hd__a31o_1 _1847_ (.A1(net243),
    .A2(_1057_),
    .A3(_1059_),
    .B1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__mux4_1 _1848_ (.A0(\mem[20][1] ),
    .A1(\mem[21][1] ),
    .A2(\mem[22][1] ),
    .A3(\mem[23][1] ),
    .S0(net331),
    .S1(net283),
    .X(_1062_));
 sky130_fd_sc_hd__nor2_1 _1849_ (.A(net224),
    .B(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__mux2_1 _1850_ (.A0(\mem[16][1] ),
    .A1(\mem[17][1] ),
    .S(net331),
    .X(_1064_));
 sky130_fd_sc_hd__nand2b_1 _1851_ (.A_N(net283),
    .B(_1064_),
    .Y(_1065_));
 sky130_fd_sc_hd__mux2_1 _1852_ (.A0(\mem[18][1] ),
    .A1(\mem[19][1] ),
    .S(net331),
    .X(_1066_));
 sky130_fd_sc_hd__nand2_1 _1853_ (.A(net283),
    .B(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__a311o_1 _1854_ (.A1(net224),
    .A2(_1065_),
    .A3(_1067_),
    .B1(_1063_),
    .C1(net236),
    .X(_1068_));
 sky130_fd_sc_hd__a311oi_4 _1855_ (.A1(net231),
    .A2(_1061_),
    .A3(_1068_),
    .B1(net219),
    .C1(_1054_),
    .Y(net54));
 sky130_fd_sc_hd__mux4_1 _1856_ (.A0(\mem[0][2] ),
    .A1(\mem[1][2] ),
    .A2(\mem[2][2] ),
    .A3(\mem[3][2] ),
    .S0(net334),
    .S1(net287),
    .X(_1069_));
 sky130_fd_sc_hd__mux4_1 _1857_ (.A0(\mem[4][2] ),
    .A1(\mem[5][2] ),
    .A2(\mem[6][2] ),
    .A3(\mem[7][2] ),
    .S0(net334),
    .S1(net287),
    .X(_1070_));
 sky130_fd_sc_hd__mux4_1 _1858_ (.A0(\mem[12][2] ),
    .A1(\mem[13][2] ),
    .A2(\mem[14][2] ),
    .A3(\mem[15][2] ),
    .S0(net334),
    .S1(net287),
    .X(_1071_));
 sky130_fd_sc_hd__mux4_1 _1859_ (.A0(\mem[8][2] ),
    .A1(\mem[9][2] ),
    .A2(\mem[10][2] ),
    .A3(\mem[11][2] ),
    .S0(net334),
    .S1(net287),
    .X(_1072_));
 sky130_fd_sc_hd__mux4_1 _1860_ (.A0(_1069_),
    .A1(_1070_),
    .A2(_1072_),
    .A3(_1071_),
    .S0(net245),
    .S1(net238),
    .X(_1073_));
 sky130_fd_sc_hd__nor2_2 _1861_ (.A(net229),
    .B(_1073_),
    .Y(_1074_));
 sky130_fd_sc_hd__mux4_1 _1862_ (.A0(\mem[24][2] ),
    .A1(\mem[25][2] ),
    .A2(\mem[26][2] ),
    .A3(\mem[27][2] ),
    .S0(net318),
    .S1(net270),
    .X(_1075_));
 sky130_fd_sc_hd__mux2_1 _1863_ (.A0(\mem[30][2] ),
    .A1(\mem[31][2] ),
    .S(net318),
    .X(_1076_));
 sky130_fd_sc_hd__nand2_1 _1864_ (.A(net270),
    .B(_1076_),
    .Y(_1077_));
 sky130_fd_sc_hd__mux2_1 _1865_ (.A0(\mem[28][2] ),
    .A1(\mem[29][2] ),
    .S(net318),
    .X(_1078_));
 sky130_fd_sc_hd__nand2b_1 _1866_ (.A_N(net270),
    .B(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__o21ai_1 _1867_ (.A1(net241),
    .A2(_1075_),
    .B1(net234),
    .Y(_1080_));
 sky130_fd_sc_hd__a31o_1 _1868_ (.A1(net241),
    .A2(_1077_),
    .A3(_1079_),
    .B1(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__mux4_1 _1869_ (.A0(\mem[20][2] ),
    .A1(\mem[21][2] ),
    .A2(\mem[22][2] ),
    .A3(\mem[23][2] ),
    .S0(net318),
    .S1(net270),
    .X(_1082_));
 sky130_fd_sc_hd__nor2_1 _1870_ (.A(net220),
    .B(_1082_),
    .Y(_1083_));
 sky130_fd_sc_hd__mux2_1 _1871_ (.A0(\mem[16][2] ),
    .A1(\mem[17][2] ),
    .S(net318),
    .X(_1084_));
 sky130_fd_sc_hd__nand2b_1 _1872_ (.A_N(net270),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__mux2_1 _1873_ (.A0(\mem[18][2] ),
    .A1(\mem[19][2] ),
    .S(net318),
    .X(_1086_));
 sky130_fd_sc_hd__nand2_1 _1874_ (.A(net270),
    .B(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__a311o_1 _1875_ (.A1(net220),
    .A2(_1085_),
    .A3(_1087_),
    .B1(_1083_),
    .C1(net234),
    .X(_1088_));
 sky130_fd_sc_hd__a311oi_4 _1876_ (.A1(net230),
    .A2(_1081_),
    .A3(_1088_),
    .B1(net218),
    .C1(_1074_),
    .Y(net65));
 sky130_fd_sc_hd__mux4_1 _1877_ (.A0(\mem[0][3] ),
    .A1(\mem[1][3] ),
    .A2(\mem[2][3] ),
    .A3(\mem[3][3] ),
    .S0(net339),
    .S1(net291),
    .X(_1089_));
 sky130_fd_sc_hd__mux4_1 _1878_ (.A0(\mem[4][3] ),
    .A1(\mem[5][3] ),
    .A2(\mem[6][3] ),
    .A3(\mem[7][3] ),
    .S0(net339),
    .S1(net291),
    .X(_1090_));
 sky130_fd_sc_hd__mux4_1 _1879_ (.A0(\mem[12][3] ),
    .A1(\mem[13][3] ),
    .A2(\mem[14][3] ),
    .A3(\mem[15][3] ),
    .S0(net339),
    .S1(net291),
    .X(_1091_));
 sky130_fd_sc_hd__mux4_1 _1880_ (.A0(\mem[8][3] ),
    .A1(\mem[9][3] ),
    .A2(\mem[10][3] ),
    .A3(\mem[11][3] ),
    .S0(net339),
    .S1(net291),
    .X(_1092_));
 sky130_fd_sc_hd__mux4_1 _1881_ (.A0(_1089_),
    .A1(_1090_),
    .A2(_1092_),
    .A3(_1091_),
    .S0(net247),
    .S1(net239),
    .X(_1093_));
 sky130_fd_sc_hd__nor2_1 _1882_ (.A(net232),
    .B(_1093_),
    .Y(_1094_));
 sky130_fd_sc_hd__mux4_1 _1883_ (.A0(\mem[24][3] ),
    .A1(\mem[25][3] ),
    .A2(\mem[26][3] ),
    .A3(\mem[27][3] ),
    .S0(net329),
    .S1(net281),
    .X(_1095_));
 sky130_fd_sc_hd__mux2_1 _1884_ (.A0(\mem[30][3] ),
    .A1(\mem[31][3] ),
    .S(net329),
    .X(_1096_));
 sky130_fd_sc_hd__nand2_1 _1885_ (.A(net281),
    .B(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__mux2_1 _1886_ (.A0(\mem[28][3] ),
    .A1(\mem[29][3] ),
    .S(net329),
    .X(_1098_));
 sky130_fd_sc_hd__nand2b_1 _1887_ (.A_N(net281),
    .B(_1098_),
    .Y(_1099_));
 sky130_fd_sc_hd__o21ai_1 _1888_ (.A1(net243),
    .A2(_1095_),
    .B1(net236),
    .Y(_1100_));
 sky130_fd_sc_hd__a31o_1 _1889_ (.A1(net243),
    .A2(_1097_),
    .A3(_1099_),
    .B1(_1100_),
    .X(_1101_));
 sky130_fd_sc_hd__mux4_1 _1890_ (.A0(\mem[20][3] ),
    .A1(\mem[21][3] ),
    .A2(\mem[22][3] ),
    .A3(\mem[23][3] ),
    .S0(net326),
    .S1(net278),
    .X(_1102_));
 sky130_fd_sc_hd__nor2_1 _1891_ (.A(net222),
    .B(_1102_),
    .Y(_1103_));
 sky130_fd_sc_hd__mux2_1 _1892_ (.A0(\mem[16][3] ),
    .A1(\mem[17][3] ),
    .S(net326),
    .X(_1104_));
 sky130_fd_sc_hd__nand2b_1 _1893_ (.A_N(net278),
    .B(_1104_),
    .Y(_1105_));
 sky130_fd_sc_hd__mux2_1 _1894_ (.A0(\mem[18][3] ),
    .A1(\mem[19][3] ),
    .S(net319),
    .X(_1106_));
 sky130_fd_sc_hd__nand2_1 _1895_ (.A(net278),
    .B(_1106_),
    .Y(_1107_));
 sky130_fd_sc_hd__a311o_2 _1896_ (.A1(net222),
    .A2(_1105_),
    .A3(_1107_),
    .B1(_1103_),
    .C1(net234),
    .X(_1108_));
 sky130_fd_sc_hd__a311oi_4 _1897_ (.A1(net232),
    .A2(_1101_),
    .A3(_1108_),
    .B1(_1026_),
    .C1(_1094_),
    .Y(net68));
 sky130_fd_sc_hd__mux4_1 _1898_ (.A0(\mem[0][4] ),
    .A1(\mem[1][4] ),
    .A2(\mem[2][4] ),
    .A3(\mem[3][4] ),
    .S0(net341),
    .S1(net293),
    .X(_1109_));
 sky130_fd_sc_hd__mux4_1 _1899_ (.A0(\mem[4][4] ),
    .A1(\mem[5][4] ),
    .A2(\mem[6][4] ),
    .A3(\mem[7][4] ),
    .S0(net341),
    .S1(net293),
    .X(_1110_));
 sky130_fd_sc_hd__mux4_1 _1900_ (.A0(\mem[12][4] ),
    .A1(\mem[13][4] ),
    .A2(\mem[14][4] ),
    .A3(\mem[15][4] ),
    .S0(net340),
    .S1(net292),
    .X(_1111_));
 sky130_fd_sc_hd__mux4_1 _1901_ (.A0(\mem[8][4] ),
    .A1(\mem[9][4] ),
    .A2(\mem[10][4] ),
    .A3(\mem[11][4] ),
    .S0(net340),
    .S1(net292),
    .X(_1112_));
 sky130_fd_sc_hd__mux4_1 _1902_ (.A0(_1109_),
    .A1(_1110_),
    .A2(_1112_),
    .A3(_1111_),
    .S0(net247),
    .S1(net239),
    .X(_1113_));
 sky130_fd_sc_hd__nor2_1 _1903_ (.A(net231),
    .B(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__mux4_1 _1904_ (.A0(\mem[24][4] ),
    .A1(\mem[25][4] ),
    .A2(\mem[26][4] ),
    .A3(\mem[27][4] ),
    .S0(net332),
    .S1(net284),
    .X(_1115_));
 sky130_fd_sc_hd__mux2_1 _1905_ (.A0(\mem[30][4] ),
    .A1(\mem[31][4] ),
    .S(net340),
    .X(_1116_));
 sky130_fd_sc_hd__nand2_1 _1906_ (.A(net284),
    .B(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__mux2_1 _1907_ (.A0(\mem[28][4] ),
    .A1(\mem[29][4] ),
    .S(net332),
    .X(_1118_));
 sky130_fd_sc_hd__nand2b_1 _1908_ (.A_N(net284),
    .B(_1118_),
    .Y(_1119_));
 sky130_fd_sc_hd__o21ai_1 _1909_ (.A1(net243),
    .A2(_1115_),
    .B1(net236),
    .Y(_1120_));
 sky130_fd_sc_hd__a31o_1 _1910_ (.A1(net247),
    .A2(_1117_),
    .A3(_1119_),
    .B1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__mux4_1 _1911_ (.A0(\mem[20][4] ),
    .A1(\mem[21][4] ),
    .A2(\mem[22][4] ),
    .A3(\mem[23][4] ),
    .S0(net331),
    .S1(net283),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_1 _1912_ (.A(net223),
    .B(_1122_),
    .Y(_1123_));
 sky130_fd_sc_hd__mux2_1 _1913_ (.A0(\mem[16][4] ),
    .A1(\mem[17][4] ),
    .S(net331),
    .X(_1124_));
 sky130_fd_sc_hd__nand2b_1 _1914_ (.A_N(net283),
    .B(_1124_),
    .Y(_1125_));
 sky130_fd_sc_hd__mux2_1 _1915_ (.A0(\mem[18][4] ),
    .A1(\mem[19][4] ),
    .S(net331),
    .X(_1126_));
 sky130_fd_sc_hd__nand2_1 _1916_ (.A(net283),
    .B(_1126_),
    .Y(_1127_));
 sky130_fd_sc_hd__a311o_1 _1917_ (.A1(net223),
    .A2(_1125_),
    .A3(_1127_),
    .B1(_1123_),
    .C1(net237),
    .X(_1128_));
 sky130_fd_sc_hd__a311oi_4 _1918_ (.A1(net231),
    .A2(_1121_),
    .A3(_1128_),
    .B1(net219),
    .C1(_1114_),
    .Y(net69));
 sky130_fd_sc_hd__mux4_1 _1919_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[2][5] ),
    .A3(\mem[3][5] ),
    .S0(net341),
    .S1(net293),
    .X(_1129_));
 sky130_fd_sc_hd__mux4_1 _1920_ (.A0(\mem[4][5] ),
    .A1(\mem[5][5] ),
    .A2(\mem[6][5] ),
    .A3(\mem[7][5] ),
    .S0(net341),
    .S1(net293),
    .X(_1130_));
 sky130_fd_sc_hd__mux4_1 _1921_ (.A0(\mem[12][5] ),
    .A1(\mem[13][5] ),
    .A2(\mem[14][5] ),
    .A3(\mem[15][5] ),
    .S0(net340),
    .S1(net292),
    .X(_1131_));
 sky130_fd_sc_hd__mux4_1 _1922_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[10][5] ),
    .A3(\mem[11][5] ),
    .S0(net340),
    .S1(net292),
    .X(_1132_));
 sky130_fd_sc_hd__mux4_1 _1923_ (.A0(_1129_),
    .A1(_1130_),
    .A2(_1132_),
    .A3(_1131_),
    .S0(net247),
    .S1(net239),
    .X(_1133_));
 sky130_fd_sc_hd__nor2_1 _1924_ (.A(net231),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__mux4_1 _1925_ (.A0(\mem[24][5] ),
    .A1(\mem[25][5] ),
    .A2(\mem[26][5] ),
    .A3(\mem[27][5] ),
    .S0(net332),
    .S1(net284),
    .X(_1135_));
 sky130_fd_sc_hd__mux2_1 _1926_ (.A0(\mem[30][5] ),
    .A1(\mem[31][5] ),
    .S(net332),
    .X(_1136_));
 sky130_fd_sc_hd__nand2_1 _1927_ (.A(net284),
    .B(_1136_),
    .Y(_1137_));
 sky130_fd_sc_hd__mux2_1 _1928_ (.A0(\mem[28][5] ),
    .A1(\mem[29][5] ),
    .S(net332),
    .X(_1138_));
 sky130_fd_sc_hd__nand2b_1 _1929_ (.A_N(net284),
    .B(_1138_),
    .Y(_1139_));
 sky130_fd_sc_hd__o21ai_1 _1930_ (.A1(net244),
    .A2(_1135_),
    .B1(net237),
    .Y(_1140_));
 sky130_fd_sc_hd__a31o_1 _1931_ (.A1(net244),
    .A2(_1137_),
    .A3(_1139_),
    .B1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__mux4_1 _1932_ (.A0(\mem[20][5] ),
    .A1(\mem[21][5] ),
    .A2(\mem[22][5] ),
    .A3(\mem[23][5] ),
    .S0(net331),
    .S1(net283),
    .X(_1142_));
 sky130_fd_sc_hd__nor2_1 _1933_ (.A(net223),
    .B(_1142_),
    .Y(_1143_));
 sky130_fd_sc_hd__mux2_1 _1934_ (.A0(\mem[16][5] ),
    .A1(\mem[17][5] ),
    .S(net331),
    .X(_1144_));
 sky130_fd_sc_hd__nand2b_1 _1935_ (.A_N(net283),
    .B(_1144_),
    .Y(_1145_));
 sky130_fd_sc_hd__mux2_1 _1936_ (.A0(\mem[18][5] ),
    .A1(\mem[19][5] ),
    .S(net332),
    .X(_1146_));
 sky130_fd_sc_hd__nand2_1 _1937_ (.A(net283),
    .B(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__a311o_1 _1938_ (.A1(net224),
    .A2(_1145_),
    .A3(_1147_),
    .B1(_1143_),
    .C1(net237),
    .X(_1148_));
 sky130_fd_sc_hd__a311oi_4 _1939_ (.A1(net231),
    .A2(_1141_),
    .A3(_1148_),
    .B1(net219),
    .C1(_1134_),
    .Y(net70));
 sky130_fd_sc_hd__mux4_1 _1940_ (.A0(\mem[0][6] ),
    .A1(\mem[1][6] ),
    .A2(\mem[2][6] ),
    .A3(\mem[3][6] ),
    .S0(net343),
    .S1(net295),
    .X(_1149_));
 sky130_fd_sc_hd__mux4_1 _1941_ (.A0(\mem[4][6] ),
    .A1(\mem[5][6] ),
    .A2(\mem[6][6] ),
    .A3(\mem[7][6] ),
    .S0(net344),
    .S1(net296),
    .X(_1150_));
 sky130_fd_sc_hd__mux4_1 _1942_ (.A0(\mem[12][6] ),
    .A1(\mem[13][6] ),
    .A2(\mem[14][6] ),
    .A3(\mem[15][6] ),
    .S0(net343),
    .S1(net295),
    .X(_1151_));
 sky130_fd_sc_hd__mux4_1 _1943_ (.A0(\mem[8][6] ),
    .A1(\mem[9][6] ),
    .A2(\mem[10][6] ),
    .A3(\mem[11][6] ),
    .S0(net343),
    .S1(net295),
    .X(_1152_));
 sky130_fd_sc_hd__mux4_2 _1944_ (.A0(_1149_),
    .A1(_1150_),
    .A2(_1152_),
    .A3(_1151_),
    .S0(net247),
    .S1(net239),
    .X(_1153_));
 sky130_fd_sc_hd__nor2_2 _1945_ (.A(net231),
    .B(_1153_),
    .Y(_1154_));
 sky130_fd_sc_hd__mux4_1 _1946_ (.A0(\mem[24][6] ),
    .A1(\mem[25][6] ),
    .A2(\mem[26][6] ),
    .A3(\mem[27][6] ),
    .S0(net330),
    .S1(net281),
    .X(_1155_));
 sky130_fd_sc_hd__mux2_1 _1947_ (.A0(\mem[30][6] ),
    .A1(\mem[31][6] ),
    .S(net331),
    .X(_1156_));
 sky130_fd_sc_hd__nand2_1 _1948_ (.A(net280),
    .B(_1156_),
    .Y(_1157_));
 sky130_fd_sc_hd__mux2_1 _1949_ (.A0(\mem[28][6] ),
    .A1(\mem[29][6] ),
    .S(net328),
    .X(_1158_));
 sky130_fd_sc_hd__nand2b_1 _1950_ (.A_N(net280),
    .B(_1158_),
    .Y(_1159_));
 sky130_fd_sc_hd__o21ai_1 _1951_ (.A1(net243),
    .A2(_1155_),
    .B1(net236),
    .Y(_1160_));
 sky130_fd_sc_hd__a31o_1 _1952_ (.A1(net244),
    .A2(_1157_),
    .A3(_1159_),
    .B1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__mux4_1 _1953_ (.A0(\mem[20][6] ),
    .A1(\mem[21][6] ),
    .A2(\mem[22][6] ),
    .A3(\mem[23][6] ),
    .S0(net328),
    .S1(net280),
    .X(_1162_));
 sky130_fd_sc_hd__nor2_1 _1954_ (.A(net223),
    .B(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__mux2_1 _1955_ (.A0(\mem[16][6] ),
    .A1(\mem[17][6] ),
    .S(net326),
    .X(_1164_));
 sky130_fd_sc_hd__nand2b_1 _1956_ (.A_N(net278),
    .B(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__mux2_1 _1957_ (.A0(\mem[18][6] ),
    .A1(\mem[19][6] ),
    .S(net328),
    .X(_1166_));
 sky130_fd_sc_hd__nand2_1 _1958_ (.A(net280),
    .B(_1166_),
    .Y(_1167_));
 sky130_fd_sc_hd__a311o_1 _1959_ (.A1(net223),
    .A2(_1165_),
    .A3(_1167_),
    .B1(_1163_),
    .C1(net237),
    .X(_1168_));
 sky130_fd_sc_hd__a311oi_4 _1960_ (.A1(net233),
    .A2(_1161_),
    .A3(_1168_),
    .B1(net219),
    .C1(_1154_),
    .Y(net71));
 sky130_fd_sc_hd__mux4_1 _1961_ (.A0(\mem[0][7] ),
    .A1(\mem[1][7] ),
    .A2(\mem[2][7] ),
    .A3(\mem[3][7] ),
    .S0(net336),
    .S1(net288),
    .X(_1169_));
 sky130_fd_sc_hd__mux4_1 _1962_ (.A0(\mem[4][7] ),
    .A1(\mem[5][7] ),
    .A2(\mem[6][7] ),
    .A3(\mem[7][7] ),
    .S0(net337),
    .S1(net289),
    .X(_1170_));
 sky130_fd_sc_hd__mux4_1 _1963_ (.A0(\mem[12][7] ),
    .A1(\mem[13][7] ),
    .A2(\mem[14][7] ),
    .A3(\mem[15][7] ),
    .S0(net337),
    .S1(net289),
    .X(_1171_));
 sky130_fd_sc_hd__mux4_1 _1964_ (.A0(\mem[8][7] ),
    .A1(\mem[9][7] ),
    .A2(\mem[10][7] ),
    .A3(\mem[11][7] ),
    .S0(net337),
    .S1(net289),
    .X(_1172_));
 sky130_fd_sc_hd__mux4_2 _1965_ (.A0(_1169_),
    .A1(_1170_),
    .A2(_1172_),
    .A3(_1171_),
    .S0(net245),
    .S1(net238),
    .X(_1173_));
 sky130_fd_sc_hd__nor2_1 _1966_ (.A(net230),
    .B(_1173_),
    .Y(_1174_));
 sky130_fd_sc_hd__mux4_1 _1967_ (.A0(\mem[24][7] ),
    .A1(\mem[25][7] ),
    .A2(\mem[26][7] ),
    .A3(\mem[27][7] ),
    .S0(net318),
    .S1(net270),
    .X(_1175_));
 sky130_fd_sc_hd__mux2_1 _1968_ (.A0(\mem[30][7] ),
    .A1(\mem[31][7] ),
    .S(net318),
    .X(_1176_));
 sky130_fd_sc_hd__nand2_1 _1969_ (.A(net270),
    .B(_1176_),
    .Y(_1177_));
 sky130_fd_sc_hd__mux2_1 _1970_ (.A0(\mem[28][7] ),
    .A1(\mem[29][7] ),
    .S(net318),
    .X(_1178_));
 sky130_fd_sc_hd__nand2b_1 _1971_ (.A_N(net270),
    .B(_1178_),
    .Y(_1179_));
 sky130_fd_sc_hd__o21ai_1 _1972_ (.A1(net241),
    .A2(_1175_),
    .B1(net234),
    .Y(_1180_));
 sky130_fd_sc_hd__a31o_1 _1973_ (.A1(net241),
    .A2(_1177_),
    .A3(_1179_),
    .B1(_1180_),
    .X(_1181_));
 sky130_fd_sc_hd__mux4_1 _1974_ (.A0(\mem[20][7] ),
    .A1(\mem[21][7] ),
    .A2(\mem[22][7] ),
    .A3(\mem[23][7] ),
    .S0(net319),
    .S1(net271),
    .X(_1182_));
 sky130_fd_sc_hd__nor2_1 _1975_ (.A(net220),
    .B(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__mux2_1 _1976_ (.A0(\mem[16][7] ),
    .A1(\mem[17][7] ),
    .S(net318),
    .X(_1184_));
 sky130_fd_sc_hd__nand2b_1 _1977_ (.A_N(net270),
    .B(_1184_),
    .Y(_1185_));
 sky130_fd_sc_hd__mux2_1 _1978_ (.A0(\mem[18][7] ),
    .A1(\mem[19][7] ),
    .S(net319),
    .X(_1186_));
 sky130_fd_sc_hd__nand2_1 _1979_ (.A(net270),
    .B(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__a311o_1 _1980_ (.A1(net220),
    .A2(_1185_),
    .A3(_1187_),
    .B1(_1183_),
    .C1(net234),
    .X(_1188_));
 sky130_fd_sc_hd__a311oi_2 _1981_ (.A1(net230),
    .A2(_1181_),
    .A3(_1188_),
    .B1(net218),
    .C1(_1174_),
    .Y(net72));
 sky130_fd_sc_hd__mux4_1 _1982_ (.A0(\mem[0][8] ),
    .A1(\mem[1][8] ),
    .A2(\mem[2][8] ),
    .A3(\mem[3][8] ),
    .S0(net336),
    .S1(net288),
    .X(_1189_));
 sky130_fd_sc_hd__mux4_1 _1983_ (.A0(\mem[4][8] ),
    .A1(\mem[5][8] ),
    .A2(\mem[6][8] ),
    .A3(\mem[7][8] ),
    .S0(net335),
    .S1(net286),
    .X(_1190_));
 sky130_fd_sc_hd__mux4_1 _1984_ (.A0(\mem[12][8] ),
    .A1(\mem[13][8] ),
    .A2(\mem[14][8] ),
    .A3(\mem[15][8] ),
    .S0(net335),
    .S1(net286),
    .X(_1191_));
 sky130_fd_sc_hd__mux4_1 _1985_ (.A0(\mem[8][8] ),
    .A1(\mem[9][8] ),
    .A2(\mem[10][8] ),
    .A3(\mem[11][8] ),
    .S0(net335),
    .S1(net286),
    .X(_1192_));
 sky130_fd_sc_hd__mux4_1 _1986_ (.A0(_1189_),
    .A1(_1190_),
    .A2(_1192_),
    .A3(_1191_),
    .S0(net245),
    .S1(net238),
    .X(_1193_));
 sky130_fd_sc_hd__nor2_1 _1987_ (.A(net229),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__mux4_1 _1988_ (.A0(\mem[24][8] ),
    .A1(\mem[25][8] ),
    .A2(\mem[26][8] ),
    .A3(\mem[27][8] ),
    .S0(net324),
    .S1(net276),
    .X(_1195_));
 sky130_fd_sc_hd__mux2_1 _1989_ (.A0(\mem[30][8] ),
    .A1(\mem[31][8] ),
    .S(net324),
    .X(_1196_));
 sky130_fd_sc_hd__nand2_1 _1990_ (.A(net276),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__mux2_1 _1991_ (.A0(\mem[28][8] ),
    .A1(\mem[29][8] ),
    .S(net335),
    .X(_1198_));
 sky130_fd_sc_hd__nand2b_1 _1992_ (.A_N(net276),
    .B(_1198_),
    .Y(_1199_));
 sky130_fd_sc_hd__o21ai_1 _1993_ (.A1(net242),
    .A2(_1195_),
    .B1(net235),
    .Y(_1200_));
 sky130_fd_sc_hd__a31o_1 _1994_ (.A1(net245),
    .A2(_1197_),
    .A3(_1199_),
    .B1(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__mux4_1 _1995_ (.A0(\mem[20][8] ),
    .A1(\mem[21][8] ),
    .A2(\mem[22][8] ),
    .A3(\mem[23][8] ),
    .S0(net324),
    .S1(net276),
    .X(_1202_));
 sky130_fd_sc_hd__nor2_1 _1996_ (.A(net221),
    .B(_1202_),
    .Y(_1203_));
 sky130_fd_sc_hd__mux2_1 _1997_ (.A0(\mem[16][8] ),
    .A1(\mem[17][8] ),
    .S(net324),
    .X(_1204_));
 sky130_fd_sc_hd__nand2b_1 _1998_ (.A_N(net276),
    .B(_1204_),
    .Y(_1205_));
 sky130_fd_sc_hd__mux2_1 _1999_ (.A0(\mem[18][8] ),
    .A1(\mem[19][8] ),
    .S(net330),
    .X(_1206_));
 sky130_fd_sc_hd__nand2_1 _2000_ (.A(net276),
    .B(_1206_),
    .Y(_1207_));
 sky130_fd_sc_hd__a311o_1 _2001_ (.A1(net221),
    .A2(_1205_),
    .A3(_1207_),
    .B1(_1203_),
    .C1(net235),
    .X(_1208_));
 sky130_fd_sc_hd__a311oi_4 _2002_ (.A1(net229),
    .A2(_1201_),
    .A3(_1208_),
    .B1(net218),
    .C1(_1194_),
    .Y(net73));
 sky130_fd_sc_hd__mux4_1 _2003_ (.A0(\mem[0][9] ),
    .A1(\mem[1][9] ),
    .A2(\mem[2][9] ),
    .A3(\mem[3][9] ),
    .S0(net337),
    .S1(net289),
    .X(_1209_));
 sky130_fd_sc_hd__mux4_1 _2004_ (.A0(\mem[4][9] ),
    .A1(\mem[5][9] ),
    .A2(\mem[6][9] ),
    .A3(\mem[7][9] ),
    .S0(net337),
    .S1(net289),
    .X(_1210_));
 sky130_fd_sc_hd__mux4_1 _2005_ (.A0(\mem[12][9] ),
    .A1(\mem[13][9] ),
    .A2(\mem[14][9] ),
    .A3(\mem[15][9] ),
    .S0(net337),
    .S1(net289),
    .X(_1211_));
 sky130_fd_sc_hd__mux4_1 _2006_ (.A0(\mem[8][9] ),
    .A1(\mem[9][9] ),
    .A2(\mem[10][9] ),
    .A3(\mem[11][9] ),
    .S0(net337),
    .S1(net289),
    .X(_1212_));
 sky130_fd_sc_hd__mux4_2 _2007_ (.A0(_1209_),
    .A1(_1210_),
    .A2(_1212_),
    .A3(_1211_),
    .S0(net245),
    .S1(net238),
    .X(_1213_));
 sky130_fd_sc_hd__nor2_1 _2008_ (.A(net230),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__mux4_1 _2009_ (.A0(\mem[24][9] ),
    .A1(\mem[25][9] ),
    .A2(\mem[26][9] ),
    .A3(\mem[27][9] ),
    .S0(net322),
    .S1(net274),
    .X(_1215_));
 sky130_fd_sc_hd__mux2_1 _2010_ (.A0(\mem[30][9] ),
    .A1(\mem[31][9] ),
    .S(net322),
    .X(_1216_));
 sky130_fd_sc_hd__nand2_1 _2011_ (.A(net274),
    .B(_1216_),
    .Y(_1217_));
 sky130_fd_sc_hd__mux2_1 _2012_ (.A0(\mem[28][9] ),
    .A1(\mem[29][9] ),
    .S(net322),
    .X(_1218_));
 sky130_fd_sc_hd__nand2b_1 _2013_ (.A_N(net274),
    .B(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__o21ai_1 _2014_ (.A1(net242),
    .A2(_1215_),
    .B1(net235),
    .Y(_1220_));
 sky130_fd_sc_hd__a31o_1 _2015_ (.A1(net242),
    .A2(_1217_),
    .A3(_1219_),
    .B1(_1220_),
    .X(_1221_));
 sky130_fd_sc_hd__mux4_1 _2016_ (.A0(\mem[20][9] ),
    .A1(\mem[21][9] ),
    .A2(\mem[22][9] ),
    .A3(\mem[23][9] ),
    .S0(net318),
    .S1(net270),
    .X(_1222_));
 sky130_fd_sc_hd__nor2_1 _2017_ (.A(net221),
    .B(_1222_),
    .Y(_1223_));
 sky130_fd_sc_hd__mux2_1 _2018_ (.A0(\mem[16][9] ),
    .A1(\mem[17][9] ),
    .S(net322),
    .X(_1224_));
 sky130_fd_sc_hd__nand2b_1 _2019_ (.A_N(net274),
    .B(_1224_),
    .Y(_1225_));
 sky130_fd_sc_hd__mux2_1 _2020_ (.A0(\mem[18][9] ),
    .A1(\mem[19][9] ),
    .S(net322),
    .X(_1226_));
 sky130_fd_sc_hd__nand2_1 _2021_ (.A(net274),
    .B(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__a311o_1 _2022_ (.A1(net221),
    .A2(_1225_),
    .A3(_1227_),
    .B1(_1223_),
    .C1(net234),
    .X(_1228_));
 sky130_fd_sc_hd__a311oi_4 _2023_ (.A1(net230),
    .A2(_1221_),
    .A3(_1228_),
    .B1(net218),
    .C1(_1214_),
    .Y(net74));
 sky130_fd_sc_hd__mux4_1 _2024_ (.A0(\mem[0][10] ),
    .A1(\mem[1][10] ),
    .A2(\mem[2][10] ),
    .A3(\mem[3][10] ),
    .S0(net343),
    .S1(net295),
    .X(_1229_));
 sky130_fd_sc_hd__mux4_1 _2025_ (.A0(\mem[4][10] ),
    .A1(\mem[5][10] ),
    .A2(\mem[6][10] ),
    .A3(\mem[7][10] ),
    .S0(net343),
    .S1(net295),
    .X(_1230_));
 sky130_fd_sc_hd__mux4_1 _2026_ (.A0(\mem[12][10] ),
    .A1(\mem[13][10] ),
    .A2(\mem[14][10] ),
    .A3(\mem[15][10] ),
    .S0(net343),
    .S1(net295),
    .X(_1231_));
 sky130_fd_sc_hd__mux4_1 _2027_ (.A0(\mem[8][10] ),
    .A1(\mem[9][10] ),
    .A2(\mem[10][10] ),
    .A3(\mem[11][10] ),
    .S0(net343),
    .S1(net295),
    .X(_1232_));
 sky130_fd_sc_hd__mux4_2 _2028_ (.A0(_1229_),
    .A1(_1230_),
    .A2(_1232_),
    .A3(_1231_),
    .S0(net247),
    .S1(net238),
    .X(_1233_));
 sky130_fd_sc_hd__nor2_1 _2029_ (.A(net230),
    .B(_1233_),
    .Y(_1234_));
 sky130_fd_sc_hd__mux4_1 _2030_ (.A0(\mem[24][10] ),
    .A1(\mem[25][10] ),
    .A2(\mem[26][10] ),
    .A3(\mem[27][10] ),
    .S0(net326),
    .S1(net279),
    .X(_1235_));
 sky130_fd_sc_hd__mux2_1 _2031_ (.A0(\mem[30][10] ),
    .A1(\mem[31][10] ),
    .S(net320),
    .X(_1236_));
 sky130_fd_sc_hd__nand2_1 _2032_ (.A(net271),
    .B(_1236_),
    .Y(_1237_));
 sky130_fd_sc_hd__mux2_1 _2033_ (.A0(\mem[28][10] ),
    .A1(\mem[29][10] ),
    .S(net320),
    .X(_1238_));
 sky130_fd_sc_hd__nand2b_1 _2034_ (.A_N(net272),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__o21ai_1 _2035_ (.A1(net241),
    .A2(_1235_),
    .B1(net234),
    .Y(_1240_));
 sky130_fd_sc_hd__a31o_1 _2036_ (.A1(net241),
    .A2(_1237_),
    .A3(_1239_),
    .B1(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__mux4_1 _2037_ (.A0(\mem[20][10] ),
    .A1(\mem[21][10] ),
    .A2(\mem[22][10] ),
    .A3(\mem[23][10] ),
    .S0(net326),
    .S1(net278),
    .X(_1242_));
 sky130_fd_sc_hd__nor2_1 _2038_ (.A(net220),
    .B(_1242_),
    .Y(_1243_));
 sky130_fd_sc_hd__mux2_1 _2039_ (.A0(\mem[16][10] ),
    .A1(\mem[17][10] ),
    .S(net320),
    .X(_1244_));
 sky130_fd_sc_hd__nand2b_1 _2040_ (.A_N(net271),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__mux2_1 _2041_ (.A0(\mem[18][10] ),
    .A1(\mem[19][10] ),
    .S(net319),
    .X(_1246_));
 sky130_fd_sc_hd__nand2_1 _2042_ (.A(net271),
    .B(_1246_),
    .Y(_1247_));
 sky130_fd_sc_hd__a311o_1 _2043_ (.A1(net220),
    .A2(_1245_),
    .A3(_1247_),
    .B1(_1243_),
    .C1(net234),
    .X(_1248_));
 sky130_fd_sc_hd__a311oi_1 _2044_ (.A1(net230),
    .A2(_1241_),
    .A3(_1248_),
    .B1(net218),
    .C1(_1234_),
    .Y(net44));
 sky130_fd_sc_hd__mux4_1 _2045_ (.A0(\mem[0][11] ),
    .A1(\mem[1][11] ),
    .A2(\mem[2][11] ),
    .A3(\mem[3][11] ),
    .S0(net337),
    .S1(net289),
    .X(_1249_));
 sky130_fd_sc_hd__mux4_1 _2046_ (.A0(\mem[4][11] ),
    .A1(\mem[5][11] ),
    .A2(\mem[6][11] ),
    .A3(\mem[7][11] ),
    .S0(net337),
    .S1(net289),
    .X(_1250_));
 sky130_fd_sc_hd__mux4_1 _2047_ (.A0(\mem[12][11] ),
    .A1(\mem[13][11] ),
    .A2(\mem[14][11] ),
    .A3(\mem[15][11] ),
    .S0(net337),
    .S1(net289),
    .X(_1251_));
 sky130_fd_sc_hd__mux4_1 _2048_ (.A0(\mem[8][11] ),
    .A1(\mem[9][11] ),
    .A2(\mem[10][11] ),
    .A3(\mem[11][11] ),
    .S0(net337),
    .S1(net289),
    .X(_1252_));
 sky130_fd_sc_hd__mux4_2 _2049_ (.A0(_1249_),
    .A1(_1250_),
    .A2(_1252_),
    .A3(_1251_),
    .S0(net246),
    .S1(net238),
    .X(_1253_));
 sky130_fd_sc_hd__nor2_1 _2050_ (.A(net229),
    .B(_1253_),
    .Y(_1254_));
 sky130_fd_sc_hd__mux4_1 _2051_ (.A0(\mem[24][11] ),
    .A1(\mem[25][11] ),
    .A2(\mem[26][11] ),
    .A3(\mem[27][11] ),
    .S0(net322),
    .S1(net275),
    .X(_1255_));
 sky130_fd_sc_hd__mux2_1 _2052_ (.A0(\mem[30][11] ),
    .A1(\mem[31][11] ),
    .S(net322),
    .X(_1256_));
 sky130_fd_sc_hd__nand2_1 _2053_ (.A(net275),
    .B(_1256_),
    .Y(_1257_));
 sky130_fd_sc_hd__mux2_1 _2054_ (.A0(\mem[28][11] ),
    .A1(\mem[29][11] ),
    .S(net322),
    .X(_1258_));
 sky130_fd_sc_hd__nand2b_1 _2055_ (.A_N(net275),
    .B(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__o21ai_1 _2056_ (.A1(net242),
    .A2(_1255_),
    .B1(net235),
    .Y(_1260_));
 sky130_fd_sc_hd__a31o_1 _2057_ (.A1(net242),
    .A2(_1257_),
    .A3(_1259_),
    .B1(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__mux4_1 _2058_ (.A0(\mem[20][11] ),
    .A1(\mem[21][11] ),
    .A2(\mem[22][11] ),
    .A3(\mem[23][11] ),
    .S0(net324),
    .S1(net276),
    .X(_1262_));
 sky130_fd_sc_hd__nor2_1 _2059_ (.A(net221),
    .B(_1262_),
    .Y(_1263_));
 sky130_fd_sc_hd__mux2_1 _2060_ (.A0(\mem[16][11] ),
    .A1(\mem[17][11] ),
    .S(net323),
    .X(_1264_));
 sky130_fd_sc_hd__nand2b_1 _2061_ (.A_N(net274),
    .B(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__mux2_1 _2062_ (.A0(\mem[18][11] ),
    .A1(\mem[19][11] ),
    .S(net322),
    .X(_1266_));
 sky130_fd_sc_hd__nand2_1 _2063_ (.A(net274),
    .B(_1266_),
    .Y(_1267_));
 sky130_fd_sc_hd__a311o_1 _2064_ (.A1(net221),
    .A2(_1265_),
    .A3(_1267_),
    .B1(_1263_),
    .C1(net235),
    .X(_1268_));
 sky130_fd_sc_hd__a311oi_4 _2065_ (.A1(net229),
    .A2(_1261_),
    .A3(_1268_),
    .B1(net218),
    .C1(_1254_),
    .Y(net45));
 sky130_fd_sc_hd__mux4_1 _2066_ (.A0(\mem[0][12] ),
    .A1(\mem[1][12] ),
    .A2(\mem[2][12] ),
    .A3(\mem[3][12] ),
    .S0(net339),
    .S1(net291),
    .X(_1269_));
 sky130_fd_sc_hd__mux4_1 _2067_ (.A0(\mem[4][12] ),
    .A1(\mem[5][12] ),
    .A2(\mem[6][12] ),
    .A3(\mem[7][12] ),
    .S0(net339),
    .S1(net291),
    .X(_1270_));
 sky130_fd_sc_hd__mux4_1 _2068_ (.A0(\mem[12][12] ),
    .A1(\mem[13][12] ),
    .A2(\mem[14][12] ),
    .A3(\mem[15][12] ),
    .S0(net339),
    .S1(net291),
    .X(_1271_));
 sky130_fd_sc_hd__mux4_1 _2069_ (.A0(\mem[8][12] ),
    .A1(\mem[9][12] ),
    .A2(\mem[10][12] ),
    .A3(\mem[11][12] ),
    .S0(net339),
    .S1(net291),
    .X(_1272_));
 sky130_fd_sc_hd__mux4_1 _2070_ (.A0(_1269_),
    .A1(_1270_),
    .A2(_1272_),
    .A3(_1271_),
    .S0(net247),
    .S1(net239),
    .X(_1273_));
 sky130_fd_sc_hd__nor2_2 _2071_ (.A(net232),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__mux4_1 _2072_ (.A0(\mem[24][12] ),
    .A1(\mem[25][12] ),
    .A2(\mem[26][12] ),
    .A3(\mem[27][12] ),
    .S0(net327),
    .S1(net279),
    .X(_1275_));
 sky130_fd_sc_hd__mux2_1 _2073_ (.A0(\mem[30][12] ),
    .A1(\mem[31][12] ),
    .S(net330),
    .X(_1276_));
 sky130_fd_sc_hd__nand2_1 _2074_ (.A(net279),
    .B(_1276_),
    .Y(_1277_));
 sky130_fd_sc_hd__mux2_1 _2075_ (.A0(\mem[28][12] ),
    .A1(\mem[29][12] ),
    .S(net327),
    .X(_1278_));
 sky130_fd_sc_hd__nand2b_1 _2076_ (.A_N(net279),
    .B(_1278_),
    .Y(_1279_));
 sky130_fd_sc_hd__o21ai_1 _2077_ (.A1(net244),
    .A2(_1275_),
    .B1(net237),
    .Y(_1280_));
 sky130_fd_sc_hd__a31o_1 _2078_ (.A1(net244),
    .A2(_1277_),
    .A3(_1279_),
    .B1(_1280_),
    .X(_1281_));
 sky130_fd_sc_hd__mux4_1 _2079_ (.A0(\mem[20][12] ),
    .A1(\mem[21][12] ),
    .A2(\mem[22][12] ),
    .A3(\mem[23][12] ),
    .S0(net326),
    .S1(net278),
    .X(_1282_));
 sky130_fd_sc_hd__nor2_1 _2080_ (.A(net223),
    .B(_1282_),
    .Y(_1283_));
 sky130_fd_sc_hd__mux2_1 _2081_ (.A0(\mem[16][12] ),
    .A1(\mem[17][12] ),
    .S(net326),
    .X(_1284_));
 sky130_fd_sc_hd__nand2b_1 _2082_ (.A_N(net278),
    .B(_1284_),
    .Y(_1285_));
 sky130_fd_sc_hd__mux2_1 _2083_ (.A0(\mem[18][12] ),
    .A1(\mem[19][12] ),
    .S(net326),
    .X(_1286_));
 sky130_fd_sc_hd__nand2_1 _2084_ (.A(net278),
    .B(_1286_),
    .Y(_1287_));
 sky130_fd_sc_hd__a311o_2 _2085_ (.A1(net223),
    .A2(_1285_),
    .A3(_1287_),
    .B1(_1283_),
    .C1(net237),
    .X(_1288_));
 sky130_fd_sc_hd__a311oi_4 _2086_ (.A1(net233),
    .A2(_1281_),
    .A3(_1288_),
    .B1(net219),
    .C1(_1274_),
    .Y(net46));
 sky130_fd_sc_hd__mux4_1 _2087_ (.A0(\mem[0][13] ),
    .A1(\mem[1][13] ),
    .A2(\mem[2][13] ),
    .A3(\mem[3][13] ),
    .S0(net336),
    .S1(net288),
    .X(_1289_));
 sky130_fd_sc_hd__mux4_1 _2088_ (.A0(\mem[4][13] ),
    .A1(\mem[5][13] ),
    .A2(\mem[6][13] ),
    .A3(\mem[7][13] ),
    .S0(net336),
    .S1(net288),
    .X(_1290_));
 sky130_fd_sc_hd__mux4_1 _2089_ (.A0(\mem[12][13] ),
    .A1(\mem[13][13] ),
    .A2(\mem[14][13] ),
    .A3(\mem[15][13] ),
    .S0(net336),
    .S1(net288),
    .X(_1291_));
 sky130_fd_sc_hd__mux4_1 _2090_ (.A0(\mem[8][13] ),
    .A1(\mem[9][13] ),
    .A2(\mem[10][13] ),
    .A3(\mem[11][13] ),
    .S0(net336),
    .S1(net288),
    .X(_1292_));
 sky130_fd_sc_hd__mux4_2 _2091_ (.A0(_1289_),
    .A1(_1290_),
    .A2(_1292_),
    .A3(_1291_),
    .S0(net246),
    .S1(net238),
    .X(_1293_));
 sky130_fd_sc_hd__nor2_1 _2092_ (.A(net229),
    .B(_1293_),
    .Y(_1294_));
 sky130_fd_sc_hd__mux4_1 _2093_ (.A0(\mem[24][13] ),
    .A1(\mem[25][13] ),
    .A2(\mem[26][13] ),
    .A3(\mem[27][13] ),
    .S0(net325),
    .S1(net276),
    .X(_1295_));
 sky130_fd_sc_hd__mux2_1 _2094_ (.A0(\mem[30][13] ),
    .A1(\mem[31][13] ),
    .S(net325),
    .X(_1296_));
 sky130_fd_sc_hd__nand2_1 _2095_ (.A(net277),
    .B(_1296_),
    .Y(_1297_));
 sky130_fd_sc_hd__mux2_1 _2096_ (.A0(\mem[28][13] ),
    .A1(\mem[29][13] ),
    .S(net325),
    .X(_1298_));
 sky130_fd_sc_hd__nand2b_1 _2097_ (.A_N(net277),
    .B(_1298_),
    .Y(_1299_));
 sky130_fd_sc_hd__o21ai_1 _2098_ (.A1(net242),
    .A2(_1295_),
    .B1(net235),
    .Y(_1300_));
 sky130_fd_sc_hd__a31o_1 _2099_ (.A1(net245),
    .A2(_1297_),
    .A3(_1299_),
    .B1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__mux4_1 _2100_ (.A0(\mem[20][13] ),
    .A1(\mem[21][13] ),
    .A2(\mem[22][13] ),
    .A3(\mem[23][13] ),
    .S0(net324),
    .S1(net276),
    .X(_1302_));
 sky130_fd_sc_hd__nor2_1 _2101_ (.A(net222),
    .B(_1302_),
    .Y(_1303_));
 sky130_fd_sc_hd__mux2_1 _2102_ (.A0(\mem[16][13] ),
    .A1(\mem[17][13] ),
    .S(net325),
    .X(_1304_));
 sky130_fd_sc_hd__nand2b_1 _2103_ (.A_N(net276),
    .B(_1304_),
    .Y(_1305_));
 sky130_fd_sc_hd__mux2_1 _2104_ (.A0(\mem[18][13] ),
    .A1(\mem[19][13] ),
    .S(net324),
    .X(_1306_));
 sky130_fd_sc_hd__nand2_1 _2105_ (.A(net276),
    .B(_1306_),
    .Y(_1307_));
 sky130_fd_sc_hd__a311o_1 _2106_ (.A1(net222),
    .A2(_1305_),
    .A3(_1307_),
    .B1(_1303_),
    .C1(net235),
    .X(_1308_));
 sky130_fd_sc_hd__a311oi_4 _2107_ (.A1(net6),
    .A2(_1301_),
    .A3(_1308_),
    .B1(net219),
    .C1(_1294_),
    .Y(net47));
 sky130_fd_sc_hd__mux4_1 _2108_ (.A0(\mem[0][14] ),
    .A1(\mem[1][14] ),
    .A2(\mem[2][14] ),
    .A3(\mem[3][14] ),
    .S0(net343),
    .S1(net295),
    .X(_1309_));
 sky130_fd_sc_hd__mux4_1 _2109_ (.A0(\mem[4][14] ),
    .A1(\mem[5][14] ),
    .A2(\mem[6][14] ),
    .A3(\mem[7][14] ),
    .S0(net343),
    .S1(net295),
    .X(_1310_));
 sky130_fd_sc_hd__mux4_1 _2110_ (.A0(\mem[12][14] ),
    .A1(\mem[13][14] ),
    .A2(\mem[14][14] ),
    .A3(\mem[15][14] ),
    .S0(net343),
    .S1(net295),
    .X(_1311_));
 sky130_fd_sc_hd__mux4_1 _2111_ (.A0(\mem[8][14] ),
    .A1(\mem[9][14] ),
    .A2(\mem[10][14] ),
    .A3(\mem[11][14] ),
    .S0(net343),
    .S1(net295),
    .X(_1312_));
 sky130_fd_sc_hd__mux4_2 _2112_ (.A0(_1309_),
    .A1(_1310_),
    .A2(_1312_),
    .A3(_1311_),
    .S0(net248),
    .S1(net239),
    .X(_1313_));
 sky130_fd_sc_hd__nor2_1 _2113_ (.A(net233),
    .B(_1313_),
    .Y(_1314_));
 sky130_fd_sc_hd__mux4_1 _2114_ (.A0(\mem[24][14] ),
    .A1(\mem[25][14] ),
    .A2(\mem[26][14] ),
    .A3(\mem[27][14] ),
    .S0(net330),
    .S1(net281),
    .X(_1315_));
 sky130_fd_sc_hd__mux2_1 _2115_ (.A0(\mem[30][14] ),
    .A1(\mem[31][14] ),
    .S(net330),
    .X(_1316_));
 sky130_fd_sc_hd__nand2_1 _2116_ (.A(net281),
    .B(_1316_),
    .Y(_1317_));
 sky130_fd_sc_hd__mux2_1 _2117_ (.A0(\mem[28][14] ),
    .A1(\mem[29][14] ),
    .S(net330),
    .X(_1318_));
 sky130_fd_sc_hd__nand2b_1 _2118_ (.A_N(net281),
    .B(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__o21ai_1 _2119_ (.A1(net243),
    .A2(_1315_),
    .B1(net236),
    .Y(_1320_));
 sky130_fd_sc_hd__a31o_1 _2120_ (.A1(net243),
    .A2(_1317_),
    .A3(_1319_),
    .B1(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__mux4_1 _2121_ (.A0(\mem[20][14] ),
    .A1(\mem[21][14] ),
    .A2(\mem[22][14] ),
    .A3(\mem[23][14] ),
    .S0(net326),
    .S1(net278),
    .X(_1322_));
 sky130_fd_sc_hd__nor2_1 _2122_ (.A(net223),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__mux2_1 _2123_ (.A0(\mem[16][14] ),
    .A1(\mem[17][14] ),
    .S(net326),
    .X(_1324_));
 sky130_fd_sc_hd__nand2b_1 _2124_ (.A_N(net278),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__mux2_1 _2125_ (.A0(\mem[18][14] ),
    .A1(\mem[19][14] ),
    .S(net326),
    .X(_1326_));
 sky130_fd_sc_hd__nand2_1 _2126_ (.A(net278),
    .B(_1326_),
    .Y(_1327_));
 sky130_fd_sc_hd__a311o_1 _2127_ (.A1(net223),
    .A2(_1325_),
    .A3(_1327_),
    .B1(_1323_),
    .C1(net237),
    .X(_1328_));
 sky130_fd_sc_hd__a311oi_2 _2128_ (.A1(net233),
    .A2(_1321_),
    .A3(_1328_),
    .B1(net219),
    .C1(_1314_),
    .Y(net48));
 sky130_fd_sc_hd__mux4_1 _2129_ (.A0(\mem[0][15] ),
    .A1(\mem[1][15] ),
    .A2(\mem[2][15] ),
    .A3(\mem[3][15] ),
    .S0(net336),
    .S1(net288),
    .X(_1329_));
 sky130_fd_sc_hd__mux4_1 _2130_ (.A0(\mem[4][15] ),
    .A1(\mem[5][15] ),
    .A2(\mem[6][15] ),
    .A3(\mem[7][15] ),
    .S0(net336),
    .S1(net288),
    .X(_1330_));
 sky130_fd_sc_hd__mux4_1 _2131_ (.A0(\mem[12][15] ),
    .A1(\mem[13][15] ),
    .A2(\mem[14][15] ),
    .A3(\mem[15][15] ),
    .S0(net336),
    .S1(net288),
    .X(_1331_));
 sky130_fd_sc_hd__mux4_1 _2132_ (.A0(\mem[8][15] ),
    .A1(\mem[9][15] ),
    .A2(\mem[10][15] ),
    .A3(\mem[11][15] ),
    .S0(net336),
    .S1(net288),
    .X(_1332_));
 sky130_fd_sc_hd__mux4_2 _2133_ (.A0(_1329_),
    .A1(_1330_),
    .A2(_1332_),
    .A3(_1331_),
    .S0(net246),
    .S1(net238),
    .X(_1333_));
 sky130_fd_sc_hd__nor2_1 _2134_ (.A(net230),
    .B(_1333_),
    .Y(_1334_));
 sky130_fd_sc_hd__mux4_1 _2135_ (.A0(\mem[24][15] ),
    .A1(\mem[25][15] ),
    .A2(\mem[26][15] ),
    .A3(\mem[27][15] ),
    .S0(net320),
    .S1(net272),
    .X(_1335_));
 sky130_fd_sc_hd__mux2_1 _2136_ (.A0(\mem[30][15] ),
    .A1(\mem[31][15] ),
    .S(net324),
    .X(_1336_));
 sky130_fd_sc_hd__nand2_1 _2137_ (.A(net272),
    .B(_1336_),
    .Y(_1337_));
 sky130_fd_sc_hd__mux2_1 _2138_ (.A0(\mem[28][15] ),
    .A1(\mem[29][15] ),
    .S(net324),
    .X(_1338_));
 sky130_fd_sc_hd__nand2b_1 _2139_ (.A_N(net272),
    .B(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__o21ai_1 _2140_ (.A1(net241),
    .A2(_1335_),
    .B1(net234),
    .Y(_1340_));
 sky130_fd_sc_hd__a31o_1 _2141_ (.A1(net241),
    .A2(_1337_),
    .A3(_1339_),
    .B1(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__mux4_1 _2142_ (.A0(\mem[20][15] ),
    .A1(\mem[21][15] ),
    .A2(\mem[22][15] ),
    .A3(\mem[23][15] ),
    .S0(net319),
    .S1(net271),
    .X(_1342_));
 sky130_fd_sc_hd__nor2_1 _2143_ (.A(net220),
    .B(_1342_),
    .Y(_1343_));
 sky130_fd_sc_hd__mux2_1 _2144_ (.A0(\mem[16][15] ),
    .A1(\mem[17][15] ),
    .S(net319),
    .X(_1344_));
 sky130_fd_sc_hd__nand2b_1 _2145_ (.A_N(net271),
    .B(_1344_),
    .Y(_1345_));
 sky130_fd_sc_hd__mux2_1 _2146_ (.A0(\mem[18][15] ),
    .A1(\mem[19][15] ),
    .S(net319),
    .X(_1346_));
 sky130_fd_sc_hd__nand2_1 _2147_ (.A(net271),
    .B(_1346_),
    .Y(_1347_));
 sky130_fd_sc_hd__a311o_1 _2148_ (.A1(net220),
    .A2(_1345_),
    .A3(_1347_),
    .B1(_1343_),
    .C1(net234),
    .X(_1348_));
 sky130_fd_sc_hd__a311oi_4 _2149_ (.A1(net230),
    .A2(_1341_),
    .A3(_1348_),
    .B1(net218),
    .C1(_1334_),
    .Y(net49));
 sky130_fd_sc_hd__mux4_1 _2150_ (.A0(\mem[0][16] ),
    .A1(\mem[1][16] ),
    .A2(\mem[2][16] ),
    .A3(\mem[3][16] ),
    .S0(net339),
    .S1(net291),
    .X(_1349_));
 sky130_fd_sc_hd__mux4_1 _2151_ (.A0(\mem[4][16] ),
    .A1(\mem[5][16] ),
    .A2(\mem[6][16] ),
    .A3(\mem[7][16] ),
    .S0(net339),
    .S1(net291),
    .X(_1350_));
 sky130_fd_sc_hd__mux4_1 _2152_ (.A0(\mem[12][16] ),
    .A1(\mem[13][16] ),
    .A2(\mem[14][16] ),
    .A3(\mem[15][16] ),
    .S0(net339),
    .S1(net291),
    .X(_1351_));
 sky130_fd_sc_hd__mux4_1 _2153_ (.A0(\mem[8][16] ),
    .A1(\mem[9][16] ),
    .A2(\mem[10][16] ),
    .A3(\mem[11][16] ),
    .S0(net339),
    .S1(net291),
    .X(_1352_));
 sky130_fd_sc_hd__mux4_1 _2154_ (.A0(_1349_),
    .A1(_1350_),
    .A2(_1352_),
    .A3(_1351_),
    .S0(net247),
    .S1(net239),
    .X(_1353_));
 sky130_fd_sc_hd__nor2_2 _2155_ (.A(net232),
    .B(_1353_),
    .Y(_1354_));
 sky130_fd_sc_hd__mux4_1 _2156_ (.A0(\mem[24][16] ),
    .A1(\mem[25][16] ),
    .A2(\mem[26][16] ),
    .A3(\mem[27][16] ),
    .S0(net327),
    .S1(net279),
    .X(_1355_));
 sky130_fd_sc_hd__mux2_1 _2157_ (.A0(\mem[30][16] ),
    .A1(\mem[31][16] ),
    .S(net327),
    .X(_1356_));
 sky130_fd_sc_hd__nand2_1 _2158_ (.A(net279),
    .B(_1356_),
    .Y(_1357_));
 sky130_fd_sc_hd__mux2_1 _2159_ (.A0(\mem[28][16] ),
    .A1(\mem[29][16] ),
    .S(net327),
    .X(_1358_));
 sky130_fd_sc_hd__nand2b_1 _2160_ (.A_N(net279),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__o21ai_1 _2161_ (.A1(net244),
    .A2(_1355_),
    .B1(net237),
    .Y(_1360_));
 sky130_fd_sc_hd__a31o_1 _2162_ (.A1(net244),
    .A2(_1357_),
    .A3(_1359_),
    .B1(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__mux4_1 _2163_ (.A0(\mem[20][16] ),
    .A1(\mem[21][16] ),
    .A2(\mem[22][16] ),
    .A3(\mem[23][16] ),
    .S0(net326),
    .S1(net278),
    .X(_1362_));
 sky130_fd_sc_hd__nor2_1 _2164_ (.A(net223),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__mux2_1 _2165_ (.A0(\mem[16][16] ),
    .A1(\mem[17][16] ),
    .S(net326),
    .X(_1364_));
 sky130_fd_sc_hd__nand2b_1 _2166_ (.A_N(net278),
    .B(_1364_),
    .Y(_1365_));
 sky130_fd_sc_hd__mux2_1 _2167_ (.A0(\mem[18][16] ),
    .A1(\mem[19][16] ),
    .S(net326),
    .X(_1366_));
 sky130_fd_sc_hd__nand2_1 _2168_ (.A(net278),
    .B(_1366_),
    .Y(_1367_));
 sky130_fd_sc_hd__a311o_1 _2169_ (.A1(net223),
    .A2(_1365_),
    .A3(_1367_),
    .B1(_1363_),
    .C1(net237),
    .X(_1368_));
 sky130_fd_sc_hd__a311oi_4 _2170_ (.A1(net233),
    .A2(_1361_),
    .A3(_1368_),
    .B1(net219),
    .C1(_1354_),
    .Y(net50));
 sky130_fd_sc_hd__mux4_1 _2171_ (.A0(\mem[0][17] ),
    .A1(\mem[1][17] ),
    .A2(\mem[2][17] ),
    .A3(\mem[3][17] ),
    .S0(net344),
    .S1(net296),
    .X(_1369_));
 sky130_fd_sc_hd__mux4_1 _2172_ (.A0(\mem[4][17] ),
    .A1(\mem[5][17] ),
    .A2(\mem[6][17] ),
    .A3(\mem[7][17] ),
    .S0(net344),
    .S1(net296),
    .X(_1370_));
 sky130_fd_sc_hd__mux4_1 _2173_ (.A0(\mem[12][17] ),
    .A1(\mem[13][17] ),
    .A2(\mem[14][17] ),
    .A3(\mem[15][17] ),
    .S0(net343),
    .S1(net295),
    .X(_1371_));
 sky130_fd_sc_hd__mux4_1 _2174_ (.A0(\mem[8][17] ),
    .A1(\mem[9][17] ),
    .A2(\mem[10][17] ),
    .A3(\mem[11][17] ),
    .S0(net344),
    .S1(net296),
    .X(_1372_));
 sky130_fd_sc_hd__mux4_2 _2175_ (.A0(_1369_),
    .A1(_1370_),
    .A2(_1372_),
    .A3(_1371_),
    .S0(net248),
    .S1(net239),
    .X(_1373_));
 sky130_fd_sc_hd__nor2_1 _2176_ (.A(net231),
    .B(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__mux4_1 _2177_ (.A0(\mem[24][17] ),
    .A1(\mem[25][17] ),
    .A2(\mem[26][17] ),
    .A3(\mem[27][17] ),
    .S0(net329),
    .S1(net281),
    .X(_1375_));
 sky130_fd_sc_hd__mux2_1 _2178_ (.A0(\mem[30][17] ),
    .A1(\mem[31][17] ),
    .S(net329),
    .X(_1376_));
 sky130_fd_sc_hd__nand2_1 _2179_ (.A(net282),
    .B(_1376_),
    .Y(_1377_));
 sky130_fd_sc_hd__mux2_1 _2180_ (.A0(\mem[28][17] ),
    .A1(\mem[29][17] ),
    .S(net329),
    .X(_1378_));
 sky130_fd_sc_hd__nand2b_1 _2181_ (.A_N(net282),
    .B(_1378_),
    .Y(_1379_));
 sky130_fd_sc_hd__o21ai_1 _2182_ (.A1(net243),
    .A2(_1375_),
    .B1(net236),
    .Y(_1380_));
 sky130_fd_sc_hd__a31o_1 _2183_ (.A1(net243),
    .A2(_1377_),
    .A3(_1379_),
    .B1(_1380_),
    .X(_1381_));
 sky130_fd_sc_hd__mux4_1 _2184_ (.A0(\mem[20][17] ),
    .A1(\mem[21][17] ),
    .A2(\mem[22][17] ),
    .A3(\mem[23][17] ),
    .S0(net330),
    .S1(net281),
    .X(_1382_));
 sky130_fd_sc_hd__nor2_1 _2185_ (.A(net224),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__mux2_1 _2186_ (.A0(\mem[16][17] ),
    .A1(\mem[17][17] ),
    .S(net329),
    .X(_1384_));
 sky130_fd_sc_hd__nand2b_1 _2187_ (.A_N(net281),
    .B(_1384_),
    .Y(_1385_));
 sky130_fd_sc_hd__mux2_1 _2188_ (.A0(\mem[18][17] ),
    .A1(\mem[19][17] ),
    .S(net330),
    .X(_1386_));
 sky130_fd_sc_hd__nand2_1 _2189_ (.A(net281),
    .B(_1386_),
    .Y(_1387_));
 sky130_fd_sc_hd__a311o_1 _2190_ (.A1(net223),
    .A2(_1385_),
    .A3(_1387_),
    .B1(_1383_),
    .C1(net236),
    .X(_1388_));
 sky130_fd_sc_hd__a311oi_4 _2191_ (.A1(net231),
    .A2(_1381_),
    .A3(_1388_),
    .B1(net219),
    .C1(_1374_),
    .Y(net51));
 sky130_fd_sc_hd__mux4_1 _2192_ (.A0(\mem[0][18] ),
    .A1(\mem[1][18] ),
    .A2(\mem[2][18] ),
    .A3(\mem[3][18] ),
    .S0(net336),
    .S1(net288),
    .X(_1389_));
 sky130_fd_sc_hd__mux4_1 _2193_ (.A0(\mem[4][18] ),
    .A1(\mem[5][18] ),
    .A2(\mem[6][18] ),
    .A3(\mem[7][18] ),
    .S0(net336),
    .S1(net288),
    .X(_1390_));
 sky130_fd_sc_hd__mux4_1 _2194_ (.A0(\mem[12][18] ),
    .A1(\mem[13][18] ),
    .A2(\mem[14][18] ),
    .A3(\mem[15][18] ),
    .S0(net335),
    .S1(net286),
    .X(_1391_));
 sky130_fd_sc_hd__mux4_1 _2195_ (.A0(\mem[8][18] ),
    .A1(\mem[9][18] ),
    .A2(\mem[10][18] ),
    .A3(\mem[11][18] ),
    .S0(net335),
    .S1(net286),
    .X(_1392_));
 sky130_fd_sc_hd__mux4_1 _2196_ (.A0(_1389_),
    .A1(_1390_),
    .A2(_1392_),
    .A3(_1391_),
    .S0(net246),
    .S1(net238),
    .X(_1393_));
 sky130_fd_sc_hd__nor2_1 _2197_ (.A(net6),
    .B(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__mux4_1 _2198_ (.A0(\mem[24][18] ),
    .A1(\mem[25][18] ),
    .A2(\mem[26][18] ),
    .A3(\mem[27][18] ),
    .S0(net325),
    .S1(net277),
    .X(_1395_));
 sky130_fd_sc_hd__mux2_1 _2199_ (.A0(\mem[30][18] ),
    .A1(\mem[31][18] ),
    .S(net325),
    .X(_1396_));
 sky130_fd_sc_hd__nand2_1 _2200_ (.A(net277),
    .B(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__mux2_1 _2201_ (.A0(\mem[28][18] ),
    .A1(\mem[29][18] ),
    .S(net325),
    .X(_1398_));
 sky130_fd_sc_hd__nand2b_1 _2202_ (.A_N(net277),
    .B(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__o21ai_1 _2203_ (.A1(net242),
    .A2(_1395_),
    .B1(net235),
    .Y(_1400_));
 sky130_fd_sc_hd__a31o_1 _2204_ (.A1(net245),
    .A2(_1397_),
    .A3(_1399_),
    .B1(_1400_),
    .X(_1401_));
 sky130_fd_sc_hd__mux4_1 _2205_ (.A0(\mem[20][18] ),
    .A1(\mem[21][18] ),
    .A2(\mem[22][18] ),
    .A3(\mem[23][18] ),
    .S0(net324),
    .S1(net276),
    .X(_1402_));
 sky130_fd_sc_hd__nor2_1 _2206_ (.A(net221),
    .B(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__mux2_1 _2207_ (.A0(\mem[16][18] ),
    .A1(\mem[17][18] ),
    .S(net325),
    .X(_1404_));
 sky130_fd_sc_hd__nand2b_1 _2208_ (.A_N(net276),
    .B(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__mux2_1 _2209_ (.A0(\mem[18][18] ),
    .A1(\mem[19][18] ),
    .S(net324),
    .X(_1406_));
 sky130_fd_sc_hd__nand2_1 _2210_ (.A(net276),
    .B(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__a311o_1 _2211_ (.A1(net221),
    .A2(_1405_),
    .A3(_1407_),
    .B1(_1403_),
    .C1(net235),
    .X(_1408_));
 sky130_fd_sc_hd__a311oi_2 _2212_ (.A1(net6),
    .A2(_1401_),
    .A3(_1408_),
    .B1(net219),
    .C1(_1394_),
    .Y(net52));
 sky130_fd_sc_hd__mux4_1 _2213_ (.A0(\mem[0][19] ),
    .A1(\mem[1][19] ),
    .A2(\mem[2][19] ),
    .A3(\mem[3][19] ),
    .S0(net344),
    .S1(net296),
    .X(_1409_));
 sky130_fd_sc_hd__mux4_1 _2214_ (.A0(\mem[4][19] ),
    .A1(\mem[5][19] ),
    .A2(\mem[6][19] ),
    .A3(\mem[7][19] ),
    .S0(net344),
    .S1(net296),
    .X(_1410_));
 sky130_fd_sc_hd__mux4_1 _2215_ (.A0(\mem[12][19] ),
    .A1(\mem[13][19] ),
    .A2(\mem[14][19] ),
    .A3(\mem[15][19] ),
    .S0(net343),
    .S1(net295),
    .X(_1411_));
 sky130_fd_sc_hd__mux4_1 _2216_ (.A0(\mem[8][19] ),
    .A1(\mem[9][19] ),
    .A2(\mem[10][19] ),
    .A3(\mem[11][19] ),
    .S0(net344),
    .S1(net296),
    .X(_1412_));
 sky130_fd_sc_hd__mux4_2 _2217_ (.A0(_1409_),
    .A1(_1410_),
    .A2(_1412_),
    .A3(_1411_),
    .S0(net248),
    .S1(net239),
    .X(_1413_));
 sky130_fd_sc_hd__nor2_1 _2218_ (.A(net232),
    .B(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__mux4_1 _2219_ (.A0(\mem[24][19] ),
    .A1(\mem[25][19] ),
    .A2(\mem[26][19] ),
    .A3(\mem[27][19] ),
    .S0(net329),
    .S1(net282),
    .X(_1415_));
 sky130_fd_sc_hd__mux2_1 _2220_ (.A0(\mem[30][19] ),
    .A1(\mem[31][19] ),
    .S(net329),
    .X(_1416_));
 sky130_fd_sc_hd__nand2_1 _2221_ (.A(net282),
    .B(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__mux2_1 _2222_ (.A0(\mem[28][19] ),
    .A1(\mem[29][19] ),
    .S(net329),
    .X(_1418_));
 sky130_fd_sc_hd__nand2b_1 _2223_ (.A_N(net282),
    .B(_1418_),
    .Y(_1419_));
 sky130_fd_sc_hd__o21ai_1 _2224_ (.A1(net243),
    .A2(_1415_),
    .B1(net236),
    .Y(_1420_));
 sky130_fd_sc_hd__a31o_1 _2225_ (.A1(net243),
    .A2(_1417_),
    .A3(_1419_),
    .B1(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__mux4_1 _2226_ (.A0(\mem[20][19] ),
    .A1(\mem[21][19] ),
    .A2(\mem[22][19] ),
    .A3(\mem[23][19] ),
    .S0(net330),
    .S1(net281),
    .X(_1422_));
 sky130_fd_sc_hd__nor2_1 _2227_ (.A(net224),
    .B(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__mux2_1 _2228_ (.A0(\mem[16][19] ),
    .A1(\mem[17][19] ),
    .S(net329),
    .X(_1424_));
 sky130_fd_sc_hd__nand2b_1 _2229_ (.A_N(net281),
    .B(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__mux2_1 _2230_ (.A0(\mem[18][19] ),
    .A1(\mem[19][19] ),
    .S(net330),
    .X(_1426_));
 sky130_fd_sc_hd__nand2_1 _2231_ (.A(net281),
    .B(_1426_),
    .Y(_1427_));
 sky130_fd_sc_hd__a311o_1 _2232_ (.A1(net224),
    .A2(_1425_),
    .A3(_1427_),
    .B1(_1423_),
    .C1(net236),
    .X(_1428_));
 sky130_fd_sc_hd__a311oi_4 _2233_ (.A1(net232),
    .A2(_1421_),
    .A3(_1428_),
    .B1(net219),
    .C1(_1414_),
    .Y(net53));
 sky130_fd_sc_hd__mux4_1 _2234_ (.A0(\mem[0][20] ),
    .A1(\mem[1][20] ),
    .A2(\mem[2][20] ),
    .A3(\mem[3][20] ),
    .S0(net343),
    .S1(net295),
    .X(_1429_));
 sky130_fd_sc_hd__mux4_1 _2235_ (.A0(\mem[4][20] ),
    .A1(\mem[5][20] ),
    .A2(\mem[6][20] ),
    .A3(\mem[7][20] ),
    .S0(net344),
    .S1(net296),
    .X(_1430_));
 sky130_fd_sc_hd__mux4_1 _2236_ (.A0(\mem[12][20] ),
    .A1(\mem[13][20] ),
    .A2(\mem[14][20] ),
    .A3(\mem[15][20] ),
    .S0(net343),
    .S1(net295),
    .X(_1431_));
 sky130_fd_sc_hd__mux4_1 _2237_ (.A0(\mem[8][20] ),
    .A1(\mem[9][20] ),
    .A2(\mem[10][20] ),
    .A3(\mem[11][20] ),
    .S0(net344),
    .S1(net296),
    .X(_1432_));
 sky130_fd_sc_hd__mux4_2 _2238_ (.A0(_1429_),
    .A1(_1430_),
    .A2(_1432_),
    .A3(_1431_),
    .S0(net248),
    .S1(net239),
    .X(_1433_));
 sky130_fd_sc_hd__nor2_2 _2239_ (.A(net231),
    .B(_1433_),
    .Y(_1434_));
 sky130_fd_sc_hd__mux4_1 _2240_ (.A0(\mem[24][20] ),
    .A1(\mem[25][20] ),
    .A2(\mem[26][20] ),
    .A3(\mem[27][20] ),
    .S0(net327),
    .S1(net279),
    .X(_1435_));
 sky130_fd_sc_hd__mux2_1 _2241_ (.A0(\mem[30][20] ),
    .A1(\mem[31][20] ),
    .S(net328),
    .X(_1436_));
 sky130_fd_sc_hd__nand2_1 _2242_ (.A(net280),
    .B(_1436_),
    .Y(_1437_));
 sky130_fd_sc_hd__mux2_1 _2243_ (.A0(\mem[28][20] ),
    .A1(\mem[29][20] ),
    .S(net328),
    .X(_1438_));
 sky130_fd_sc_hd__nand2b_1 _2244_ (.A_N(net280),
    .B(_1438_),
    .Y(_1439_));
 sky130_fd_sc_hd__o21ai_1 _2245_ (.A1(net244),
    .A2(_1435_),
    .B1(net237),
    .Y(_1440_));
 sky130_fd_sc_hd__a31o_1 _2246_ (.A1(net244),
    .A2(_1437_),
    .A3(_1439_),
    .B1(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__mux4_1 _2247_ (.A0(\mem[20][20] ),
    .A1(\mem[21][20] ),
    .A2(\mem[22][20] ),
    .A3(\mem[23][20] ),
    .S0(net328),
    .S1(net280),
    .X(_1442_));
 sky130_fd_sc_hd__nor2_1 _2248_ (.A(net223),
    .B(_1442_),
    .Y(_1443_));
 sky130_fd_sc_hd__mux2_1 _2249_ (.A0(\mem[16][20] ),
    .A1(\mem[17][20] ),
    .S(net328),
    .X(_1444_));
 sky130_fd_sc_hd__nand2b_1 _2250_ (.A_N(net280),
    .B(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__mux2_1 _2251_ (.A0(\mem[18][20] ),
    .A1(\mem[19][20] ),
    .S(net328),
    .X(_1446_));
 sky130_fd_sc_hd__nand2_1 _2252_ (.A(net280),
    .B(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__a311o_1 _2253_ (.A1(net223),
    .A2(_1445_),
    .A3(_1447_),
    .B1(_1443_),
    .C1(net237),
    .X(_1448_));
 sky130_fd_sc_hd__a311oi_4 _2254_ (.A1(net233),
    .A2(_1441_),
    .A3(_1448_),
    .B1(net219),
    .C1(_1434_),
    .Y(net55));
 sky130_fd_sc_hd__mux4_1 _2255_ (.A0(\mem[0][21] ),
    .A1(\mem[1][21] ),
    .A2(\mem[2][21] ),
    .A3(\mem[3][21] ),
    .S0(net338),
    .S1(net290),
    .X(_1449_));
 sky130_fd_sc_hd__mux4_1 _2256_ (.A0(\mem[4][21] ),
    .A1(\mem[5][21] ),
    .A2(\mem[6][21] ),
    .A3(\mem[7][21] ),
    .S0(net338),
    .S1(net290),
    .X(_1450_));
 sky130_fd_sc_hd__mux4_1 _2257_ (.A0(\mem[12][21] ),
    .A1(\mem[13][21] ),
    .A2(\mem[14][21] ),
    .A3(\mem[15][21] ),
    .S0(net336),
    .S1(net288),
    .X(_1451_));
 sky130_fd_sc_hd__mux4_1 _2258_ (.A0(\mem[8][21] ),
    .A1(\mem[9][21] ),
    .A2(\mem[10][21] ),
    .A3(\mem[11][21] ),
    .S0(net338),
    .S1(net290),
    .X(_1452_));
 sky130_fd_sc_hd__mux4_2 _2259_ (.A0(_1449_),
    .A1(_1450_),
    .A2(_1452_),
    .A3(_1451_),
    .S0(net246),
    .S1(net238),
    .X(_1453_));
 sky130_fd_sc_hd__nor2_1 _2260_ (.A(net230),
    .B(_1453_),
    .Y(_1454_));
 sky130_fd_sc_hd__mux4_1 _2261_ (.A0(\mem[24][21] ),
    .A1(\mem[25][21] ),
    .A2(\mem[26][21] ),
    .A3(\mem[27][21] ),
    .S0(net320),
    .S1(net272),
    .X(_1455_));
 sky130_fd_sc_hd__mux2_1 _2262_ (.A0(\mem[30][21] ),
    .A1(\mem[31][21] ),
    .S(net324),
    .X(_1456_));
 sky130_fd_sc_hd__nand2_1 _2263_ (.A(net272),
    .B(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__mux2_1 _2264_ (.A0(\mem[28][21] ),
    .A1(\mem[29][21] ),
    .S(net324),
    .X(_1458_));
 sky130_fd_sc_hd__nand2b_1 _2265_ (.A_N(net272),
    .B(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__o21ai_1 _2266_ (.A1(net241),
    .A2(_1455_),
    .B1(net234),
    .Y(_1460_));
 sky130_fd_sc_hd__a31o_1 _2267_ (.A1(net241),
    .A2(_1457_),
    .A3(_1459_),
    .B1(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__mux4_1 _2268_ (.A0(\mem[20][21] ),
    .A1(\mem[21][21] ),
    .A2(\mem[22][21] ),
    .A3(\mem[23][21] ),
    .S0(net320),
    .S1(net272),
    .X(_1462_));
 sky130_fd_sc_hd__nor2_1 _2269_ (.A(net221),
    .B(_1462_),
    .Y(_1463_));
 sky130_fd_sc_hd__mux2_1 _2270_ (.A0(\mem[16][21] ),
    .A1(\mem[17][21] ),
    .S(net324),
    .X(_1464_));
 sky130_fd_sc_hd__nand2b_1 _2271_ (.A_N(net272),
    .B(_1464_),
    .Y(_1465_));
 sky130_fd_sc_hd__mux2_1 _2272_ (.A0(\mem[18][21] ),
    .A1(\mem[19][21] ),
    .S(net320),
    .X(_1466_));
 sky130_fd_sc_hd__nand2_1 _2273_ (.A(net272),
    .B(_1466_),
    .Y(_1467_));
 sky130_fd_sc_hd__a311o_1 _2274_ (.A1(net221),
    .A2(_1465_),
    .A3(_1467_),
    .B1(_1463_),
    .C1(net235),
    .X(_1468_));
 sky130_fd_sc_hd__a311oi_2 _2275_ (.A1(net230),
    .A2(_1461_),
    .A3(_1468_),
    .B1(net218),
    .C1(_1454_),
    .Y(net56));
 sky130_fd_sc_hd__mux4_1 _2276_ (.A0(\mem[0][22] ),
    .A1(\mem[1][22] ),
    .A2(\mem[2][22] ),
    .A3(\mem[3][22] ),
    .S0(net336),
    .S1(net288),
    .X(_1469_));
 sky130_fd_sc_hd__mux4_1 _2277_ (.A0(\mem[4][22] ),
    .A1(\mem[5][22] ),
    .A2(\mem[6][22] ),
    .A3(\mem[7][22] ),
    .S0(net337),
    .S1(net289),
    .X(_1470_));
 sky130_fd_sc_hd__mux4_1 _2278_ (.A0(\mem[12][22] ),
    .A1(\mem[13][22] ),
    .A2(\mem[14][22] ),
    .A3(\mem[15][22] ),
    .S0(net337),
    .S1(net289),
    .X(_1471_));
 sky130_fd_sc_hd__mux4_1 _2279_ (.A0(\mem[8][22] ),
    .A1(\mem[9][22] ),
    .A2(\mem[10][22] ),
    .A3(\mem[11][22] ),
    .S0(net336),
    .S1(net288),
    .X(_1472_));
 sky130_fd_sc_hd__mux4_2 _2280_ (.A0(_1469_),
    .A1(_1470_),
    .A2(_1472_),
    .A3(_1471_),
    .S0(net246),
    .S1(net240),
    .X(_1473_));
 sky130_fd_sc_hd__nor2_1 _2281_ (.A(net229),
    .B(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__mux4_1 _2282_ (.A0(\mem[24][22] ),
    .A1(\mem[25][22] ),
    .A2(\mem[26][22] ),
    .A3(\mem[27][22] ),
    .S0(net323),
    .S1(net275),
    .X(_1475_));
 sky130_fd_sc_hd__mux2_1 _2283_ (.A0(\mem[30][22] ),
    .A1(\mem[31][22] ),
    .S(net325),
    .X(_1476_));
 sky130_fd_sc_hd__nand2_1 _2284_ (.A(net277),
    .B(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__mux2_1 _2285_ (.A0(\mem[28][22] ),
    .A1(\mem[29][22] ),
    .S(net335),
    .X(_1478_));
 sky130_fd_sc_hd__nand2b_1 _2286_ (.A_N(net277),
    .B(_1478_),
    .Y(_1479_));
 sky130_fd_sc_hd__o21ai_1 _2287_ (.A1(net242),
    .A2(_1475_),
    .B1(net235),
    .Y(_1480_));
 sky130_fd_sc_hd__a31o_1 _2288_ (.A1(net245),
    .A2(_1477_),
    .A3(_1479_),
    .B1(_1480_),
    .X(_1481_));
 sky130_fd_sc_hd__mux4_1 _2289_ (.A0(\mem[20][22] ),
    .A1(\mem[21][22] ),
    .A2(\mem[22][22] ),
    .A3(\mem[23][22] ),
    .S0(net322),
    .S1(net274),
    .X(_1482_));
 sky130_fd_sc_hd__nor2_1 _2290_ (.A(net221),
    .B(_1482_),
    .Y(_1483_));
 sky130_fd_sc_hd__mux2_1 _2291_ (.A0(\mem[16][22] ),
    .A1(\mem[17][22] ),
    .S(net322),
    .X(_1484_));
 sky130_fd_sc_hd__nand2b_1 _2292_ (.A_N(net274),
    .B(_1484_),
    .Y(_1485_));
 sky130_fd_sc_hd__mux2_1 _2293_ (.A0(\mem[18][22] ),
    .A1(\mem[19][22] ),
    .S(net322),
    .X(_1486_));
 sky130_fd_sc_hd__nand2_1 _2294_ (.A(net274),
    .B(_1486_),
    .Y(_1487_));
 sky130_fd_sc_hd__a311o_1 _2295_ (.A1(net221),
    .A2(_1485_),
    .A3(_1487_),
    .B1(_1483_),
    .C1(net235),
    .X(_1488_));
 sky130_fd_sc_hd__a311oi_4 _2296_ (.A1(net229),
    .A2(_1481_),
    .A3(_1488_),
    .B1(net218),
    .C1(_1474_),
    .Y(net57));
 sky130_fd_sc_hd__mux4_1 _2297_ (.A0(\mem[0][23] ),
    .A1(\mem[1][23] ),
    .A2(\mem[2][23] ),
    .A3(\mem[3][23] ),
    .S0(net338),
    .S1(net290),
    .X(_1489_));
 sky130_fd_sc_hd__mux4_1 _2298_ (.A0(\mem[4][23] ),
    .A1(\mem[5][23] ),
    .A2(\mem[6][23] ),
    .A3(\mem[7][23] ),
    .S0(net337),
    .S1(net289),
    .X(_1490_));
 sky130_fd_sc_hd__mux4_1 _2299_ (.A0(\mem[12][23] ),
    .A1(\mem[13][23] ),
    .A2(\mem[14][23] ),
    .A3(\mem[15][23] ),
    .S0(net337),
    .S1(net289),
    .X(_1491_));
 sky130_fd_sc_hd__mux4_1 _2300_ (.A0(\mem[8][23] ),
    .A1(\mem[9][23] ),
    .A2(\mem[10][23] ),
    .A3(\mem[11][23] ),
    .S0(net336),
    .S1(net288),
    .X(_1492_));
 sky130_fd_sc_hd__mux4_2 _2301_ (.A0(_1489_),
    .A1(_1490_),
    .A2(_1492_),
    .A3(_1491_),
    .S0(net246),
    .S1(net240),
    .X(_1493_));
 sky130_fd_sc_hd__nor2_1 _2302_ (.A(net229),
    .B(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__mux4_1 _2303_ (.A0(\mem[24][23] ),
    .A1(\mem[25][23] ),
    .A2(\mem[26][23] ),
    .A3(\mem[27][23] ),
    .S0(net323),
    .S1(net275),
    .X(_1495_));
 sky130_fd_sc_hd__mux2_1 _2304_ (.A0(\mem[30][23] ),
    .A1(\mem[31][23] ),
    .S(net323),
    .X(_1496_));
 sky130_fd_sc_hd__nand2_1 _2305_ (.A(net275),
    .B(_1496_),
    .Y(_1497_));
 sky130_fd_sc_hd__mux2_1 _2306_ (.A0(\mem[28][23] ),
    .A1(\mem[29][23] ),
    .S(net323),
    .X(_1498_));
 sky130_fd_sc_hd__nand2b_1 _2307_ (.A_N(net274),
    .B(_1498_),
    .Y(_1499_));
 sky130_fd_sc_hd__o21ai_1 _2308_ (.A1(net242),
    .A2(_1495_),
    .B1(net240),
    .Y(_1500_));
 sky130_fd_sc_hd__a31o_1 _2309_ (.A1(net242),
    .A2(_1497_),
    .A3(_1499_),
    .B1(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__mux4_1 _2310_ (.A0(\mem[20][23] ),
    .A1(\mem[21][23] ),
    .A2(\mem[22][23] ),
    .A3(\mem[23][23] ),
    .S0(net324),
    .S1(net276),
    .X(_1502_));
 sky130_fd_sc_hd__nor2_1 _2311_ (.A(net221),
    .B(_1502_),
    .Y(_1503_));
 sky130_fd_sc_hd__mux2_1 _2312_ (.A0(\mem[16][23] ),
    .A1(\mem[17][23] ),
    .S(net325),
    .X(_1504_));
 sky130_fd_sc_hd__nand2b_1 _2313_ (.A_N(net277),
    .B(_1504_),
    .Y(_1505_));
 sky130_fd_sc_hd__mux2_1 _2314_ (.A0(\mem[18][23] ),
    .A1(\mem[19][23] ),
    .S(net324),
    .X(_1506_));
 sky130_fd_sc_hd__nand2_1 _2315_ (.A(net276),
    .B(_1506_),
    .Y(_1507_));
 sky130_fd_sc_hd__a311o_1 _2316_ (.A1(net221),
    .A2(_1505_),
    .A3(_1507_),
    .B1(_1503_),
    .C1(net240),
    .X(_1508_));
 sky130_fd_sc_hd__a311oi_4 _2317_ (.A1(net6),
    .A2(_1501_),
    .A3(_1508_),
    .B1(net218),
    .C1(_1494_),
    .Y(net58));
 sky130_fd_sc_hd__mux4_1 _2318_ (.A0(\mem[0][24] ),
    .A1(\mem[1][24] ),
    .A2(\mem[2][24] ),
    .A3(\mem[3][24] ),
    .S0(net334),
    .S1(net287),
    .X(_1509_));
 sky130_fd_sc_hd__mux4_1 _2319_ (.A0(\mem[4][24] ),
    .A1(\mem[5][24] ),
    .A2(\mem[6][24] ),
    .A3(\mem[7][24] ),
    .S0(net334),
    .S1(net287),
    .X(_1510_));
 sky130_fd_sc_hd__mux4_1 _2320_ (.A0(\mem[12][24] ),
    .A1(\mem[13][24] ),
    .A2(\mem[14][24] ),
    .A3(\mem[15][24] ),
    .S0(net334),
    .S1(net287),
    .X(_1511_));
 sky130_fd_sc_hd__mux4_1 _2321_ (.A0(\mem[8][24] ),
    .A1(\mem[9][24] ),
    .A2(\mem[10][24] ),
    .A3(\mem[11][24] ),
    .S0(net334),
    .S1(net287),
    .X(_1512_));
 sky130_fd_sc_hd__mux4_2 _2322_ (.A0(_1509_),
    .A1(_1510_),
    .A2(_1512_),
    .A3(_1511_),
    .S0(net245),
    .S1(net238),
    .X(_1513_));
 sky130_fd_sc_hd__nor2_2 _2323_ (.A(net229),
    .B(_1513_),
    .Y(_1514_));
 sky130_fd_sc_hd__mux4_1 _2324_ (.A0(\mem[24][24] ),
    .A1(\mem[25][24] ),
    .A2(\mem[26][24] ),
    .A3(\mem[27][24] ),
    .S0(net322),
    .S1(net274),
    .X(_1515_));
 sky130_fd_sc_hd__mux2_1 _2325_ (.A0(\mem[30][24] ),
    .A1(\mem[31][24] ),
    .S(net322),
    .X(_1516_));
 sky130_fd_sc_hd__nand2_1 _2326_ (.A(net274),
    .B(_1516_),
    .Y(_1517_));
 sky130_fd_sc_hd__mux2_1 _2327_ (.A0(\mem[28][24] ),
    .A1(\mem[29][24] ),
    .S(net322),
    .X(_1518_));
 sky130_fd_sc_hd__nand2b_1 _2328_ (.A_N(net274),
    .B(_1518_),
    .Y(_1519_));
 sky130_fd_sc_hd__o21ai_1 _2329_ (.A1(net242),
    .A2(_1515_),
    .B1(net240),
    .Y(_1520_));
 sky130_fd_sc_hd__a31o_1 _2330_ (.A1(net242),
    .A2(_1517_),
    .A3(_1519_),
    .B1(_1520_),
    .X(_1521_));
 sky130_fd_sc_hd__mux4_1 _2331_ (.A0(\mem[20][24] ),
    .A1(\mem[21][24] ),
    .A2(\mem[22][24] ),
    .A3(\mem[23][24] ),
    .S0(net318),
    .S1(net270),
    .X(_1522_));
 sky130_fd_sc_hd__nor2_1 _2332_ (.A(net220),
    .B(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__mux2_1 _2333_ (.A0(\mem[16][24] ),
    .A1(\mem[17][24] ),
    .S(net318),
    .X(_1524_));
 sky130_fd_sc_hd__nand2b_1 _2334_ (.A_N(net270),
    .B(_1524_),
    .Y(_1525_));
 sky130_fd_sc_hd__mux2_1 _2335_ (.A0(\mem[18][24] ),
    .A1(\mem[19][24] ),
    .S(net318),
    .X(_1526_));
 sky130_fd_sc_hd__nand2_1 _2336_ (.A(net270),
    .B(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__a311o_2 _2337_ (.A1(net220),
    .A2(_1525_),
    .A3(_1527_),
    .B1(_1523_),
    .C1(net234),
    .X(_1528_));
 sky130_fd_sc_hd__a311oi_4 _2338_ (.A1(net230),
    .A2(_1521_),
    .A3(_1528_),
    .B1(net218),
    .C1(_1514_),
    .Y(net59));
 sky130_fd_sc_hd__mux4_1 _2339_ (.A0(\mem[0][25] ),
    .A1(\mem[1][25] ),
    .A2(\mem[2][25] ),
    .A3(\mem[3][25] ),
    .S0(net335),
    .S1(net286),
    .X(_1529_));
 sky130_fd_sc_hd__mux4_1 _2340_ (.A0(\mem[4][25] ),
    .A1(\mem[5][25] ),
    .A2(\mem[6][25] ),
    .A3(\mem[7][25] ),
    .S0(net334),
    .S1(net287),
    .X(_1530_));
 sky130_fd_sc_hd__mux4_1 _2341_ (.A0(\mem[12][25] ),
    .A1(\mem[13][25] ),
    .A2(\mem[14][25] ),
    .A3(\mem[15][25] ),
    .S0(net334),
    .S1(net287),
    .X(_1531_));
 sky130_fd_sc_hd__mux4_1 _2342_ (.A0(\mem[8][25] ),
    .A1(\mem[9][25] ),
    .A2(\mem[10][25] ),
    .A3(\mem[11][25] ),
    .S0(net334),
    .S1(net287),
    .X(_1532_));
 sky130_fd_sc_hd__mux4_1 _2343_ (.A0(_1529_),
    .A1(_1530_),
    .A2(_1532_),
    .A3(_1531_),
    .S0(net246),
    .S1(net240),
    .X(_1533_));
 sky130_fd_sc_hd__nor2_1 _2344_ (.A(net229),
    .B(_1533_),
    .Y(_1534_));
 sky130_fd_sc_hd__mux4_1 _2345_ (.A0(\mem[24][25] ),
    .A1(\mem[25][25] ),
    .A2(\mem[26][25] ),
    .A3(\mem[27][25] ),
    .S0(net323),
    .S1(net275),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_1 _2346_ (.A0(\mem[30][25] ),
    .A1(\mem[31][25] ),
    .S(net323),
    .X(_1536_));
 sky130_fd_sc_hd__nand2_1 _2347_ (.A(net275),
    .B(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__mux2_1 _2348_ (.A0(\mem[28][25] ),
    .A1(\mem[29][25] ),
    .S(net334),
    .X(_1538_));
 sky130_fd_sc_hd__nand2b_1 _2349_ (.A_N(net275),
    .B(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__o21ai_1 _2350_ (.A1(net245),
    .A2(_1535_),
    .B1(net238),
    .Y(_1540_));
 sky130_fd_sc_hd__a31o_1 _2351_ (.A1(net245),
    .A2(_1537_),
    .A3(_1539_),
    .B1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__mux4_1 _2352_ (.A0(\mem[20][25] ),
    .A1(\mem[21][25] ),
    .A2(\mem[22][25] ),
    .A3(\mem[23][25] ),
    .S0(net322),
    .S1(net274),
    .X(_1542_));
 sky130_fd_sc_hd__nor2_1 _2353_ (.A(net221),
    .B(_1542_),
    .Y(_1543_));
 sky130_fd_sc_hd__mux2_1 _2354_ (.A0(\mem[16][25] ),
    .A1(\mem[17][25] ),
    .S(net323),
    .X(_1544_));
 sky130_fd_sc_hd__nand2b_1 _2355_ (.A_N(net275),
    .B(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__mux2_1 _2356_ (.A0(\mem[18][25] ),
    .A1(\mem[19][25] ),
    .S(net323),
    .X(_1546_));
 sky130_fd_sc_hd__nand2_1 _2357_ (.A(net274),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__a311o_1 _2358_ (.A1(net221),
    .A2(_1545_),
    .A3(_1547_),
    .B1(_1543_),
    .C1(net240),
    .X(_1548_));
 sky130_fd_sc_hd__a311oi_4 _2359_ (.A1(net229),
    .A2(_1541_),
    .A3(_1548_),
    .B1(net218),
    .C1(_1534_),
    .Y(net60));
 sky130_fd_sc_hd__mux4_1 _2360_ (.A0(\mem[0][26] ),
    .A1(\mem[1][26] ),
    .A2(\mem[2][26] ),
    .A3(\mem[3][26] ),
    .S0(net335),
    .S1(net286),
    .X(_1549_));
 sky130_fd_sc_hd__mux4_1 _2361_ (.A0(\mem[4][26] ),
    .A1(\mem[5][26] ),
    .A2(\mem[6][26] ),
    .A3(\mem[7][26] ),
    .S0(net335),
    .S1(net286),
    .X(_1550_));
 sky130_fd_sc_hd__mux4_1 _2362_ (.A0(\mem[12][26] ),
    .A1(\mem[13][26] ),
    .A2(\mem[14][26] ),
    .A3(\mem[15][26] ),
    .S0(net335),
    .S1(net286),
    .X(_1551_));
 sky130_fd_sc_hd__mux4_1 _2363_ (.A0(\mem[8][26] ),
    .A1(\mem[9][26] ),
    .A2(\mem[10][26] ),
    .A3(\mem[11][26] ),
    .S0(net335),
    .S1(net286),
    .X(_1552_));
 sky130_fd_sc_hd__mux4_1 _2364_ (.A0(_1549_),
    .A1(_1550_),
    .A2(_1552_),
    .A3(_1551_),
    .S0(net245),
    .S1(net238),
    .X(_1553_));
 sky130_fd_sc_hd__nor2_1 _2365_ (.A(net229),
    .B(_1553_),
    .Y(_1554_));
 sky130_fd_sc_hd__mux4_1 _2366_ (.A0(\mem[24][26] ),
    .A1(\mem[25][26] ),
    .A2(\mem[26][26] ),
    .A3(\mem[27][26] ),
    .S0(net323),
    .S1(net275),
    .X(_1555_));
 sky130_fd_sc_hd__mux2_1 _2367_ (.A0(\mem[30][26] ),
    .A1(\mem[31][26] ),
    .S(net323),
    .X(_1556_));
 sky130_fd_sc_hd__nand2_1 _2368_ (.A(net275),
    .B(_1556_),
    .Y(_1557_));
 sky130_fd_sc_hd__mux2_1 _2369_ (.A0(\mem[28][26] ),
    .A1(\mem[29][26] ),
    .S(net323),
    .X(_1558_));
 sky130_fd_sc_hd__nand2b_1 _2370_ (.A_N(net275),
    .B(_1558_),
    .Y(_1559_));
 sky130_fd_sc_hd__o21ai_1 _2371_ (.A1(net242),
    .A2(_1555_),
    .B1(net240),
    .Y(_1560_));
 sky130_fd_sc_hd__a31o_1 _2372_ (.A1(net245),
    .A2(_1557_),
    .A3(_1559_),
    .B1(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__mux4_1 _2373_ (.A0(\mem[20][26] ),
    .A1(\mem[21][26] ),
    .A2(\mem[22][26] ),
    .A3(\mem[23][26] ),
    .S0(net319),
    .S1(net271),
    .X(_1562_));
 sky130_fd_sc_hd__nor2_1 _2374_ (.A(net222),
    .B(_1562_),
    .Y(_1563_));
 sky130_fd_sc_hd__mux2_1 _2375_ (.A0(\mem[16][26] ),
    .A1(\mem[17][26] ),
    .S(net319),
    .X(_1564_));
 sky130_fd_sc_hd__nand2b_1 _2376_ (.A_N(net271),
    .B(_1564_),
    .Y(_1565_));
 sky130_fd_sc_hd__mux2_1 _2377_ (.A0(\mem[18][26] ),
    .A1(\mem[19][26] ),
    .S(net319),
    .X(_1566_));
 sky130_fd_sc_hd__nand2_1 _2378_ (.A(net271),
    .B(_1566_),
    .Y(_1567_));
 sky130_fd_sc_hd__a311o_2 _2379_ (.A1(net220),
    .A2(_1565_),
    .A3(_1567_),
    .B1(_1563_),
    .C1(net235),
    .X(_1568_));
 sky130_fd_sc_hd__a311oi_2 _2380_ (.A1(net229),
    .A2(_1561_),
    .A3(_1568_),
    .B1(net218),
    .C1(_1554_),
    .Y(net61));
 sky130_fd_sc_hd__mux4_1 _2381_ (.A0(\mem[0][27] ),
    .A1(\mem[1][27] ),
    .A2(\mem[2][27] ),
    .A3(\mem[3][27] ),
    .S0(net339),
    .S1(net291),
    .X(_1569_));
 sky130_fd_sc_hd__mux4_1 _2382_ (.A0(\mem[4][27] ),
    .A1(\mem[5][27] ),
    .A2(\mem[6][27] ),
    .A3(\mem[7][27] ),
    .S0(net341),
    .S1(net293),
    .X(_1570_));
 sky130_fd_sc_hd__mux4_1 _2383_ (.A0(\mem[12][27] ),
    .A1(\mem[13][27] ),
    .A2(\mem[14][27] ),
    .A3(\mem[15][27] ),
    .S0(net339),
    .S1(net291),
    .X(_1571_));
 sky130_fd_sc_hd__mux4_1 _2384_ (.A0(\mem[8][27] ),
    .A1(\mem[9][27] ),
    .A2(\mem[10][27] ),
    .A3(\mem[11][27] ),
    .S0(net341),
    .S1(net293),
    .X(_1572_));
 sky130_fd_sc_hd__mux4_2 _2385_ (.A0(_1569_),
    .A1(_1570_),
    .A2(_1572_),
    .A3(_1571_),
    .S0(net248),
    .S1(net240),
    .X(_1573_));
 sky130_fd_sc_hd__nor2_2 _2386_ (.A(net231),
    .B(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__mux4_1 _2387_ (.A0(\mem[24][27] ),
    .A1(\mem[25][27] ),
    .A2(\mem[26][27] ),
    .A3(\mem[27][27] ),
    .S0(net327),
    .S1(net279),
    .X(_1575_));
 sky130_fd_sc_hd__mux2_1 _2388_ (.A0(\mem[30][27] ),
    .A1(\mem[31][27] ),
    .S(net327),
    .X(_1576_));
 sky130_fd_sc_hd__nand2_1 _2389_ (.A(net279),
    .B(_1576_),
    .Y(_1577_));
 sky130_fd_sc_hd__mux2_1 _2390_ (.A0(\mem[28][27] ),
    .A1(\mem[29][27] ),
    .S(net327),
    .X(_1578_));
 sky130_fd_sc_hd__nand2b_1 _2391_ (.A_N(net279),
    .B(_1578_),
    .Y(_1579_));
 sky130_fd_sc_hd__o21ai_1 _2392_ (.A1(net244),
    .A2(_1575_),
    .B1(net237),
    .Y(_1580_));
 sky130_fd_sc_hd__a31o_1 _2393_ (.A1(net244),
    .A2(_1577_),
    .A3(_1579_),
    .B1(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__mux4_1 _2394_ (.A0(\mem[20][27] ),
    .A1(\mem[21][27] ),
    .A2(\mem[22][27] ),
    .A3(\mem[23][27] ),
    .S0(net326),
    .S1(net278),
    .X(_1582_));
 sky130_fd_sc_hd__nor2_1 _2395_ (.A(net223),
    .B(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__mux2_1 _2396_ (.A0(\mem[16][27] ),
    .A1(\mem[17][27] ),
    .S(net326),
    .X(_1584_));
 sky130_fd_sc_hd__nand2b_1 _2397_ (.A_N(net278),
    .B(_1584_),
    .Y(_1585_));
 sky130_fd_sc_hd__mux2_1 _2398_ (.A0(\mem[18][27] ),
    .A1(\mem[19][27] ),
    .S(net328),
    .X(_1586_));
 sky130_fd_sc_hd__nand2_1 _2399_ (.A(net280),
    .B(_1586_),
    .Y(_1587_));
 sky130_fd_sc_hd__a311o_1 _2400_ (.A1(net223),
    .A2(_1585_),
    .A3(_1587_),
    .B1(_1583_),
    .C1(net237),
    .X(_1588_));
 sky130_fd_sc_hd__a311oi_4 _2401_ (.A1(net233),
    .A2(_1581_),
    .A3(_1588_),
    .B1(net219),
    .C1(_1574_),
    .Y(net62));
 sky130_fd_sc_hd__mux4_1 _2402_ (.A0(\mem[0][28] ),
    .A1(\mem[1][28] ),
    .A2(\mem[2][28] ),
    .A3(\mem[3][28] ),
    .S0(net338),
    .S1(net286),
    .X(_1589_));
 sky130_fd_sc_hd__mux4_1 _2403_ (.A0(\mem[4][28] ),
    .A1(\mem[5][28] ),
    .A2(\mem[6][28] ),
    .A3(\mem[7][28] ),
    .S0(net335),
    .S1(net286),
    .X(_1590_));
 sky130_fd_sc_hd__mux4_1 _2404_ (.A0(\mem[12][28] ),
    .A1(\mem[13][28] ),
    .A2(\mem[14][28] ),
    .A3(\mem[15][28] ),
    .S0(net335),
    .S1(net286),
    .X(_1591_));
 sky130_fd_sc_hd__mux4_1 _2405_ (.A0(\mem[8][28] ),
    .A1(\mem[9][28] ),
    .A2(\mem[10][28] ),
    .A3(\mem[11][28] ),
    .S0(net335),
    .S1(net286),
    .X(_1592_));
 sky130_fd_sc_hd__mux4_1 _2406_ (.A0(_1589_),
    .A1(_1590_),
    .A2(_1592_),
    .A3(_1591_),
    .S0(net245),
    .S1(net238),
    .X(_1593_));
 sky130_fd_sc_hd__nor2_1 _2407_ (.A(net6),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__mux4_1 _2408_ (.A0(\mem[24][28] ),
    .A1(\mem[25][28] ),
    .A2(\mem[26][28] ),
    .A3(\mem[27][28] ),
    .S0(net320),
    .S1(net272),
    .X(_1595_));
 sky130_fd_sc_hd__mux2_1 _2409_ (.A0(\mem[30][28] ),
    .A1(\mem[31][28] ),
    .S(net320),
    .X(_1596_));
 sky130_fd_sc_hd__nand2_1 _2410_ (.A(net272),
    .B(_1596_),
    .Y(_1597_));
 sky130_fd_sc_hd__mux2_1 _2411_ (.A0(\mem[28][28] ),
    .A1(\mem[29][28] ),
    .S(net320),
    .X(_1598_));
 sky130_fd_sc_hd__nand2b_1 _2412_ (.A_N(net272),
    .B(_1598_),
    .Y(_1599_));
 sky130_fd_sc_hd__o21ai_1 _2413_ (.A1(net241),
    .A2(_1595_),
    .B1(net235),
    .Y(_1600_));
 sky130_fd_sc_hd__a31o_1 _2414_ (.A1(net241),
    .A2(_1597_),
    .A3(_1599_),
    .B1(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__mux4_1 _2415_ (.A0(\mem[20][28] ),
    .A1(\mem[21][28] ),
    .A2(\mem[22][28] ),
    .A3(\mem[23][28] ),
    .S0(net319),
    .S1(net271),
    .X(_1602_));
 sky130_fd_sc_hd__nor2_1 _2416_ (.A(net222),
    .B(_1602_),
    .Y(_1603_));
 sky130_fd_sc_hd__mux2_1 _2417_ (.A0(\mem[16][28] ),
    .A1(\mem[17][28] ),
    .S(net319),
    .X(_1604_));
 sky130_fd_sc_hd__nand2b_1 _2418_ (.A_N(net271),
    .B(_1604_),
    .Y(_1605_));
 sky130_fd_sc_hd__mux2_1 _2419_ (.A0(\mem[18][28] ),
    .A1(\mem[19][28] ),
    .S(net319),
    .X(_1606_));
 sky130_fd_sc_hd__nand2_1 _2420_ (.A(net271),
    .B(_1606_),
    .Y(_1607_));
 sky130_fd_sc_hd__a311o_1 _2421_ (.A1(net220),
    .A2(_1605_),
    .A3(_1607_),
    .B1(_1603_),
    .C1(net235),
    .X(_1608_));
 sky130_fd_sc_hd__a311oi_2 _2422_ (.A1(net230),
    .A2(_1601_),
    .A3(_1608_),
    .B1(net218),
    .C1(_1594_),
    .Y(net63));
 sky130_fd_sc_hd__mux4_1 _2423_ (.A0(\mem[0][29] ),
    .A1(\mem[1][29] ),
    .A2(\mem[2][29] ),
    .A3(\mem[3][29] ),
    .S0(net338),
    .S1(net286),
    .X(_1609_));
 sky130_fd_sc_hd__mux4_1 _2424_ (.A0(\mem[4][29] ),
    .A1(\mem[5][29] ),
    .A2(\mem[6][29] ),
    .A3(\mem[7][29] ),
    .S0(net334),
    .S1(net287),
    .X(_1610_));
 sky130_fd_sc_hd__mux4_1 _2425_ (.A0(\mem[12][29] ),
    .A1(\mem[13][29] ),
    .A2(\mem[14][29] ),
    .A3(\mem[15][29] ),
    .S0(net338),
    .S1(net287),
    .X(_1611_));
 sky130_fd_sc_hd__mux4_1 _2426_ (.A0(\mem[8][29] ),
    .A1(\mem[9][29] ),
    .A2(\mem[10][29] ),
    .A3(\mem[11][29] ),
    .S0(net334),
    .S1(net287),
    .X(_1612_));
 sky130_fd_sc_hd__mux4_2 _2427_ (.A0(_1609_),
    .A1(_1610_),
    .A2(_1612_),
    .A3(_1611_),
    .S0(net245),
    .S1(net238),
    .X(_1613_));
 sky130_fd_sc_hd__nor2_2 _2428_ (.A(net229),
    .B(_1613_),
    .Y(_1614_));
 sky130_fd_sc_hd__mux4_1 _2429_ (.A0(\mem[24][29] ),
    .A1(\mem[25][29] ),
    .A2(\mem[26][29] ),
    .A3(\mem[27][29] ),
    .S0(net318),
    .S1(net270),
    .X(_1615_));
 sky130_fd_sc_hd__mux2_1 _2430_ (.A0(\mem[30][29] ),
    .A1(\mem[31][29] ),
    .S(net318),
    .X(_1616_));
 sky130_fd_sc_hd__nand2_1 _2431_ (.A(net273),
    .B(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__mux2_1 _2432_ (.A0(\mem[28][29] ),
    .A1(\mem[29][29] ),
    .S(net321),
    .X(_1618_));
 sky130_fd_sc_hd__nand2b_1 _2433_ (.A_N(net273),
    .B(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__o21ai_1 _2434_ (.A1(net241),
    .A2(_1615_),
    .B1(net234),
    .Y(_1620_));
 sky130_fd_sc_hd__a31o_1 _2435_ (.A1(net241),
    .A2(_1617_),
    .A3(_1619_),
    .B1(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__mux4_1 _2436_ (.A0(\mem[20][29] ),
    .A1(\mem[21][29] ),
    .A2(\mem[22][29] ),
    .A3(\mem[23][29] ),
    .S0(net320),
    .S1(net272),
    .X(_1622_));
 sky130_fd_sc_hd__nor2_1 _2437_ (.A(net220),
    .B(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__mux2_1 _2438_ (.A0(\mem[16][29] ),
    .A1(\mem[17][29] ),
    .S(net321),
    .X(_1624_));
 sky130_fd_sc_hd__nand2b_1 _2439_ (.A_N(net273),
    .B(_1624_),
    .Y(_1625_));
 sky130_fd_sc_hd__mux2_1 _2440_ (.A0(\mem[18][29] ),
    .A1(\mem[19][29] ),
    .S(net321),
    .X(_1626_));
 sky130_fd_sc_hd__nand2_1 _2441_ (.A(net273),
    .B(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__a311o_1 _2442_ (.A1(net220),
    .A2(_1625_),
    .A3(_1627_),
    .B1(_1623_),
    .C1(net234),
    .X(_1628_));
 sky130_fd_sc_hd__a311oi_4 _2443_ (.A1(net230),
    .A2(_1621_),
    .A3(_1628_),
    .B1(net218),
    .C1(_1614_),
    .Y(net64));
 sky130_fd_sc_hd__mux4_1 _2444_ (.A0(\mem[0][30] ),
    .A1(\mem[1][30] ),
    .A2(\mem[2][30] ),
    .A3(\mem[3][30] ),
    .S0(net338),
    .S1(net290),
    .X(_1629_));
 sky130_fd_sc_hd__mux4_1 _2445_ (.A0(\mem[4][30] ),
    .A1(\mem[5][30] ),
    .A2(\mem[6][30] ),
    .A3(\mem[7][30] ),
    .S0(net335),
    .S1(net286),
    .X(_1630_));
 sky130_fd_sc_hd__mux4_1 _2446_ (.A0(\mem[12][30] ),
    .A1(\mem[13][30] ),
    .A2(\mem[14][30] ),
    .A3(\mem[15][30] ),
    .S0(net334),
    .S1(net287),
    .X(_1631_));
 sky130_fd_sc_hd__mux4_1 _2447_ (.A0(\mem[8][30] ),
    .A1(\mem[9][30] ),
    .A2(\mem[10][30] ),
    .A3(\mem[11][30] ),
    .S0(net334),
    .S1(net287),
    .X(_1632_));
 sky130_fd_sc_hd__mux4_1 _2448_ (.A0(_1629_),
    .A1(_1630_),
    .A2(_1632_),
    .A3(_1631_),
    .S0(net245),
    .S1(net238),
    .X(_1633_));
 sky130_fd_sc_hd__nor2_2 _2449_ (.A(net229),
    .B(_1633_),
    .Y(_1634_));
 sky130_fd_sc_hd__mux4_1 _2450_ (.A0(\mem[24][30] ),
    .A1(\mem[25][30] ),
    .A2(\mem[26][30] ),
    .A3(\mem[27][30] ),
    .S0(net321),
    .S1(net273),
    .X(_1635_));
 sky130_fd_sc_hd__mux2_1 _2451_ (.A0(\mem[30][30] ),
    .A1(\mem[31][30] ),
    .S(net321),
    .X(_1636_));
 sky130_fd_sc_hd__nand2_1 _2452_ (.A(net273),
    .B(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__mux2_1 _2453_ (.A0(\mem[28][30] ),
    .A1(\mem[29][30] ),
    .S(net321),
    .X(_1638_));
 sky130_fd_sc_hd__nand2b_1 _2454_ (.A_N(net273),
    .B(_1638_),
    .Y(_1639_));
 sky130_fd_sc_hd__o21ai_1 _2455_ (.A1(net241),
    .A2(_1635_),
    .B1(net234),
    .Y(_1640_));
 sky130_fd_sc_hd__a31o_1 _2456_ (.A1(net241),
    .A2(_1637_),
    .A3(_1639_),
    .B1(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__mux4_1 _2457_ (.A0(\mem[20][30] ),
    .A1(\mem[21][30] ),
    .A2(\mem[22][30] ),
    .A3(\mem[23][30] ),
    .S0(net319),
    .S1(net271),
    .X(_1642_));
 sky130_fd_sc_hd__nor2_1 _2458_ (.A(net220),
    .B(_1642_),
    .Y(_1643_));
 sky130_fd_sc_hd__mux2_1 _2459_ (.A0(\mem[16][30] ),
    .A1(\mem[17][30] ),
    .S(net319),
    .X(_1644_));
 sky130_fd_sc_hd__nand2b_1 _2460_ (.A_N(net271),
    .B(_1644_),
    .Y(_1645_));
 sky130_fd_sc_hd__mux2_1 _2461_ (.A0(\mem[18][30] ),
    .A1(\mem[19][30] ),
    .S(net319),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_1 _2462_ (.A(net271),
    .B(_1646_),
    .Y(_1647_));
 sky130_fd_sc_hd__a311o_1 _2463_ (.A1(net220),
    .A2(_1645_),
    .A3(_1647_),
    .B1(_1643_),
    .C1(net234),
    .X(_1648_));
 sky130_fd_sc_hd__a311oi_4 _2464_ (.A1(net230),
    .A2(_1641_),
    .A3(_1648_),
    .B1(net218),
    .C1(_1634_),
    .Y(net66));
 sky130_fd_sc_hd__mux4_1 _2465_ (.A0(\mem[0][31] ),
    .A1(\mem[1][31] ),
    .A2(\mem[2][31] ),
    .A3(\mem[3][31] ),
    .S0(net342),
    .S1(net294),
    .X(_1649_));
 sky130_fd_sc_hd__mux4_1 _2466_ (.A0(\mem[4][31] ),
    .A1(\mem[5][31] ),
    .A2(\mem[6][31] ),
    .A3(\mem[7][31] ),
    .S0(net343),
    .S1(net295),
    .X(_1650_));
 sky130_fd_sc_hd__mux4_1 _2467_ (.A0(\mem[12][31] ),
    .A1(\mem[13][31] ),
    .A2(\mem[14][31] ),
    .A3(\mem[15][31] ),
    .S0(net342),
    .S1(net294),
    .X(_1651_));
 sky130_fd_sc_hd__mux4_1 _2468_ (.A0(\mem[8][31] ),
    .A1(\mem[9][31] ),
    .A2(\mem[10][31] ),
    .A3(\mem[11][31] ),
    .S0(net342),
    .S1(net294),
    .X(_1652_));
 sky130_fd_sc_hd__mux4_1 _2469_ (.A0(_1649_),
    .A1(_1650_),
    .A2(_1652_),
    .A3(_1651_),
    .S0(net248),
    .S1(net240),
    .X(_1653_));
 sky130_fd_sc_hd__nor2_1 _2470_ (.A(net232),
    .B(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__mux4_1 _2471_ (.A0(\mem[24][31] ),
    .A1(\mem[25][31] ),
    .A2(\mem[26][31] ),
    .A3(\mem[27][31] ),
    .S0(net329),
    .S1(net282),
    .X(_1655_));
 sky130_fd_sc_hd__mux2_1 _2472_ (.A0(\mem[30][31] ),
    .A1(\mem[31][31] ),
    .S(net329),
    .X(_1656_));
 sky130_fd_sc_hd__nand2_1 _2473_ (.A(net282),
    .B(_1656_),
    .Y(_1657_));
 sky130_fd_sc_hd__mux2_1 _2474_ (.A0(\mem[28][31] ),
    .A1(\mem[29][31] ),
    .S(net329),
    .X(_1658_));
 sky130_fd_sc_hd__nand2b_1 _2475_ (.A_N(net282),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__o21ai_1 _2476_ (.A1(net243),
    .A2(_1655_),
    .B1(net236),
    .Y(_1660_));
 sky130_fd_sc_hd__a31o_1 _2477_ (.A1(net247),
    .A2(_1657_),
    .A3(_1659_),
    .B1(_1660_),
    .X(_1661_));
 sky130_fd_sc_hd__mux4_1 _2478_ (.A0(\mem[20][31] ),
    .A1(\mem[21][31] ),
    .A2(\mem[22][31] ),
    .A3(\mem[23][31] ),
    .S0(net327),
    .S1(net279),
    .X(_1662_));
 sky130_fd_sc_hd__nor2_1 _2479_ (.A(net224),
    .B(_1662_),
    .Y(_1663_));
 sky130_fd_sc_hd__mux2_1 _2480_ (.A0(\mem[16][31] ),
    .A1(\mem[17][31] ),
    .S(net330),
    .X(_1664_));
 sky130_fd_sc_hd__nand2b_1 _2481_ (.A_N(net281),
    .B(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__mux2_1 _2482_ (.A0(\mem[18][31] ),
    .A1(\mem[19][31] ),
    .S(net330),
    .X(_1666_));
 sky130_fd_sc_hd__nand2_1 _2483_ (.A(net281),
    .B(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__a311o_2 _2484_ (.A1(net224),
    .A2(_1665_),
    .A3(_1667_),
    .B1(_1663_),
    .C1(net236),
    .X(_1668_));
 sky130_fd_sc_hd__a311oi_4 _2485_ (.A1(net232),
    .A2(_1661_),
    .A3(_1668_),
    .B1(net219),
    .C1(_1654_),
    .Y(net67));
 sky130_fd_sc_hd__and3b_1 _2486_ (.A_N(net369),
    .B(net7),
    .C(net40),
    .X(_0573_));
 sky130_fd_sc_hd__and4b_2 _2487_ (.A_N(net369),
    .B(net41),
    .C(net7),
    .D(net40),
    .X(_1669_));
 sky130_fd_sc_hd__and3b_4 _2488_ (.A_N(net292),
    .B(net340),
    .C(net216),
    .X(_1670_));
 sky130_fd_sc_hd__and4b_1 _2489_ (.A_N(net283),
    .B(net331),
    .C(_1028_),
    .D(net217),
    .X(_1671_));
 sky130_fd_sc_hd__nand2_1 _2490_ (.A(_1028_),
    .B(_1670_),
    .Y(_1672_));
 sky130_fd_sc_hd__nor2_1 _2491_ (.A(net365),
    .B(net215),
    .Y(_1673_));
 sky130_fd_sc_hd__or2_2 _2492_ (.A(net365),
    .B(net215),
    .X(_1674_));
 sky130_fd_sc_hd__o22a_1 _2493_ (.A1(net228),
    .A2(_1672_),
    .B1(_1674_),
    .B2(net476),
    .X(_0541_));
 sky130_fd_sc_hd__o22a_1 _2494_ (.A1(net345),
    .A2(_1672_),
    .B1(_1674_),
    .B2(net388),
    .X(_0542_));
 sky130_fd_sc_hd__a22o_1 _2495_ (.A1(net268),
    .A2(net214),
    .B1(net150),
    .B2(net618),
    .X(_0543_));
 sky130_fd_sc_hd__a22o_1 _2496_ (.A1(net263),
    .A2(net215),
    .B1(net151),
    .B2(net874),
    .X(_0544_));
 sky130_fd_sc_hd__o22a_1 _2497_ (.A1(net260),
    .A2(_1672_),
    .B1(_1674_),
    .B2(net448),
    .X(_0545_));
 sky130_fd_sc_hd__o22a_1 _2498_ (.A1(net257),
    .A2(_1672_),
    .B1(_1674_),
    .B2(net528),
    .X(_0546_));
 sky130_fd_sc_hd__a22o_1 _2499_ (.A1(net255),
    .A2(net215),
    .B1(net151),
    .B2(net1428),
    .X(_0547_));
 sky130_fd_sc_hd__a22o_1 _2500_ (.A1(net253),
    .A2(net214),
    .B1(net150),
    .B2(net1330),
    .X(_0548_));
 sky130_fd_sc_hd__a22o_1 _2501_ (.A1(net251),
    .A2(net214),
    .B1(net151),
    .B2(net2394),
    .X(_0549_));
 sky130_fd_sc_hd__a22o_1 _2502_ (.A1(net249),
    .A2(net214),
    .B1(net150),
    .B2(net1284),
    .X(_0550_));
 sky130_fd_sc_hd__a22o_1 _2503_ (.A1(net225),
    .A2(net215),
    .B1(net151),
    .B2(net614),
    .X(_0551_));
 sky130_fd_sc_hd__a22o_1 _2504_ (.A1(net363),
    .A2(net214),
    .B1(net150),
    .B2(net1638),
    .X(_0552_));
 sky130_fd_sc_hd__a22o_1 _2505_ (.A1(net361),
    .A2(net215),
    .B1(net151),
    .B2(net1660),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_1 _2506_ (.A1(net359),
    .A2(net214),
    .B1(net150),
    .B2(net2396),
    .X(_0554_));
 sky130_fd_sc_hd__a22o_1 _2507_ (.A1(net357),
    .A2(net215),
    .B1(net151),
    .B2(net1450),
    .X(_0555_));
 sky130_fd_sc_hd__a22o_1 _2508_ (.A1(net355),
    .A2(net214),
    .B1(net150),
    .B2(net2086),
    .X(_0556_));
 sky130_fd_sc_hd__a22o_1 _2509_ (.A1(net353),
    .A2(net215),
    .B1(net151),
    .B2(net2220),
    .X(_0557_));
 sky130_fd_sc_hd__a22o_1 _2510_ (.A1(net351),
    .A2(net215),
    .B1(net151),
    .B2(net766),
    .X(_0558_));
 sky130_fd_sc_hd__a22o_1 _2511_ (.A1(net349),
    .A2(net214),
    .B1(net150),
    .B2(net1866),
    .X(_0559_));
 sky130_fd_sc_hd__a22o_1 _2512_ (.A1(net347),
    .A2(net215),
    .B1(net151),
    .B2(net1664),
    .X(_0560_));
 sky130_fd_sc_hd__a22o_1 _2513_ (.A1(net316),
    .A2(net215),
    .B1(net151),
    .B2(net2326),
    .X(_0561_));
 sky130_fd_sc_hd__a22o_1 _2514_ (.A1(net314),
    .A2(net214),
    .B1(net150),
    .B2(net938),
    .X(_0562_));
 sky130_fd_sc_hd__a22o_1 _2515_ (.A1(net312),
    .A2(net214),
    .B1(net150),
    .B2(net2006),
    .X(_0563_));
 sky130_fd_sc_hd__a22o_1 _2516_ (.A1(net310),
    .A2(net215),
    .B1(net150),
    .B2(net984),
    .X(_0564_));
 sky130_fd_sc_hd__a22o_1 _2517_ (.A1(net308),
    .A2(net214),
    .B1(net150),
    .B2(net2116),
    .X(_0565_));
 sky130_fd_sc_hd__a22o_1 _2518_ (.A1(net306),
    .A2(net214),
    .B1(net150),
    .B2(net1558),
    .X(_0566_));
 sky130_fd_sc_hd__a22o_1 _2519_ (.A1(net305),
    .A2(net214),
    .B1(net150),
    .B2(net858),
    .X(_0567_));
 sky130_fd_sc_hd__a22o_1 _2520_ (.A1(net301),
    .A2(net215),
    .B1(net151),
    .B2(net678),
    .X(_0568_));
 sky130_fd_sc_hd__a22o_1 _2521_ (.A1(net299),
    .A2(net214),
    .B1(net150),
    .B2(net912),
    .X(_0569_));
 sky130_fd_sc_hd__a22o_1 _2522_ (.A1(net297),
    .A2(net214),
    .B1(net150),
    .B2(net842),
    .X(_0570_));
 sky130_fd_sc_hd__a22o_1 _2523_ (.A1(net266),
    .A2(net214),
    .B1(net150),
    .B2(net1502),
    .X(_0571_));
 sky130_fd_sc_hd__a22o_1 _2524_ (.A1(net265),
    .A2(net215),
    .B1(net151),
    .B2(net1072),
    .X(_0572_));
 sky130_fd_sc_hd__and2b_2 _2525_ (.A_N(net332),
    .B(net284),
    .X(_1675_));
 sky130_fd_sc_hd__and2_4 _2526_ (.A(net216),
    .B(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__and3_1 _2527_ (.A(_1028_),
    .B(net217),
    .C(_1675_),
    .X(_1677_));
 sky130_fd_sc_hd__nand2_1 _2528_ (.A(_1028_),
    .B(_1676_),
    .Y(_1678_));
 sky130_fd_sc_hd__nor2_1 _2529_ (.A(net367),
    .B(net213),
    .Y(_1679_));
 sky130_fd_sc_hd__or2_2 _2530_ (.A(net365),
    .B(net213),
    .X(_1680_));
 sky130_fd_sc_hd__o22a_1 _2531_ (.A1(net228),
    .A2(_1678_),
    .B1(_1680_),
    .B2(net566),
    .X(_0574_));
 sky130_fd_sc_hd__o22a_1 _2532_ (.A1(net345),
    .A2(_1678_),
    .B1(_1680_),
    .B2(net442),
    .X(_0575_));
 sky130_fd_sc_hd__a22o_1 _2533_ (.A1(net268),
    .A2(net212),
    .B1(net148),
    .B2(net856),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _2534_ (.A1(net263),
    .A2(net213),
    .B1(net149),
    .B2(net1874),
    .X(_0577_));
 sky130_fd_sc_hd__o22a_1 _2535_ (.A1(net260),
    .A2(_1678_),
    .B1(_1680_),
    .B2(net586),
    .X(_0578_));
 sky130_fd_sc_hd__o22a_1 _2536_ (.A1(net257),
    .A2(_1678_),
    .B1(_1680_),
    .B2(net896),
    .X(_0579_));
 sky130_fd_sc_hd__a22o_1 _2537_ (.A1(net255),
    .A2(net213),
    .B1(net149),
    .B2(net852),
    .X(_0580_));
 sky130_fd_sc_hd__a22o_1 _2538_ (.A1(net253),
    .A2(net212),
    .B1(net148),
    .B2(net1460),
    .X(_0581_));
 sky130_fd_sc_hd__a22o_1 _2539_ (.A1(net251),
    .A2(net213),
    .B1(net148),
    .B2(net2304),
    .X(_0582_));
 sky130_fd_sc_hd__a22o_1 _2540_ (.A1(net249),
    .A2(net212),
    .B1(net148),
    .B2(net1626),
    .X(_0583_));
 sky130_fd_sc_hd__a22o_1 _2541_ (.A1(net225),
    .A2(net213),
    .B1(net149),
    .B2(net1180),
    .X(_0584_));
 sky130_fd_sc_hd__a22o_1 _2542_ (.A1(net363),
    .A2(net212),
    .B1(net148),
    .B2(net1134),
    .X(_0585_));
 sky130_fd_sc_hd__a22o_1 _2543_ (.A1(net361),
    .A2(net213),
    .B1(net149),
    .B2(net1742),
    .X(_0586_));
 sky130_fd_sc_hd__a22o_1 _2544_ (.A1(net359),
    .A2(net212),
    .B1(net148),
    .B2(net2180),
    .X(_0587_));
 sky130_fd_sc_hd__a22o_1 _2545_ (.A1(net357),
    .A2(net213),
    .B1(net149),
    .B2(net1930),
    .X(_0588_));
 sky130_fd_sc_hd__a22o_1 _2546_ (.A1(net355),
    .A2(net212),
    .B1(net148),
    .B2(net1602),
    .X(_0589_));
 sky130_fd_sc_hd__a22o_1 _2547_ (.A1(net353),
    .A2(net213),
    .B1(net149),
    .B2(net1256),
    .X(_0590_));
 sky130_fd_sc_hd__a22o_1 _2548_ (.A1(net351),
    .A2(net213),
    .B1(net149),
    .B2(net1498),
    .X(_0591_));
 sky130_fd_sc_hd__a22o_1 _2549_ (.A1(net349),
    .A2(net212),
    .B1(net149),
    .B2(net1598),
    .X(_0592_));
 sky130_fd_sc_hd__a22o_1 _2550_ (.A1(net347),
    .A2(net213),
    .B1(net149),
    .B2(net2094),
    .X(_0593_));
 sky130_fd_sc_hd__a22o_1 _2551_ (.A1(net316),
    .A2(net213),
    .B1(net149),
    .B2(net1954),
    .X(_0594_));
 sky130_fd_sc_hd__a22o_1 _2552_ (.A1(net314),
    .A2(net212),
    .B1(net148),
    .B2(net2248),
    .X(_0595_));
 sky130_fd_sc_hd__a22o_1 _2553_ (.A1(net312),
    .A2(net212),
    .B1(net148),
    .B2(net1746),
    .X(_0596_));
 sky130_fd_sc_hd__a22o_1 _2554_ (.A1(net310),
    .A2(net212),
    .B1(net148),
    .B2(net1222),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _2555_ (.A1(net308),
    .A2(net212),
    .B1(net148),
    .B2(net646),
    .X(_0598_));
 sky130_fd_sc_hd__a22o_1 _2556_ (.A1(net306),
    .A2(net212),
    .B1(net148),
    .B2(net2110),
    .X(_0599_));
 sky130_fd_sc_hd__a22o_1 _2557_ (.A1(net305),
    .A2(net212),
    .B1(net148),
    .B2(net1802),
    .X(_0600_));
 sky130_fd_sc_hd__a22o_1 _2558_ (.A1(net301),
    .A2(net213),
    .B1(net149),
    .B2(net1524),
    .X(_0601_));
 sky130_fd_sc_hd__a22o_1 _2559_ (.A1(net299),
    .A2(net212),
    .B1(net148),
    .B2(net2198),
    .X(_0602_));
 sky130_fd_sc_hd__a22o_1 _2560_ (.A1(net297),
    .A2(net212),
    .B1(net148),
    .B2(net1872),
    .X(_0603_));
 sky130_fd_sc_hd__a22o_1 _2561_ (.A1(net266),
    .A2(net212),
    .B1(net148),
    .B2(net900),
    .X(_0604_));
 sky130_fd_sc_hd__a22o_1 _2562_ (.A1(net265),
    .A2(net213),
    .B1(net149),
    .B2(net1582),
    .X(_0605_));
 sky130_fd_sc_hd__and3_2 _2563_ (.A(net231),
    .B(net237),
    .C(net244),
    .X(_1681_));
 sky130_fd_sc_hd__and3_2 _2564_ (.A(net217),
    .B(_1675_),
    .C(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__nand2_2 _2565_ (.A(_1676_),
    .B(_1681_),
    .Y(_1683_));
 sky130_fd_sc_hd__nor2_1 _2566_ (.A(net367),
    .B(net210),
    .Y(_1684_));
 sky130_fd_sc_hd__or2_2 _2567_ (.A(net366),
    .B(net211),
    .X(_1685_));
 sky130_fd_sc_hd__o22a_1 _2568_ (.A1(net227),
    .A2(_1683_),
    .B1(_1685_),
    .B2(net444),
    .X(_0606_));
 sky130_fd_sc_hd__o22a_1 _2569_ (.A1(net345),
    .A2(_1683_),
    .B1(_1685_),
    .B2(net452),
    .X(_0607_));
 sky130_fd_sc_hd__a22o_1 _2570_ (.A1(net268),
    .A2(net210),
    .B1(net146),
    .B2(net708),
    .X(_0608_));
 sky130_fd_sc_hd__a22o_1 _2571_ (.A1(net261),
    .A2(net211),
    .B1(net146),
    .B2(net2078),
    .X(_0609_));
 sky130_fd_sc_hd__o22a_1 _2572_ (.A1(net260),
    .A2(_1683_),
    .B1(_1685_),
    .B2(net416),
    .X(_0610_));
 sky130_fd_sc_hd__o22a_1 _2573_ (.A1(net257),
    .A2(_1683_),
    .B1(_1685_),
    .B2(net468),
    .X(_0611_));
 sky130_fd_sc_hd__a22o_1 _2574_ (.A1(net255),
    .A2(net211),
    .B1(net147),
    .B2(net732),
    .X(_0612_));
 sky130_fd_sc_hd__a22o_1 _2575_ (.A1(net253),
    .A2(net210),
    .B1(net146),
    .B2(net1332),
    .X(_0613_));
 sky130_fd_sc_hd__a22o_1 _2576_ (.A1(net251),
    .A2(net211),
    .B1(net147),
    .B2(net2352),
    .X(_0614_));
 sky130_fd_sc_hd__a22o_1 _2577_ (.A1(net249),
    .A2(net210),
    .B1(net146),
    .B2(net1652),
    .X(_0615_));
 sky130_fd_sc_hd__a22o_1 _2578_ (.A1(net225),
    .A2(net211),
    .B1(net147),
    .B2(net1296),
    .X(_0616_));
 sky130_fd_sc_hd__a22o_1 _2579_ (.A1(net363),
    .A2(net210),
    .B1(net146),
    .B2(net1454),
    .X(_0617_));
 sky130_fd_sc_hd__a22o_1 _2580_ (.A1(net361),
    .A2(net211),
    .B1(net147),
    .B2(net2138),
    .X(_0618_));
 sky130_fd_sc_hd__a22o_1 _2581_ (.A1(net359),
    .A2(net210),
    .B1(net146),
    .B2(net1970),
    .X(_0619_));
 sky130_fd_sc_hd__a22o_1 _2582_ (.A1(net357),
    .A2(net211),
    .B1(net147),
    .B2(net1302),
    .X(_0620_));
 sky130_fd_sc_hd__a22o_1 _2583_ (.A1(net355),
    .A2(net211),
    .B1(net147),
    .B2(net2278),
    .X(_0621_));
 sky130_fd_sc_hd__a22o_1 _2584_ (.A1(net353),
    .A2(net211),
    .B1(net147),
    .B2(net1796),
    .X(_0622_));
 sky130_fd_sc_hd__a22o_1 _2585_ (.A1(net351),
    .A2(net211),
    .B1(net147),
    .B2(net1020),
    .X(_0623_));
 sky130_fd_sc_hd__a22o_1 _2586_ (.A1(net349),
    .A2(net210),
    .B1(net146),
    .B2(net1690),
    .X(_0624_));
 sky130_fd_sc_hd__a22o_1 _2587_ (.A1(net347),
    .A2(net211),
    .B1(net147),
    .B2(net1042),
    .X(_0625_));
 sky130_fd_sc_hd__a22o_1 _2588_ (.A1(net316),
    .A2(net211),
    .B1(net147),
    .B2(net1376),
    .X(_0626_));
 sky130_fd_sc_hd__a22o_1 _2589_ (.A1(net314),
    .A2(net210),
    .B1(net146),
    .B2(net1448),
    .X(_0627_));
 sky130_fd_sc_hd__a22o_1 _2590_ (.A1(net312),
    .A2(net210),
    .B1(net146),
    .B2(net1772),
    .X(_0628_));
 sky130_fd_sc_hd__a22o_1 _2591_ (.A1(net310),
    .A2(net210),
    .B1(net146),
    .B2(net680),
    .X(_0629_));
 sky130_fd_sc_hd__a22o_1 _2592_ (.A1(net308),
    .A2(net210),
    .B1(net146),
    .B2(net2000),
    .X(_0630_));
 sky130_fd_sc_hd__a22o_1 _2593_ (.A1(net306),
    .A2(net210),
    .B1(net146),
    .B2(net1128),
    .X(_0631_));
 sky130_fd_sc_hd__a22o_1 _2594_ (.A1(net304),
    .A2(net210),
    .B1(net146),
    .B2(net752),
    .X(_0632_));
 sky130_fd_sc_hd__a22o_1 _2595_ (.A1(net301),
    .A2(net211),
    .B1(net147),
    .B2(net1682),
    .X(_0633_));
 sky130_fd_sc_hd__a22o_1 _2596_ (.A1(net299),
    .A2(net210),
    .B1(net146),
    .B2(net2060),
    .X(_0634_));
 sky130_fd_sc_hd__a22o_1 _2597_ (.A1(net297),
    .A2(net210),
    .B1(net146),
    .B2(net968),
    .X(_0635_));
 sky130_fd_sc_hd__a22o_1 _2598_ (.A1(net266),
    .A2(net210),
    .B1(net146),
    .B2(net1560),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_1 _2599_ (.A1(net264),
    .A2(net211),
    .B1(net147),
    .B2(net610),
    .X(_0637_));
 sky130_fd_sc_hd__and3b_2 _2600_ (.A_N(net231),
    .B(net239),
    .C(net247),
    .X(_1686_));
 sky130_fd_sc_hd__and3_4 _2601_ (.A(net292),
    .B(net340),
    .C(net216),
    .X(_1687_));
 sky130_fd_sc_hd__and4_1 _2602_ (.A(net291),
    .B(net339),
    .C(net216),
    .D(_1686_),
    .X(_1688_));
 sky130_fd_sc_hd__nand2_2 _2603_ (.A(_1686_),
    .B(_1687_),
    .Y(_1689_));
 sky130_fd_sc_hd__nor2_1 _2604_ (.A(net368),
    .B(net208),
    .Y(_1690_));
 sky130_fd_sc_hd__or2_2 _2605_ (.A(net366),
    .B(net208),
    .X(_1691_));
 sky130_fd_sc_hd__o22a_1 _2606_ (.A1(net227),
    .A2(_1689_),
    .B1(_1691_),
    .B2(net480),
    .X(_0638_));
 sky130_fd_sc_hd__o22a_1 _2607_ (.A1(net346),
    .A2(_1689_),
    .B1(_1691_),
    .B2(net420),
    .X(_0639_));
 sky130_fd_sc_hd__a22o_1 _2608_ (.A1(net269),
    .A2(net209),
    .B1(net144),
    .B2(net1178),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_1 _2609_ (.A1(net261),
    .A2(net208),
    .B1(net145),
    .B2(net1362),
    .X(_0641_));
 sky130_fd_sc_hd__o22a_1 _2610_ (.A1(net259),
    .A2(_1689_),
    .B1(_1691_),
    .B2(net422),
    .X(_0642_));
 sky130_fd_sc_hd__o22a_1 _2611_ (.A1(net258),
    .A2(_1689_),
    .B1(_1691_),
    .B2(net626),
    .X(_0643_));
 sky130_fd_sc_hd__a22o_1 _2612_ (.A1(net256),
    .A2(net208),
    .B1(net145),
    .B2(net1352),
    .X(_0644_));
 sky130_fd_sc_hd__a22o_1 _2613_ (.A1(net254),
    .A2(net209),
    .B1(net144),
    .B2(net1646),
    .X(_0645_));
 sky130_fd_sc_hd__a22o_1 _2614_ (.A1(net252),
    .A2(net208),
    .B1(net144),
    .B2(net1140),
    .X(_0646_));
 sky130_fd_sc_hd__a22o_1 _2615_ (.A1(net250),
    .A2(net209),
    .B1(net144),
    .B2(net1654),
    .X(_0647_));
 sky130_fd_sc_hd__a22o_1 _2616_ (.A1(net226),
    .A2(net208),
    .B1(net145),
    .B2(net1234),
    .X(_0648_));
 sky130_fd_sc_hd__a22o_1 _2617_ (.A1(net364),
    .A2(net209),
    .B1(net144),
    .B2(net2324),
    .X(_0649_));
 sky130_fd_sc_hd__a22o_1 _2618_ (.A1(net362),
    .A2(net208),
    .B1(net145),
    .B2(net1118),
    .X(_0650_));
 sky130_fd_sc_hd__a22o_1 _2619_ (.A1(net360),
    .A2(net209),
    .B1(net144),
    .B2(net744),
    .X(_0651_));
 sky130_fd_sc_hd__a22o_1 _2620_ (.A1(net358),
    .A2(net208),
    .B1(net145),
    .B2(net2254),
    .X(_0652_));
 sky130_fd_sc_hd__a22o_1 _2621_ (.A1(net356),
    .A2(net208),
    .B1(net145),
    .B2(net2022),
    .X(_0653_));
 sky130_fd_sc_hd__a22o_1 _2622_ (.A1(net354),
    .A2(net209),
    .B1(net145),
    .B2(net1618),
    .X(_0654_));
 sky130_fd_sc_hd__a22o_1 _2623_ (.A1(net352),
    .A2(net208),
    .B1(net145),
    .B2(net918),
    .X(_0655_));
 sky130_fd_sc_hd__a22o_1 _2624_ (.A1(net350),
    .A2(net209),
    .B1(net144),
    .B2(net2136),
    .X(_0656_));
 sky130_fd_sc_hd__a22o_1 _2625_ (.A1(net348),
    .A2(net208),
    .B1(net145),
    .B2(net1310),
    .X(_0657_));
 sky130_fd_sc_hd__a22o_1 _2626_ (.A1(net317),
    .A2(net208),
    .B1(net145),
    .B2(net850),
    .X(_0658_));
 sky130_fd_sc_hd__a22o_1 _2627_ (.A1(net315),
    .A2(net208),
    .B1(net144),
    .B2(net1272),
    .X(_0659_));
 sky130_fd_sc_hd__a22o_1 _2628_ (.A1(net313),
    .A2(net209),
    .B1(net144),
    .B2(net2286),
    .X(_0660_));
 sky130_fd_sc_hd__a22o_1 _2629_ (.A1(net311),
    .A2(net209),
    .B1(net144),
    .B2(net828),
    .X(_0661_));
 sky130_fd_sc_hd__a22o_1 _2630_ (.A1(net309),
    .A2(net209),
    .B1(net144),
    .B2(net1410),
    .X(_0662_));
 sky130_fd_sc_hd__a22o_1 _2631_ (.A1(net307),
    .A2(net209),
    .B1(net144),
    .B2(net1278),
    .X(_0663_));
 sky130_fd_sc_hd__a22o_1 _2632_ (.A1(net303),
    .A2(net208),
    .B1(net144),
    .B2(net1324),
    .X(_0664_));
 sky130_fd_sc_hd__a22o_1 _2633_ (.A1(net302),
    .A2(net208),
    .B1(net145),
    .B2(net630),
    .X(_0665_));
 sky130_fd_sc_hd__a22o_1 _2634_ (.A1(net300),
    .A2(net209),
    .B1(net144),
    .B2(net1292),
    .X(_0666_));
 sky130_fd_sc_hd__a22o_1 _2635_ (.A1(net298),
    .A2(net209),
    .B1(net144),
    .B2(net1518),
    .X(_0667_));
 sky130_fd_sc_hd__a22o_1 _2636_ (.A1(net267),
    .A2(net209),
    .B1(net144),
    .B2(net992),
    .X(_0668_));
 sky130_fd_sc_hd__a22o_1 _2637_ (.A1(net264),
    .A2(net208),
    .B1(net145),
    .B2(net1000),
    .X(_0669_));
 sky130_fd_sc_hd__and3b_2 _2638_ (.A_N(net244),
    .B(net237),
    .C(net231),
    .X(_1692_));
 sky130_fd_sc_hd__nor2_4 _2639_ (.A(net282),
    .B(net329),
    .Y(_1693_));
 sky130_fd_sc_hd__and2_4 _2640_ (.A(net216),
    .B(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__and3_1 _2641_ (.A(net217),
    .B(_1692_),
    .C(_1693_),
    .X(_1695_));
 sky130_fd_sc_hd__nand2_2 _2642_ (.A(_1692_),
    .B(_1694_),
    .Y(_1696_));
 sky130_fd_sc_hd__nor2_1 _2643_ (.A(net365),
    .B(net206),
    .Y(_1697_));
 sky130_fd_sc_hd__or2_2 _2644_ (.A(net366),
    .B(net206),
    .X(_1698_));
 sky130_fd_sc_hd__o22a_1 _2645_ (.A1(net228),
    .A2(_1696_),
    .B1(_1698_),
    .B2(net542),
    .X(_0670_));
 sky130_fd_sc_hd__o22a_1 _2646_ (.A1(net345),
    .A2(_1696_),
    .B1(_1698_),
    .B2(net496),
    .X(_0671_));
 sky130_fd_sc_hd__a22o_1 _2647_ (.A1(net268),
    .A2(net207),
    .B1(net142),
    .B2(net1568),
    .X(_0672_));
 sky130_fd_sc_hd__a22o_1 _2648_ (.A1(net261),
    .A2(net206),
    .B1(net142),
    .B2(net2204),
    .X(_0673_));
 sky130_fd_sc_hd__o22a_1 _2649_ (.A1(net260),
    .A2(_1696_),
    .B1(_1698_),
    .B2(net484),
    .X(_0674_));
 sky130_fd_sc_hd__o22a_1 _2650_ (.A1(net257),
    .A2(_1696_),
    .B1(_1698_),
    .B2(net534),
    .X(_0675_));
 sky130_fd_sc_hd__a22o_1 _2651_ (.A1(net255),
    .A2(net206),
    .B1(net143),
    .B2(net650),
    .X(_0676_));
 sky130_fd_sc_hd__a22o_1 _2652_ (.A1(net253),
    .A2(net207),
    .B1(net142),
    .B2(net1246),
    .X(_0677_));
 sky130_fd_sc_hd__a22o_1 _2653_ (.A1(net251),
    .A2(net206),
    .B1(net142),
    .B2(net1504),
    .X(_0678_));
 sky130_fd_sc_hd__a22o_1 _2654_ (.A1(net249),
    .A2(net207),
    .B1(net142),
    .B2(net2002),
    .X(_0679_));
 sky130_fd_sc_hd__a22o_1 _2655_ (.A1(net225),
    .A2(net206),
    .B1(net143),
    .B2(net882),
    .X(_0680_));
 sky130_fd_sc_hd__a22o_1 _2656_ (.A1(net363),
    .A2(net207),
    .B1(net142),
    .B2(net1950),
    .X(_0681_));
 sky130_fd_sc_hd__a22o_1 _2657_ (.A1(net361),
    .A2(net207),
    .B1(net143),
    .B2(net2050),
    .X(_0682_));
 sky130_fd_sc_hd__a22o_1 _2658_ (.A1(net359),
    .A2(net206),
    .B1(net143),
    .B2(net1860),
    .X(_0683_));
 sky130_fd_sc_hd__a22o_1 _2659_ (.A1(net357),
    .A2(net206),
    .B1(net143),
    .B2(net1392),
    .X(_0684_));
 sky130_fd_sc_hd__a22o_1 _2660_ (.A1(net355),
    .A2(net206),
    .B1(net143),
    .B2(net2320),
    .X(_0685_));
 sky130_fd_sc_hd__a22o_1 _2661_ (.A1(net353),
    .A2(net206),
    .B1(net143),
    .B2(net1116),
    .X(_0686_));
 sky130_fd_sc_hd__a22o_1 _2662_ (.A1(net351),
    .A2(net206),
    .B1(net143),
    .B2(net1268),
    .X(_0687_));
 sky130_fd_sc_hd__a22o_1 _2663_ (.A1(net349),
    .A2(net207),
    .B1(net142),
    .B2(net2280),
    .X(_0688_));
 sky130_fd_sc_hd__a22o_1 _2664_ (.A1(net347),
    .A2(net206),
    .B1(net143),
    .B2(net1674),
    .X(_0689_));
 sky130_fd_sc_hd__a22o_1 _2665_ (.A1(net316),
    .A2(net206),
    .B1(net143),
    .B2(net588),
    .X(_0690_));
 sky130_fd_sc_hd__a22o_1 _2666_ (.A1(net314),
    .A2(net207),
    .B1(net142),
    .B2(net982),
    .X(_0691_));
 sky130_fd_sc_hd__a22o_1 _2667_ (.A1(net312),
    .A2(net207),
    .B1(net142),
    .B2(net1286),
    .X(_0692_));
 sky130_fd_sc_hd__a22o_1 _2668_ (.A1(net310),
    .A2(net207),
    .B1(net142),
    .B2(net640),
    .X(_0693_));
 sky130_fd_sc_hd__a22o_1 _2669_ (.A1(net308),
    .A2(net207),
    .B1(net142),
    .B2(net1642),
    .X(_0694_));
 sky130_fd_sc_hd__a22o_1 _2670_ (.A1(net306),
    .A2(net207),
    .B1(net142),
    .B2(net2106),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _2671_ (.A1(net304),
    .A2(net207),
    .B1(net142),
    .B2(net1710),
    .X(_0696_));
 sky130_fd_sc_hd__a22o_1 _2672_ (.A1(net301),
    .A2(net206),
    .B1(net143),
    .B2(net804),
    .X(_0697_));
 sky130_fd_sc_hd__a22o_1 _2673_ (.A1(net299),
    .A2(net206),
    .B1(net142),
    .B2(net1274),
    .X(_0698_));
 sky130_fd_sc_hd__a22o_1 _2674_ (.A1(net297),
    .A2(net207),
    .B1(net142),
    .B2(net1972),
    .X(_0699_));
 sky130_fd_sc_hd__a22o_1 _2675_ (.A1(net266),
    .A2(net207),
    .B1(net142),
    .B2(net622),
    .X(_0700_));
 sky130_fd_sc_hd__a22o_1 _2676_ (.A1(net264),
    .A2(net206),
    .B1(net143),
    .B2(net1316),
    .X(_0701_));
 sky130_fd_sc_hd__and4_2 _2677_ (.A(net284),
    .B(net332),
    .C(net217),
    .D(_1681_),
    .X(_1699_));
 sky130_fd_sc_hd__nand2_2 _2678_ (.A(_1681_),
    .B(_1687_),
    .Y(_1700_));
 sky130_fd_sc_hd__nor2_1 _2679_ (.A(net367),
    .B(net204),
    .Y(_1701_));
 sky130_fd_sc_hd__or2_2 _2680_ (.A(net366),
    .B(net205),
    .X(_1702_));
 sky130_fd_sc_hd__o22a_1 _2681_ (.A1(net227),
    .A2(_1700_),
    .B1(_1702_),
    .B2(net446),
    .X(_0702_));
 sky130_fd_sc_hd__o22a_1 _2682_ (.A1(net345),
    .A2(_1700_),
    .B1(_1702_),
    .B2(net636),
    .X(_0703_));
 sky130_fd_sc_hd__a22o_1 _2683_ (.A1(net268),
    .A2(net204),
    .B1(net140),
    .B2(net2404),
    .X(_0704_));
 sky130_fd_sc_hd__a22o_1 _2684_ (.A1(net261),
    .A2(net205),
    .B1(net140),
    .B2(net2380),
    .X(_0705_));
 sky130_fd_sc_hd__o22a_1 _2685_ (.A1(net259),
    .A2(_1700_),
    .B1(_1702_),
    .B2(net578),
    .X(_0706_));
 sky130_fd_sc_hd__o22a_1 _2686_ (.A1(net257),
    .A2(_1700_),
    .B1(_1702_),
    .B2(net490),
    .X(_0707_));
 sky130_fd_sc_hd__a22o_1 _2687_ (.A1(net255),
    .A2(net205),
    .B1(net141),
    .B2(net1594),
    .X(_0708_));
 sky130_fd_sc_hd__a22o_1 _2688_ (.A1(net253),
    .A2(net204),
    .B1(net140),
    .B2(net1656),
    .X(_0709_));
 sky130_fd_sc_hd__a22o_1 _2689_ (.A1(net251),
    .A2(net205),
    .B1(net141),
    .B2(net2308),
    .X(_0710_));
 sky130_fd_sc_hd__a22o_1 _2690_ (.A1(net249),
    .A2(net204),
    .B1(net140),
    .B2(net2032),
    .X(_0711_));
 sky130_fd_sc_hd__a22o_1 _2691_ (.A1(net225),
    .A2(net205),
    .B1(net141),
    .B2(net1824),
    .X(_0712_));
 sky130_fd_sc_hd__a22o_1 _2692_ (.A1(net363),
    .A2(net204),
    .B1(net140),
    .B2(net1994),
    .X(_0713_));
 sky130_fd_sc_hd__a22o_1 _2693_ (.A1(net361),
    .A2(net205),
    .B1(net141),
    .B2(net2126),
    .X(_0714_));
 sky130_fd_sc_hd__a22o_1 _2694_ (.A1(net359),
    .A2(net204),
    .B1(net140),
    .B2(net2342),
    .X(_0715_));
 sky130_fd_sc_hd__a22o_1 _2695_ (.A1(net357),
    .A2(net205),
    .B1(net141),
    .B2(net2370),
    .X(_0716_));
 sky130_fd_sc_hd__a22o_1 _2696_ (.A1(net355),
    .A2(net205),
    .B1(net141),
    .B2(net2328),
    .X(_0717_));
 sky130_fd_sc_hd__a22o_1 _2697_ (.A1(net353),
    .A2(net205),
    .B1(net141),
    .B2(net1306),
    .X(_0718_));
 sky130_fd_sc_hd__a22o_1 _2698_ (.A1(net351),
    .A2(net205),
    .B1(net141),
    .B2(net2252),
    .X(_0719_));
 sky130_fd_sc_hd__a22o_1 _2699_ (.A1(net349),
    .A2(net204),
    .B1(net140),
    .B2(net2150),
    .X(_0720_));
 sky130_fd_sc_hd__a22o_1 _2700_ (.A1(net347),
    .A2(net205),
    .B1(net141),
    .B2(net1702),
    .X(_0721_));
 sky130_fd_sc_hd__a22o_1 _2701_ (.A1(net316),
    .A2(net205),
    .B1(net141),
    .B2(net2350),
    .X(_0722_));
 sky130_fd_sc_hd__a22o_1 _2702_ (.A1(net314),
    .A2(net204),
    .B1(net140),
    .B2(net1774),
    .X(_0723_));
 sky130_fd_sc_hd__a22o_1 _2703_ (.A1(net312),
    .A2(net204),
    .B1(net140),
    .B2(net1550),
    .X(_0724_));
 sky130_fd_sc_hd__a22o_1 _2704_ (.A1(net310),
    .A2(net204),
    .B1(net140),
    .B2(net1778),
    .X(_0725_));
 sky130_fd_sc_hd__a22o_1 _2705_ (.A1(net308),
    .A2(net204),
    .B1(net140),
    .B2(net2186),
    .X(_0726_));
 sky130_fd_sc_hd__a22o_1 _2706_ (.A1(net306),
    .A2(net204),
    .B1(net140),
    .B2(net1692),
    .X(_0727_));
 sky130_fd_sc_hd__a22o_1 _2707_ (.A1(net304),
    .A2(net204),
    .B1(net140),
    .B2(net2100),
    .X(_0728_));
 sky130_fd_sc_hd__a22o_1 _2708_ (.A1(net301),
    .A2(net205),
    .B1(net141),
    .B2(net1298),
    .X(_0729_));
 sky130_fd_sc_hd__a22o_1 _2709_ (.A1(net299),
    .A2(net204),
    .B1(net140),
    .B2(net2160),
    .X(_0730_));
 sky130_fd_sc_hd__a22o_1 _2710_ (.A1(net297),
    .A2(net204),
    .B1(net140),
    .B2(net1986),
    .X(_0731_));
 sky130_fd_sc_hd__a22o_1 _2711_ (.A1(net266),
    .A2(net204),
    .B1(net140),
    .B2(net2386),
    .X(_0732_));
 sky130_fd_sc_hd__a22o_1 _2712_ (.A1(net264),
    .A2(net205),
    .B1(net141),
    .B2(net1920),
    .X(_0733_));
 sky130_fd_sc_hd__and4b_1 _2713_ (.A_N(net282),
    .B(net329),
    .C(net217),
    .D(_1692_),
    .X(_1703_));
 sky130_fd_sc_hd__nand2_1 _2714_ (.A(_1670_),
    .B(_1692_),
    .Y(_1704_));
 sky130_fd_sc_hd__nor2_1 _2715_ (.A(net365),
    .B(net202),
    .Y(_1705_));
 sky130_fd_sc_hd__or2_2 _2716_ (.A(net365),
    .B(net202),
    .X(_1706_));
 sky130_fd_sc_hd__o22a_1 _2717_ (.A1(net228),
    .A2(_1704_),
    .B1(_1706_),
    .B2(net424),
    .X(_0734_));
 sky130_fd_sc_hd__o22a_1 _2718_ (.A1(net345),
    .A2(_1704_),
    .B1(_1706_),
    .B2(net396),
    .X(_0735_));
 sky130_fd_sc_hd__a22o_1 _2719_ (.A1(net268),
    .A2(net203),
    .B1(net138),
    .B2(net794),
    .X(_0736_));
 sky130_fd_sc_hd__a22o_1 _2720_ (.A1(net261),
    .A2(net202),
    .B1(net138),
    .B2(net2218),
    .X(_0737_));
 sky130_fd_sc_hd__o22a_1 _2721_ (.A1(net260),
    .A2(_1704_),
    .B1(_1706_),
    .B2(net412),
    .X(_0738_));
 sky130_fd_sc_hd__o22a_1 _2722_ (.A1(net257),
    .A2(_1704_),
    .B1(_1706_),
    .B2(net402),
    .X(_0739_));
 sky130_fd_sc_hd__a22o_1 _2723_ (.A1(net255),
    .A2(net202),
    .B1(net139),
    .B2(net956),
    .X(_0740_));
 sky130_fd_sc_hd__a22o_1 _2724_ (.A1(net253),
    .A2(net203),
    .B1(net138),
    .B2(net1158),
    .X(_0741_));
 sky130_fd_sc_hd__a22o_1 _2725_ (.A1(net251),
    .A2(net202),
    .B1(net138),
    .B2(net2054),
    .X(_0742_));
 sky130_fd_sc_hd__a22o_1 _2726_ (.A1(net249),
    .A2(net203),
    .B1(net138),
    .B2(net1414),
    .X(_0743_));
 sky130_fd_sc_hd__a22o_1 _2727_ (.A1(net225),
    .A2(net202),
    .B1(net139),
    .B2(net1224),
    .X(_0744_));
 sky130_fd_sc_hd__a22o_1 _2728_ (.A1(net363),
    .A2(net203),
    .B1(net138),
    .B2(net1090),
    .X(_0745_));
 sky130_fd_sc_hd__a22o_1 _2729_ (.A1(net361),
    .A2(net203),
    .B1(net139),
    .B2(net1394),
    .X(_0746_));
 sky130_fd_sc_hd__a22o_1 _2730_ (.A1(net359),
    .A2(net202),
    .B1(net139),
    .B2(net2108),
    .X(_0747_));
 sky130_fd_sc_hd__a22o_1 _2731_ (.A1(net357),
    .A2(net202),
    .B1(net139),
    .B2(net2224),
    .X(_0748_));
 sky130_fd_sc_hd__a22o_1 _2732_ (.A1(net355),
    .A2(net202),
    .B1(net139),
    .B2(net1080),
    .X(_0749_));
 sky130_fd_sc_hd__a22o_1 _2733_ (.A1(net353),
    .A2(net202),
    .B1(net139),
    .B2(net2166),
    .X(_0750_));
 sky130_fd_sc_hd__a22o_1 _2734_ (.A1(net351),
    .A2(net202),
    .B1(net139),
    .B2(net928),
    .X(_0751_));
 sky130_fd_sc_hd__a22o_1 _2735_ (.A1(net349),
    .A2(net203),
    .B1(net138),
    .B2(net1942),
    .X(_0752_));
 sky130_fd_sc_hd__a22o_1 _2736_ (.A1(net347),
    .A2(net202),
    .B1(net139),
    .B2(net686),
    .X(_0753_));
 sky130_fd_sc_hd__a22o_1 _2737_ (.A1(net316),
    .A2(net202),
    .B1(net139),
    .B2(net1540),
    .X(_0754_));
 sky130_fd_sc_hd__a22o_1 _2738_ (.A1(net314),
    .A2(net203),
    .B1(net138),
    .B2(net700),
    .X(_0755_));
 sky130_fd_sc_hd__a22o_1 _2739_ (.A1(net312),
    .A2(net203),
    .B1(net138),
    .B2(net638),
    .X(_0756_));
 sky130_fd_sc_hd__a22o_1 _2740_ (.A1(net310),
    .A2(net203),
    .B1(net138),
    .B2(net1078),
    .X(_0757_));
 sky130_fd_sc_hd__a22o_1 _2741_ (.A1(net308),
    .A2(net203),
    .B1(net138),
    .B2(net1864),
    .X(_0758_));
 sky130_fd_sc_hd__a22o_1 _2742_ (.A1(net306),
    .A2(net203),
    .B1(net138),
    .B2(net1010),
    .X(_0759_));
 sky130_fd_sc_hd__a22o_1 _2743_ (.A1(net304),
    .A2(net203),
    .B1(net138),
    .B2(net1130),
    .X(_0760_));
 sky130_fd_sc_hd__a22o_1 _2744_ (.A1(net301),
    .A2(net202),
    .B1(net139),
    .B2(net2042),
    .X(_0761_));
 sky130_fd_sc_hd__a22o_1 _2745_ (.A1(net299),
    .A2(net202),
    .B1(net138),
    .B2(net2036),
    .X(_0762_));
 sky130_fd_sc_hd__a22o_1 _2746_ (.A1(net297),
    .A2(net203),
    .B1(net138),
    .B2(net1936),
    .X(_0763_));
 sky130_fd_sc_hd__a22o_1 _2747_ (.A1(net266),
    .A2(net203),
    .B1(net138),
    .B2(net1360),
    .X(_0764_));
 sky130_fd_sc_hd__a22o_1 _2748_ (.A1(net264),
    .A2(net202),
    .B1(net139),
    .B2(net1152),
    .X(_0765_));
 sky130_fd_sc_hd__and4_1 _2749_ (.A(net282),
    .B(net330),
    .C(net217),
    .D(_1692_),
    .X(_1707_));
 sky130_fd_sc_hd__nand2_1 _2750_ (.A(_1687_),
    .B(_1692_),
    .Y(_1708_));
 sky130_fd_sc_hd__nor2_1 _2751_ (.A(net365),
    .B(net201),
    .Y(_1709_));
 sky130_fd_sc_hd__or2_2 _2752_ (.A(net365),
    .B(net200),
    .X(_1710_));
 sky130_fd_sc_hd__o22a_1 _2753_ (.A1(net228),
    .A2(_1708_),
    .B1(_1710_),
    .B2(net532),
    .X(_0766_));
 sky130_fd_sc_hd__o22a_1 _2754_ (.A1(net345),
    .A2(_1708_),
    .B1(_1710_),
    .B2(net380),
    .X(_0767_));
 sky130_fd_sc_hd__a22o_1 _2755_ (.A1(net268),
    .A2(net200),
    .B1(net136),
    .B2(net916),
    .X(_0768_));
 sky130_fd_sc_hd__a22o_1 _2756_ (.A1(net261),
    .A2(net201),
    .B1(net136),
    .B2(net1974),
    .X(_0769_));
 sky130_fd_sc_hd__o22a_1 _2757_ (.A1(net260),
    .A2(_1708_),
    .B1(_1710_),
    .B2(net404),
    .X(_0770_));
 sky130_fd_sc_hd__o22a_1 _2758_ (.A1(net257),
    .A2(_1708_),
    .B1(_1710_),
    .B2(net576),
    .X(_0771_));
 sky130_fd_sc_hd__a22o_1 _2759_ (.A1(net255),
    .A2(net201),
    .B1(net137),
    .B2(net806),
    .X(_0772_));
 sky130_fd_sc_hd__a22o_1 _2760_ (.A1(net253),
    .A2(net200),
    .B1(net136),
    .B2(net1214),
    .X(_0773_));
 sky130_fd_sc_hd__a22o_1 _2761_ (.A1(net251),
    .A2(net201),
    .B1(net136),
    .B2(net1852),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _2762_ (.A1(net249),
    .A2(net200),
    .B1(net136),
    .B2(net1364),
    .X(_0775_));
 sky130_fd_sc_hd__a22o_1 _2763_ (.A1(net225),
    .A2(net201),
    .B1(net137),
    .B2(net624),
    .X(_0776_));
 sky130_fd_sc_hd__a22o_1 _2764_ (.A1(net363),
    .A2(net200),
    .B1(net136),
    .B2(net1384),
    .X(_0777_));
 sky130_fd_sc_hd__a22o_1 _2765_ (.A1(net361),
    .A2(net201),
    .B1(net137),
    .B2(net1270),
    .X(_0778_));
 sky130_fd_sc_hd__a22o_1 _2766_ (.A1(net359),
    .A2(net200),
    .B1(net137),
    .B2(net2330),
    .X(_0779_));
 sky130_fd_sc_hd__a22o_1 _2767_ (.A1(net357),
    .A2(net201),
    .B1(net137),
    .B2(net2014),
    .X(_0780_));
 sky130_fd_sc_hd__a22o_1 _2768_ (.A1(net355),
    .A2(net201),
    .B1(net137),
    .B2(net892),
    .X(_0781_));
 sky130_fd_sc_hd__a22o_1 _2769_ (.A1(net353),
    .A2(net201),
    .B1(net137),
    .B2(net714),
    .X(_0782_));
 sky130_fd_sc_hd__a22o_1 _2770_ (.A1(net351),
    .A2(net200),
    .B1(net137),
    .B2(net1724),
    .X(_0783_));
 sky130_fd_sc_hd__a22o_1 _2771_ (.A1(net349),
    .A2(net200),
    .B1(net136),
    .B2(net1992),
    .X(_0784_));
 sky130_fd_sc_hd__a22o_1 _2772_ (.A1(net347),
    .A2(net201),
    .B1(net137),
    .B2(net1024),
    .X(_0785_));
 sky130_fd_sc_hd__a22o_1 _2773_ (.A1(net316),
    .A2(net201),
    .B1(net137),
    .B2(net1408),
    .X(_0786_));
 sky130_fd_sc_hd__a22o_1 _2774_ (.A1(net314),
    .A2(net200),
    .B1(net136),
    .B2(net1544),
    .X(_0787_));
 sky130_fd_sc_hd__a22o_1 _2775_ (.A1(net312),
    .A2(net200),
    .B1(net136),
    .B2(net1578),
    .X(_0788_));
 sky130_fd_sc_hd__a22o_1 _2776_ (.A1(net310),
    .A2(net200),
    .B1(net136),
    .B2(net1148),
    .X(_0789_));
 sky130_fd_sc_hd__a22o_1 _2777_ (.A1(net308),
    .A2(net200),
    .B1(net136),
    .B2(net2088),
    .X(_0790_));
 sky130_fd_sc_hd__a22o_1 _2778_ (.A1(net306),
    .A2(net200),
    .B1(net136),
    .B2(net1648),
    .X(_0791_));
 sky130_fd_sc_hd__a22o_1 _2779_ (.A1(net304),
    .A2(net200),
    .B1(net136),
    .B2(net2232),
    .X(_0792_));
 sky130_fd_sc_hd__a22o_1 _2780_ (.A1(net301),
    .A2(net201),
    .B1(net137),
    .B2(net632),
    .X(_0793_));
 sky130_fd_sc_hd__a22o_1 _2781_ (.A1(net299),
    .A2(net201),
    .B1(net136),
    .B2(net1212),
    .X(_0794_));
 sky130_fd_sc_hd__a22o_1 _2782_ (.A1(net297),
    .A2(net200),
    .B1(net136),
    .B2(net666),
    .X(_0795_));
 sky130_fd_sc_hd__a22o_1 _2783_ (.A1(net266),
    .A2(net200),
    .B1(net136),
    .B2(net662),
    .X(_0796_));
 sky130_fd_sc_hd__a22o_1 _2784_ (.A1(net265),
    .A2(net201),
    .B1(net137),
    .B2(net2152),
    .X(_0797_));
 sky130_fd_sc_hd__nor3_4 _2785_ (.A(net232),
    .B(net239),
    .C(net247),
    .Y(_1711_));
 sky130_fd_sc_hd__and4_1 _2786_ (.A(net294),
    .B(net342),
    .C(net216),
    .D(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__nand2_1 _2787_ (.A(_1687_),
    .B(_1711_),
    .Y(_1713_));
 sky130_fd_sc_hd__nor2_1 _2788_ (.A(net369),
    .B(net199),
    .Y(_1714_));
 sky130_fd_sc_hd__or2_2 _2789_ (.A(net366),
    .B(net199),
    .X(_1715_));
 sky130_fd_sc_hd__o22a_1 _2790_ (.A1(net227),
    .A2(_1713_),
    .B1(_1715_),
    .B2(net410),
    .X(_0798_));
 sky130_fd_sc_hd__o22a_1 _2791_ (.A1(net346),
    .A2(_1713_),
    .B1(_1715_),
    .B2(net372),
    .X(_0799_));
 sky130_fd_sc_hd__a22o_1 _2792_ (.A1(net269),
    .A2(net198),
    .B1(net134),
    .B2(net1840),
    .X(_0800_));
 sky130_fd_sc_hd__a22o_1 _2793_ (.A1(net261),
    .A2(net199),
    .B1(net135),
    .B2(net692),
    .X(_0801_));
 sky130_fd_sc_hd__o22a_1 _2794_ (.A1(net259),
    .A2(_1713_),
    .B1(_1715_),
    .B2(net460),
    .X(_0802_));
 sky130_fd_sc_hd__o22a_1 _2795_ (.A1(net258),
    .A2(_1713_),
    .B1(_1715_),
    .B2(net458),
    .X(_0803_));
 sky130_fd_sc_hd__a22o_1 _2796_ (.A1(net256),
    .A2(net199),
    .B1(net135),
    .B2(net1658),
    .X(_0804_));
 sky130_fd_sc_hd__a22o_1 _2797_ (.A1(net254),
    .A2(net198),
    .B1(net134),
    .B2(net1694),
    .X(_0805_));
 sky130_fd_sc_hd__a22o_1 _2798_ (.A1(net252),
    .A2(net198),
    .B1(net134),
    .B2(net1644),
    .X(_0806_));
 sky130_fd_sc_hd__a22o_1 _2799_ (.A1(net250),
    .A2(net198),
    .B1(net134),
    .B2(net758),
    .X(_0807_));
 sky130_fd_sc_hd__a22o_1 _2800_ (.A1(net226),
    .A2(net199),
    .B1(net135),
    .B2(net860),
    .X(_0808_));
 sky130_fd_sc_hd__a22o_1 _2801_ (.A1(net364),
    .A2(net198),
    .B1(net134),
    .B2(net868),
    .X(_0809_));
 sky130_fd_sc_hd__a22o_1 _2802_ (.A1(net362),
    .A2(net199),
    .B1(net135),
    .B2(net1100),
    .X(_0810_));
 sky130_fd_sc_hd__a22o_1 _2803_ (.A1(net360),
    .A2(net199),
    .B1(net134),
    .B2(net1486),
    .X(_0811_));
 sky130_fd_sc_hd__a22o_1 _2804_ (.A1(net358),
    .A2(net199),
    .B1(net135),
    .B2(net2112),
    .X(_0812_));
 sky130_fd_sc_hd__a22o_1 _2805_ (.A1(net356),
    .A2(net198),
    .B1(net135),
    .B2(net1012),
    .X(_0813_));
 sky130_fd_sc_hd__a22o_1 _2806_ (.A1(net354),
    .A2(net199),
    .B1(net135),
    .B2(net722),
    .X(_0814_));
 sky130_fd_sc_hd__a22o_1 _2807_ (.A1(net352),
    .A2(net199),
    .B1(net135),
    .B2(net1752),
    .X(_0815_));
 sky130_fd_sc_hd__a22o_1 _2808_ (.A1(net350),
    .A2(net198),
    .B1(net134),
    .B2(net1468),
    .X(_0816_));
 sky130_fd_sc_hd__a22o_1 _2809_ (.A1(net348),
    .A2(net199),
    .B1(net135),
    .B2(net1662),
    .X(_0817_));
 sky130_fd_sc_hd__a22o_1 _2810_ (.A1(net317),
    .A2(net199),
    .B1(net135),
    .B2(net1996),
    .X(_0818_));
 sky130_fd_sc_hd__a22o_1 _2811_ (.A1(net315),
    .A2(net198),
    .B1(net134),
    .B2(net770),
    .X(_0819_));
 sky130_fd_sc_hd__a22o_1 _2812_ (.A1(net313),
    .A2(net198),
    .B1(net134),
    .B2(net2120),
    .X(_0820_));
 sky130_fd_sc_hd__a22o_1 _2813_ (.A1(net311),
    .A2(net198),
    .B1(net134),
    .B2(net1952),
    .X(_0821_));
 sky130_fd_sc_hd__a22o_1 _2814_ (.A1(net309),
    .A2(net198),
    .B1(net134),
    .B2(net2084),
    .X(_0822_));
 sky130_fd_sc_hd__a22o_1 _2815_ (.A1(net307),
    .A2(net198),
    .B1(net134),
    .B2(net1390),
    .X(_0823_));
 sky130_fd_sc_hd__a22o_1 _2816_ (.A1(net303),
    .A2(net198),
    .B1(net134),
    .B2(net1110),
    .X(_0824_));
 sky130_fd_sc_hd__a22o_1 _2817_ (.A1(net302),
    .A2(net199),
    .B1(net135),
    .B2(net1898),
    .X(_0825_));
 sky130_fd_sc_hd__a22o_1 _2818_ (.A1(net300),
    .A2(net198),
    .B1(net134),
    .B2(net1910),
    .X(_0826_));
 sky130_fd_sc_hd__a22o_1 _2819_ (.A1(net298),
    .A2(net198),
    .B1(net134),
    .B2(net1168),
    .X(_0827_));
 sky130_fd_sc_hd__a22o_1 _2820_ (.A1(net267),
    .A2(net198),
    .B1(net134),
    .B2(net1614),
    .X(_0828_));
 sky130_fd_sc_hd__a22o_1 _2821_ (.A1(net264),
    .A2(net199),
    .B1(net135),
    .B2(net2162),
    .X(_0829_));
 sky130_fd_sc_hd__and3_2 _2822_ (.A(net217),
    .B(_1681_),
    .C(_1693_),
    .X(_1716_));
 sky130_fd_sc_hd__nand2_1 _2823_ (.A(_1681_),
    .B(_1694_),
    .Y(_1717_));
 sky130_fd_sc_hd__nor2_1 _2824_ (.A(net367),
    .B(net197),
    .Y(_1718_));
 sky130_fd_sc_hd__or2_1 _2825_ (.A(net365),
    .B(net197),
    .X(_1719_));
 sky130_fd_sc_hd__o22a_1 _2826_ (.A1(net228),
    .A2(_1717_),
    .B1(_1719_),
    .B2(net558),
    .X(_0830_));
 sky130_fd_sc_hd__o22a_1 _2827_ (.A1(net345),
    .A2(_1717_),
    .B1(_1719_),
    .B2(net464),
    .X(_0831_));
 sky130_fd_sc_hd__a22o_1 _2828_ (.A1(net268),
    .A2(net196),
    .B1(net132),
    .B2(net690),
    .X(_0832_));
 sky130_fd_sc_hd__a22o_1 _2829_ (.A1(net261),
    .A2(net196),
    .B1(net132),
    .B2(net2406),
    .X(_0833_));
 sky130_fd_sc_hd__o22a_1 _2830_ (.A1(net260),
    .A2(_1717_),
    .B1(_1719_),
    .B2(net564),
    .X(_0834_));
 sky130_fd_sc_hd__o22a_1 _2831_ (.A1(net257),
    .A2(_1717_),
    .B1(_1719_),
    .B2(net560),
    .X(_0835_));
 sky130_fd_sc_hd__a22o_1 _2832_ (.A1(net255),
    .A2(net197),
    .B1(net133),
    .B2(net1382),
    .X(_0836_));
 sky130_fd_sc_hd__a22o_1 _2833_ (.A1(net253),
    .A2(net196),
    .B1(net132),
    .B2(net2098),
    .X(_0837_));
 sky130_fd_sc_hd__a22o_1 _2834_ (.A1(net251),
    .A2(net197),
    .B1(net133),
    .B2(net2356),
    .X(_0838_));
 sky130_fd_sc_hd__a22o_1 _2835_ (.A1(net249),
    .A2(net196),
    .B1(net132),
    .B2(net2114),
    .X(_0839_));
 sky130_fd_sc_hd__a22o_1 _2836_ (.A1(net225),
    .A2(net197),
    .B1(net133),
    .B2(net1526),
    .X(_0840_));
 sky130_fd_sc_hd__a22o_1 _2837_ (.A1(net363),
    .A2(net196),
    .B1(net132),
    .B2(net1600),
    .X(_0841_));
 sky130_fd_sc_hd__a22o_1 _2838_ (.A1(net361),
    .A2(net197),
    .B1(net133),
    .B2(net1370),
    .X(_0842_));
 sky130_fd_sc_hd__a22o_1 _2839_ (.A1(net359),
    .A2(net196),
    .B1(net132),
    .B2(net2012),
    .X(_0843_));
 sky130_fd_sc_hd__a22o_1 _2840_ (.A1(net357),
    .A2(net197),
    .B1(net133),
    .B2(net1984),
    .X(_0844_));
 sky130_fd_sc_hd__a22o_1 _2841_ (.A1(net355),
    .A2(net197),
    .B1(net133),
    .B2(net2298),
    .X(_0845_));
 sky130_fd_sc_hd__a22o_1 _2842_ (.A1(net353),
    .A2(net197),
    .B1(net133),
    .B2(net1850),
    .X(_0846_));
 sky130_fd_sc_hd__a22o_1 _2843_ (.A1(net351),
    .A2(net197),
    .B1(net133),
    .B2(net1138),
    .X(_0847_));
 sky130_fd_sc_hd__a22o_1 _2844_ (.A1(net349),
    .A2(net196),
    .B1(net132),
    .B2(net2264),
    .X(_0848_));
 sky130_fd_sc_hd__a22o_1 _2845_ (.A1(net347),
    .A2(net197),
    .B1(net133),
    .B2(net1464),
    .X(_0849_));
 sky130_fd_sc_hd__a22o_1 _2846_ (.A1(net316),
    .A2(net197),
    .B1(net133),
    .B2(net2034),
    .X(_0850_));
 sky130_fd_sc_hd__a22o_1 _2847_ (.A1(net314),
    .A2(net196),
    .B1(net132),
    .B2(net2270),
    .X(_0851_));
 sky130_fd_sc_hd__a22o_1 _2848_ (.A1(net312),
    .A2(net196),
    .B1(net132),
    .B2(net2068),
    .X(_0852_));
 sky130_fd_sc_hd__a22o_1 _2849_ (.A1(net310),
    .A2(net196),
    .B1(net132),
    .B2(net1512),
    .X(_0853_));
 sky130_fd_sc_hd__a22o_1 _2850_ (.A1(net308),
    .A2(net196),
    .B1(net132),
    .B2(net1536),
    .X(_0854_));
 sky130_fd_sc_hd__a22o_1 _2851_ (.A1(net306),
    .A2(net196),
    .B1(net132),
    .B2(net2040),
    .X(_0855_));
 sky130_fd_sc_hd__a22o_1 _2852_ (.A1(net303),
    .A2(net196),
    .B1(net132),
    .B2(net1940),
    .X(_0856_));
 sky130_fd_sc_hd__a22o_1 _2853_ (.A1(net301),
    .A2(net197),
    .B1(net133),
    .B2(net1884),
    .X(_0857_));
 sky130_fd_sc_hd__a22o_1 _2854_ (.A1(net299),
    .A2(net196),
    .B1(net132),
    .B2(net792),
    .X(_0858_));
 sky130_fd_sc_hd__a22o_1 _2855_ (.A1(net297),
    .A2(net196),
    .B1(net132),
    .B2(net2212),
    .X(_0859_));
 sky130_fd_sc_hd__a22o_1 _2856_ (.A1(net266),
    .A2(net196),
    .B1(net132),
    .B2(net1556),
    .X(_0860_));
 sky130_fd_sc_hd__a22o_1 _2857_ (.A1(net264),
    .A2(net197),
    .B1(net133),
    .B2(net1262),
    .X(_0861_));
 sky130_fd_sc_hd__and3_1 _2858_ (.A(net216),
    .B(_1675_),
    .C(_1711_),
    .X(_1720_));
 sky130_fd_sc_hd__nand2_2 _2859_ (.A(_1676_),
    .B(_1711_),
    .Y(_1721_));
 sky130_fd_sc_hd__nor2_1 _2860_ (.A(net369),
    .B(net195),
    .Y(_1722_));
 sky130_fd_sc_hd__or2_2 _2861_ (.A(net366),
    .B(net195),
    .X(_1723_));
 sky130_fd_sc_hd__o22a_1 _2862_ (.A1(net227),
    .A2(_1721_),
    .B1(_1723_),
    .B2(net510),
    .X(_0862_));
 sky130_fd_sc_hd__o22a_1 _2863_ (.A1(net346),
    .A2(_1721_),
    .B1(_1723_),
    .B2(net390),
    .X(_0863_));
 sky130_fd_sc_hd__a22o_1 _2864_ (.A1(net269),
    .A2(net194),
    .B1(net130),
    .B2(net634),
    .X(_0864_));
 sky130_fd_sc_hd__a22o_1 _2865_ (.A1(net261),
    .A2(net195),
    .B1(net131),
    .B2(net986),
    .X(_0865_));
 sky130_fd_sc_hd__o22a_1 _2866_ (.A1(net259),
    .A2(_1721_),
    .B1(_1723_),
    .B2(net590),
    .X(_0866_));
 sky130_fd_sc_hd__o22a_1 _2867_ (.A1(net258),
    .A2(_1721_),
    .B1(_1723_),
    .B2(net550),
    .X(_0867_));
 sky130_fd_sc_hd__a22o_1 _2868_ (.A1(net256),
    .A2(net195),
    .B1(net131),
    .B2(net1530),
    .X(_0868_));
 sky130_fd_sc_hd__a22o_1 _2869_ (.A1(net254),
    .A2(net194),
    .B1(net130),
    .B2(net1904),
    .X(_0869_));
 sky130_fd_sc_hd__a22o_1 _2870_ (.A1(net252),
    .A2(net194),
    .B1(net130),
    .B2(net728),
    .X(_0870_));
 sky130_fd_sc_hd__a22o_1 _2871_ (.A1(net250),
    .A2(net194),
    .B1(net130),
    .B2(net612),
    .X(_0871_));
 sky130_fd_sc_hd__a22o_1 _2872_ (.A1(net226),
    .A2(net195),
    .B1(net131),
    .B2(net1744),
    .X(_0872_));
 sky130_fd_sc_hd__a22o_1 _2873_ (.A1(net364),
    .A2(net194),
    .B1(net130),
    .B2(net1354),
    .X(_0873_));
 sky130_fd_sc_hd__a22o_1 _2874_ (.A1(net362),
    .A2(net195),
    .B1(net131),
    .B2(net654),
    .X(_0874_));
 sky130_fd_sc_hd__a22o_1 _2875_ (.A1(net360),
    .A2(net195),
    .B1(net130),
    .B2(net1114),
    .X(_0875_));
 sky130_fd_sc_hd__a22o_1 _2876_ (.A1(net358),
    .A2(net195),
    .B1(net131),
    .B2(net1832),
    .X(_0876_));
 sky130_fd_sc_hd__a22o_1 _2877_ (.A1(net356),
    .A2(net194),
    .B1(net131),
    .B2(net1240),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _2878_ (.A1(net354),
    .A2(net195),
    .B1(net131),
    .B2(net820),
    .X(_0878_));
 sky130_fd_sc_hd__a22o_1 _2879_ (.A1(net352),
    .A2(net195),
    .B1(net131),
    .B2(net1476),
    .X(_0879_));
 sky130_fd_sc_hd__a22o_1 _2880_ (.A1(net350),
    .A2(net194),
    .B1(net130),
    .B2(net1624),
    .X(_0880_));
 sky130_fd_sc_hd__a22o_1 _2881_ (.A1(net348),
    .A2(net195),
    .B1(net131),
    .B2(net2256),
    .X(_0881_));
 sky130_fd_sc_hd__a22o_1 _2882_ (.A1(net317),
    .A2(net195),
    .B1(net131),
    .B2(net1490),
    .X(_0882_));
 sky130_fd_sc_hd__a22o_1 _2883_ (.A1(net315),
    .A2(net194),
    .B1(net130),
    .B2(net802),
    .X(_0883_));
 sky130_fd_sc_hd__a22o_1 _2884_ (.A1(net313),
    .A2(net194),
    .B1(net130),
    .B2(net1894),
    .X(_0884_));
 sky130_fd_sc_hd__a22o_1 _2885_ (.A1(net311),
    .A2(net194),
    .B1(net130),
    .B2(net1442),
    .X(_0885_));
 sky130_fd_sc_hd__a22o_1 _2886_ (.A1(net309),
    .A2(net194),
    .B1(net130),
    .B2(net1336),
    .X(_0886_));
 sky130_fd_sc_hd__a22o_1 _2887_ (.A1(net307),
    .A2(net194),
    .B1(net130),
    .B2(net1902),
    .X(_0887_));
 sky130_fd_sc_hd__a22o_1 _2888_ (.A1(net303),
    .A2(net194),
    .B1(net130),
    .B2(net2070),
    .X(_0888_));
 sky130_fd_sc_hd__a22o_1 _2889_ (.A1(net302),
    .A2(net195),
    .B1(net131),
    .B2(net1500),
    .X(_0889_));
 sky130_fd_sc_hd__a22o_1 _2890_ (.A1(net300),
    .A2(net194),
    .B1(net130),
    .B2(net958),
    .X(_0890_));
 sky130_fd_sc_hd__a22o_1 _2891_ (.A1(net298),
    .A2(net194),
    .B1(net130),
    .B2(net1016),
    .X(_0891_));
 sky130_fd_sc_hd__a22o_1 _2892_ (.A1(net267),
    .A2(net194),
    .B1(net130),
    .B2(net1726),
    .X(_0892_));
 sky130_fd_sc_hd__a22o_1 _2893_ (.A1(net264),
    .A2(net195),
    .B1(net131),
    .B2(net1720),
    .X(_0893_));
 sky130_fd_sc_hd__and4_2 _2894_ (.A(net283),
    .B(net331),
    .C(_1027_),
    .D(net217),
    .X(_1724_));
 sky130_fd_sc_hd__nand2_2 _2895_ (.A(_1027_),
    .B(_1687_),
    .Y(_1725_));
 sky130_fd_sc_hd__nor2_1 _2896_ (.A(net367),
    .B(net193),
    .Y(_1726_));
 sky130_fd_sc_hd__or2_2 _2897_ (.A(net365),
    .B(net193),
    .X(_1727_));
 sky130_fd_sc_hd__o22a_1 _2898_ (.A1(net228),
    .A2(_1725_),
    .B1(_1727_),
    .B2(net482),
    .X(_0894_));
 sky130_fd_sc_hd__o22a_1 _2899_ (.A1(net345),
    .A2(_1725_),
    .B1(_1727_),
    .B2(net502),
    .X(_0895_));
 sky130_fd_sc_hd__a22o_1 _2900_ (.A1(net268),
    .A2(net192),
    .B1(net128),
    .B2(net2412),
    .X(_0896_));
 sky130_fd_sc_hd__a22o_1 _2901_ (.A1(net263),
    .A2(net193),
    .B1(net129),
    .B2(net2302),
    .X(_0897_));
 sky130_fd_sc_hd__o22a_1 _2902_ (.A1(net260),
    .A2(_1725_),
    .B1(_1727_),
    .B2(net572),
    .X(_0898_));
 sky130_fd_sc_hd__o22a_1 _2903_ (.A1(net257),
    .A2(_1725_),
    .B1(_1727_),
    .B2(net454),
    .X(_0899_));
 sky130_fd_sc_hd__a22o_1 _2904_ (.A1(net255),
    .A2(net193),
    .B1(net129),
    .B2(net1570),
    .X(_0900_));
 sky130_fd_sc_hd__a22o_1 _2905_ (.A1(net253),
    .A2(net192),
    .B1(net128),
    .B2(net2294),
    .X(_0901_));
 sky130_fd_sc_hd__a22o_1 _2906_ (.A1(net251),
    .A2(net193),
    .B1(net129),
    .B2(net1882),
    .X(_0902_));
 sky130_fd_sc_hd__a22o_1 _2907_ (.A1(net249),
    .A2(net192),
    .B1(net128),
    .B2(net2378),
    .X(_0903_));
 sky130_fd_sc_hd__a22o_1 _2908_ (.A1(net225),
    .A2(net193),
    .B1(net129),
    .B2(net1616),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _2909_ (.A1(net363),
    .A2(net192),
    .B1(net128),
    .B2(net2392),
    .X(_0905_));
 sky130_fd_sc_hd__a22o_1 _2910_ (.A1(net361),
    .A2(net193),
    .B1(net129),
    .B2(net1070),
    .X(_0906_));
 sky130_fd_sc_hd__a22o_1 _2911_ (.A1(net359),
    .A2(net192),
    .B1(net128),
    .B2(net2376),
    .X(_0907_));
 sky130_fd_sc_hd__a22o_1 _2912_ (.A1(net357),
    .A2(net193),
    .B1(net129),
    .B2(net2234),
    .X(_0908_));
 sky130_fd_sc_hd__a22o_1 _2913_ (.A1(net355),
    .A2(net192),
    .B1(net128),
    .B2(net2368),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _2914_ (.A1(net353),
    .A2(net193),
    .B1(net129),
    .B2(net1962),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _2915_ (.A1(net351),
    .A2(net193),
    .B1(net129),
    .B2(net1612),
    .X(_0911_));
 sky130_fd_sc_hd__a22o_1 _2916_ (.A1(net349),
    .A2(net192),
    .B1(net128),
    .B2(net2216),
    .X(_0912_));
 sky130_fd_sc_hd__a22o_1 _2917_ (.A1(net347),
    .A2(net193),
    .B1(net129),
    .B2(net2306),
    .X(_0913_));
 sky130_fd_sc_hd__a22o_1 _2918_ (.A1(net316),
    .A2(net193),
    .B1(net129),
    .B2(net2402),
    .X(_0914_));
 sky130_fd_sc_hd__a22o_1 _2919_ (.A1(net314),
    .A2(net192),
    .B1(net128),
    .B2(net1812),
    .X(_0915_));
 sky130_fd_sc_hd__a22o_1 _2920_ (.A1(net312),
    .A2(net192),
    .B1(net128),
    .B2(net2122),
    .X(_0916_));
 sky130_fd_sc_hd__a22o_1 _2921_ (.A1(net310),
    .A2(net192),
    .B1(net128),
    .B2(net2200),
    .X(_0917_));
 sky130_fd_sc_hd__a22o_1 _2922_ (.A1(net308),
    .A2(net192),
    .B1(net128),
    .B2(net972),
    .X(_0918_));
 sky130_fd_sc_hd__a22o_1 _2923_ (.A1(net306),
    .A2(net192),
    .B1(net128),
    .B2(net2382),
    .X(_0919_));
 sky130_fd_sc_hd__a22o_1 _2924_ (.A1(net305),
    .A2(net192),
    .B1(net128),
    .B2(net1050),
    .X(_0920_));
 sky130_fd_sc_hd__a22o_1 _2925_ (.A1(net301),
    .A2(net193),
    .B1(net129),
    .B2(net866),
    .X(_0921_));
 sky130_fd_sc_hd__a22o_1 _2926_ (.A1(net299),
    .A2(net192),
    .B1(net128),
    .B2(net1534),
    .X(_0922_));
 sky130_fd_sc_hd__a22o_1 _2927_ (.A1(net297),
    .A2(net192),
    .B1(net128),
    .B2(net1736),
    .X(_0923_));
 sky130_fd_sc_hd__a22o_1 _2928_ (.A1(net266),
    .A2(net192),
    .B1(net128),
    .B2(net1716),
    .X(_0924_));
 sky130_fd_sc_hd__a22o_1 _2929_ (.A1(net265),
    .A2(net193),
    .B1(net129),
    .B2(net2338),
    .X(_0925_));
 sky130_fd_sc_hd__and4b_1 _2930_ (.A_N(net283),
    .B(net331),
    .C(_1027_),
    .D(net217),
    .X(_1728_));
 sky130_fd_sc_hd__nand2_2 _2931_ (.A(_1027_),
    .B(_1670_),
    .Y(_1729_));
 sky130_fd_sc_hd__nor2_1 _2932_ (.A(net367),
    .B(net190),
    .Y(_1730_));
 sky130_fd_sc_hd__or2_2 _2933_ (.A(net365),
    .B(net191),
    .X(_1731_));
 sky130_fd_sc_hd__o22a_1 _2934_ (.A1(net228),
    .A2(_1729_),
    .B1(_1731_),
    .B2(net1076),
    .X(_0926_));
 sky130_fd_sc_hd__o22a_1 _2935_ (.A1(net345),
    .A2(_1729_),
    .B1(_1731_),
    .B2(net478),
    .X(_0927_));
 sky130_fd_sc_hd__a22o_1 _2936_ (.A1(net268),
    .A2(net190),
    .B1(net126),
    .B2(net2154),
    .X(_0928_));
 sky130_fd_sc_hd__a22o_1 _2937_ (.A1(net263),
    .A2(net191),
    .B1(net127),
    .B2(net2236),
    .X(_0929_));
 sky130_fd_sc_hd__o22a_1 _2938_ (.A1(net260),
    .A2(_1729_),
    .B1(_1731_),
    .B2(net526),
    .X(_0930_));
 sky130_fd_sc_hd__o22a_1 _2939_ (.A1(net257),
    .A2(_1729_),
    .B1(_1731_),
    .B2(net602),
    .X(_0931_));
 sky130_fd_sc_hd__a22o_1 _2940_ (.A1(net255),
    .A2(net191),
    .B1(net127),
    .B2(net1878),
    .X(_0932_));
 sky130_fd_sc_hd__a22o_1 _2941_ (.A1(net253),
    .A2(net190),
    .B1(net126),
    .B2(net2292),
    .X(_0933_));
 sky130_fd_sc_hd__a22o_1 _2942_ (.A1(net251),
    .A2(net190),
    .B1(net126),
    .B2(net2400),
    .X(_0934_));
 sky130_fd_sc_hd__a22o_1 _2943_ (.A1(net249),
    .A2(net190),
    .B1(net126),
    .B2(net2038),
    .X(_0935_));
 sky130_fd_sc_hd__a22o_1 _2944_ (.A1(net225),
    .A2(net190),
    .B1(net127),
    .B2(net2090),
    .X(_0936_));
 sky130_fd_sc_hd__a22o_1 _2945_ (.A1(net363),
    .A2(net190),
    .B1(net126),
    .B2(net1552),
    .X(_0937_));
 sky130_fd_sc_hd__a22o_1 _2946_ (.A1(net361),
    .A2(net191),
    .B1(net127),
    .B2(net1680),
    .X(_0938_));
 sky130_fd_sc_hd__a22o_1 _2947_ (.A1(net359),
    .A2(net191),
    .B1(net126),
    .B2(net2398),
    .X(_0939_));
 sky130_fd_sc_hd__a22o_1 _2948_ (.A1(net357),
    .A2(net191),
    .B1(net127),
    .B2(net1934),
    .X(_0940_));
 sky130_fd_sc_hd__a22o_1 _2949_ (.A1(net355),
    .A2(net190),
    .B1(net126),
    .B2(net2188),
    .X(_0941_));
 sky130_fd_sc_hd__a22o_1 _2950_ (.A1(net353),
    .A2(net191),
    .B1(net127),
    .B2(net1926),
    .X(_0942_));
 sky130_fd_sc_hd__a22o_1 _2951_ (.A1(net351),
    .A2(net191),
    .B1(net127),
    .B2(net1474),
    .X(_0943_));
 sky130_fd_sc_hd__a22o_1 _2952_ (.A1(net349),
    .A2(net191),
    .B1(net126),
    .B2(net2184),
    .X(_0944_));
 sky130_fd_sc_hd__a22o_1 _2953_ (.A1(net347),
    .A2(net191),
    .B1(net127),
    .B2(net2072),
    .X(_0945_));
 sky130_fd_sc_hd__a22o_1 _2954_ (.A1(net316),
    .A2(net191),
    .B1(net127),
    .B2(net2274),
    .X(_0946_));
 sky130_fd_sc_hd__a22o_1 _2955_ (.A1(net314),
    .A2(net191),
    .B1(net127),
    .B2(net2414),
    .X(_0947_));
 sky130_fd_sc_hd__a22o_1 _2956_ (.A1(net312),
    .A2(net190),
    .B1(net126),
    .B2(net1808),
    .X(_0948_));
 sky130_fd_sc_hd__a22o_1 _2957_ (.A1(net310),
    .A2(net190),
    .B1(net126),
    .B2(net1346),
    .X(_0949_));
 sky130_fd_sc_hd__a22o_1 _2958_ (.A1(net308),
    .A2(net190),
    .B1(net126),
    .B2(net2130),
    .X(_0950_));
 sky130_fd_sc_hd__a22o_1 _2959_ (.A1(net306),
    .A2(net190),
    .B1(net126),
    .B2(net2390),
    .X(_0951_));
 sky130_fd_sc_hd__a22o_1 _2960_ (.A1(net305),
    .A2(net190),
    .B1(net126),
    .B2(net1438),
    .X(_0952_));
 sky130_fd_sc_hd__a22o_1 _2961_ (.A1(net301),
    .A2(net191),
    .B1(net127),
    .B2(net898),
    .X(_0953_));
 sky130_fd_sc_hd__a22o_1 _2962_ (.A1(net299),
    .A2(net190),
    .B1(net126),
    .B2(net1446),
    .X(_0954_));
 sky130_fd_sc_hd__a22o_1 _2963_ (.A1(net297),
    .A2(net190),
    .B1(net126),
    .B2(net1814),
    .X(_0955_));
 sky130_fd_sc_hd__a22o_1 _2964_ (.A1(net266),
    .A2(net190),
    .B1(net126),
    .B2(net1966),
    .X(_0956_));
 sky130_fd_sc_hd__a22o_1 _2965_ (.A1(net265),
    .A2(net191),
    .B1(net127),
    .B2(net2372),
    .X(_0957_));
 sky130_fd_sc_hd__nor3b_4 _2966_ (.A(net232),
    .B(net239),
    .C_N(net247),
    .Y(_1732_));
 sky130_fd_sc_hd__and3_1 _2967_ (.A(net216),
    .B(_1675_),
    .C(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__nand2_1 _2968_ (.A(_1676_),
    .B(_1732_),
    .Y(_1734_));
 sky130_fd_sc_hd__nor2_1 _2969_ (.A(net368),
    .B(net189),
    .Y(_1735_));
 sky130_fd_sc_hd__or2_1 _2970_ (.A(net368),
    .B(net189),
    .X(_1736_));
 sky130_fd_sc_hd__o22a_1 _2971_ (.A1(net227),
    .A2(_1734_),
    .B1(_1736_),
    .B2(net880),
    .X(_0958_));
 sky130_fd_sc_hd__o22a_1 _2972_ (.A1(net346),
    .A2(_1734_),
    .B1(_1736_),
    .B2(net580),
    .X(_0959_));
 sky130_fd_sc_hd__a22o_1 _2973_ (.A1(net269),
    .A2(net188),
    .B1(net124),
    .B2(net970),
    .X(_0960_));
 sky130_fd_sc_hd__a22o_1 _2974_ (.A1(net261),
    .A2(net189),
    .B1(net125),
    .B2(net1406),
    .X(_0961_));
 sky130_fd_sc_hd__o22a_1 _2975_ (.A1(net259),
    .A2(_1734_),
    .B1(_1736_),
    .B2(net516),
    .X(_0962_));
 sky130_fd_sc_hd__o22a_1 _2976_ (.A1(net258),
    .A2(_1734_),
    .B1(_1736_),
    .B2(net604),
    .X(_0963_));
 sky130_fd_sc_hd__a22o_1 _2977_ (.A1(net256),
    .A2(net189),
    .B1(net124),
    .B2(net1960),
    .X(_0964_));
 sky130_fd_sc_hd__a22o_1 _2978_ (.A1(net254),
    .A2(net188),
    .B1(net124),
    .B2(net684),
    .X(_0965_));
 sky130_fd_sc_hd__a22o_1 _2979_ (.A1(net252),
    .A2(net189),
    .B1(net124),
    .B2(net746),
    .X(_0966_));
 sky130_fd_sc_hd__a22o_1 _2980_ (.A1(net250),
    .A2(net188),
    .B1(net124),
    .B2(net1008),
    .X(_0967_));
 sky130_fd_sc_hd__a22o_1 _2981_ (.A1(net226),
    .A2(net189),
    .B1(net125),
    .B2(net1750),
    .X(_0968_));
 sky130_fd_sc_hd__a22o_1 _2982_ (.A1(net364),
    .A2(net188),
    .B1(net124),
    .B2(net1684),
    .X(_0969_));
 sky130_fd_sc_hd__a22o_1 _2983_ (.A1(net362),
    .A2(net189),
    .B1(net125),
    .B2(net616),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _2984_ (.A1(net360),
    .A2(net188),
    .B1(net124),
    .B2(net1290),
    .X(_0971_));
 sky130_fd_sc_hd__a22o_1 _2985_ (.A1(net358),
    .A2(net189),
    .B1(net125),
    .B2(net2282),
    .X(_0972_));
 sky130_fd_sc_hd__a22o_1 _2986_ (.A1(net356),
    .A2(net188),
    .B1(net125),
    .B2(net1422),
    .X(_0973_));
 sky130_fd_sc_hd__a22o_1 _2987_ (.A1(net354),
    .A2(net189),
    .B1(net125),
    .B2(net674),
    .X(_0974_));
 sky130_fd_sc_hd__a22o_1 _2988_ (.A1(net352),
    .A2(net189),
    .B1(net125),
    .B2(net1174),
    .X(_0975_));
 sky130_fd_sc_hd__a22o_1 _2989_ (.A1(net350),
    .A2(net188),
    .B1(net124),
    .B2(net2358),
    .X(_0976_));
 sky130_fd_sc_hd__a22o_1 _2990_ (.A1(net348),
    .A2(net189),
    .B1(net125),
    .B2(net1068),
    .X(_0977_));
 sky130_fd_sc_hd__a22o_1 _2991_ (.A1(net317),
    .A2(net189),
    .B1(net125),
    .B2(net2046),
    .X(_0978_));
 sky130_fd_sc_hd__a22o_1 _2992_ (.A1(net315),
    .A2(net188),
    .B1(net124),
    .B2(net1220),
    .X(_0979_));
 sky130_fd_sc_hd__a22o_1 _2993_ (.A1(net313),
    .A2(net188),
    .B1(net124),
    .B2(net2028),
    .X(_0980_));
 sky130_fd_sc_hd__a22o_1 _2994_ (.A1(net311),
    .A2(net188),
    .B1(net124),
    .B2(net1484),
    .X(_0981_));
 sky130_fd_sc_hd__a22o_1 _2995_ (.A1(net309),
    .A2(net188),
    .B1(net124),
    .B2(net2312),
    .X(_0982_));
 sky130_fd_sc_hd__a22o_1 _2996_ (.A1(net307),
    .A2(net188),
    .B1(net124),
    .B2(net2366),
    .X(_0983_));
 sky130_fd_sc_hd__a22o_1 _2997_ (.A1(net303),
    .A2(net188),
    .B1(net125),
    .B2(net2170),
    .X(_0984_));
 sky130_fd_sc_hd__a22o_1 _2998_ (.A1(net302),
    .A2(net189),
    .B1(net125),
    .B2(net740),
    .X(_0985_));
 sky130_fd_sc_hd__a22o_1 _2999_ (.A1(net300),
    .A2(net188),
    .B1(net124),
    .B2(net738),
    .X(_0986_));
 sky130_fd_sc_hd__a22o_1 _3000_ (.A1(net298),
    .A2(net188),
    .B1(net124),
    .B2(net2144),
    .X(_0987_));
 sky130_fd_sc_hd__a22o_1 _3001_ (.A1(net267),
    .A2(net188),
    .B1(net124),
    .B2(net1622),
    .X(_0988_));
 sky130_fd_sc_hd__a22o_1 _3002_ (.A1(net264),
    .A2(net189),
    .B1(net125),
    .B2(net786),
    .X(_0989_));
 sky130_fd_sc_hd__and4b_2 _3003_ (.A_N(net284),
    .B(net332),
    .C(net217),
    .D(_1681_),
    .X(_1737_));
 sky130_fd_sc_hd__nand2_1 _3004_ (.A(_1670_),
    .B(_1681_),
    .Y(_1738_));
 sky130_fd_sc_hd__nor2_1 _3005_ (.A(net367),
    .B(net186),
    .Y(_1739_));
 sky130_fd_sc_hd__or2_1 _3006_ (.A(net365),
    .B(net187),
    .X(_1740_));
 sky130_fd_sc_hd__o22a_1 _3007_ (.A1(net228),
    .A2(_1738_),
    .B1(_1740_),
    .B2(net508),
    .X(_0990_));
 sky130_fd_sc_hd__o22a_1 _3008_ (.A1(net345),
    .A2(_1738_),
    .B1(_1740_),
    .B2(net466),
    .X(_0991_));
 sky130_fd_sc_hd__a22o_1 _3009_ (.A1(net268),
    .A2(net186),
    .B1(net122),
    .B2(net1880),
    .X(_0992_));
 sky130_fd_sc_hd__a22o_1 _3010_ (.A1(net261),
    .A2(net187),
    .B1(net122),
    .B2(net2226),
    .X(_0993_));
 sky130_fd_sc_hd__o22a_1 _3011_ (.A1(net260),
    .A2(_1738_),
    .B1(_1740_),
    .B2(net582),
    .X(_0994_));
 sky130_fd_sc_hd__o22a_1 _3012_ (.A1(net257),
    .A2(_1738_),
    .B1(_1740_),
    .B2(net726),
    .X(_0995_));
 sky130_fd_sc_hd__a22o_1 _3013_ (.A1(net255),
    .A2(net187),
    .B1(net123),
    .B2(net2314),
    .X(_0996_));
 sky130_fd_sc_hd__a22o_1 _3014_ (.A1(net253),
    .A2(net186),
    .B1(net122),
    .B2(net1958),
    .X(_0997_));
 sky130_fd_sc_hd__a22o_1 _3015_ (.A1(net251),
    .A2(net187),
    .B1(net123),
    .B2(net2416),
    .X(_0998_));
 sky130_fd_sc_hd__a22o_1 _3016_ (.A1(net249),
    .A2(net186),
    .B1(net122),
    .B2(net2142),
    .X(_0999_));
 sky130_fd_sc_hd__a22o_1 _3017_ (.A1(net225),
    .A2(net187),
    .B1(net123),
    .B2(net1672),
    .X(_1000_));
 sky130_fd_sc_hd__a22o_1 _3018_ (.A1(net363),
    .A2(net186),
    .B1(net122),
    .B2(net1610),
    .X(_1001_));
 sky130_fd_sc_hd__a22o_1 _3019_ (.A1(net361),
    .A2(net187),
    .B1(net123),
    .B2(net1386),
    .X(_1002_));
 sky130_fd_sc_hd__a22o_1 _3020_ (.A1(net359),
    .A2(net186),
    .B1(net122),
    .B2(net2348),
    .X(_1003_));
 sky130_fd_sc_hd__a22o_1 _3021_ (.A1(net357),
    .A2(net187),
    .B1(net123),
    .B2(net2360),
    .X(_1004_));
 sky130_fd_sc_hd__a22o_1 _3022_ (.A1(net355),
    .A2(net187),
    .B1(net123),
    .B2(net2332),
    .X(_1005_));
 sky130_fd_sc_hd__a22o_1 _3023_ (.A1(net353),
    .A2(net187),
    .B1(net123),
    .B2(net1862),
    .X(_1006_));
 sky130_fd_sc_hd__a22o_1 _3024_ (.A1(net351),
    .A2(net187),
    .B1(net123),
    .B2(net1982),
    .X(_1007_));
 sky130_fd_sc_hd__a22o_1 _3025_ (.A1(net349),
    .A2(net186),
    .B1(net122),
    .B2(net2158),
    .X(_1008_));
 sky130_fd_sc_hd__a22o_1 _3026_ (.A1(net347),
    .A2(net187),
    .B1(net123),
    .B2(net2076),
    .X(_1009_));
 sky130_fd_sc_hd__a22o_1 _3027_ (.A1(net316),
    .A2(net187),
    .B1(net123),
    .B2(net2238),
    .X(_1010_));
 sky130_fd_sc_hd__a22o_1 _3028_ (.A1(net314),
    .A2(net186),
    .B1(net122),
    .B2(net2300),
    .X(_1011_));
 sky130_fd_sc_hd__a22o_1 _3029_ (.A1(net312),
    .A2(net186),
    .B1(net122),
    .B2(net818),
    .X(_1012_));
 sky130_fd_sc_hd__a22o_1 _3030_ (.A1(net310),
    .A2(net186),
    .B1(net122),
    .B2(net1820),
    .X(_1013_));
 sky130_fd_sc_hd__a22o_1 _3031_ (.A1(net308),
    .A2(net186),
    .B1(net122),
    .B2(net2334),
    .X(_1014_));
 sky130_fd_sc_hd__a22o_1 _3032_ (.A1(net306),
    .A2(net186),
    .B1(net122),
    .B2(net1676),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_1 _3033_ (.A1(net303),
    .A2(net186),
    .B1(net122),
    .B2(net1458),
    .X(_1016_));
 sky130_fd_sc_hd__a22o_1 _3034_ (.A1(net301),
    .A2(net187),
    .B1(net123),
    .B2(net1788),
    .X(_1017_));
 sky130_fd_sc_hd__a22o_1 _3035_ (.A1(net299),
    .A2(net186),
    .B1(net122),
    .B2(net2214),
    .X(_1018_));
 sky130_fd_sc_hd__a22o_1 _3036_ (.A1(net297),
    .A2(net186),
    .B1(net122),
    .B2(net1932),
    .X(_1019_));
 sky130_fd_sc_hd__a22o_1 _3037_ (.A1(net266),
    .A2(net186),
    .B1(net122),
    .B2(net1478),
    .X(_1020_));
 sky130_fd_sc_hd__a22o_1 _3038_ (.A1(net264),
    .A2(net187),
    .B1(net123),
    .B2(net2364),
    .X(_1021_));
 sky130_fd_sc_hd__nor3b_4 _3039_ (.A(net232),
    .B(net247),
    .C_N(net239),
    .Y(_1741_));
 sky130_fd_sc_hd__and3_1 _3040_ (.A(net216),
    .B(_1693_),
    .C(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__nand2_2 _3041_ (.A(_1694_),
    .B(_1741_),
    .Y(_1743_));
 sky130_fd_sc_hd__nor2_1 _3042_ (.A(net368),
    .B(net185),
    .Y(_1744_));
 sky130_fd_sc_hd__or2_2 _3043_ (.A(net366),
    .B(net185),
    .X(_1745_));
 sky130_fd_sc_hd__o22a_1 _3044_ (.A1(net227),
    .A2(_1743_),
    .B1(_1745_),
    .B2(net522),
    .X(_1022_));
 sky130_fd_sc_hd__o22a_1 _3045_ (.A1(net346),
    .A2(_1743_),
    .B1(_1745_),
    .B2(net486),
    .X(_1023_));
 sky130_fd_sc_hd__a22o_1 _3046_ (.A1(net269),
    .A2(net184),
    .B1(net120),
    .B2(net1356),
    .X(_1024_));
 sky130_fd_sc_hd__a22o_1 _3047_ (.A1(net261),
    .A2(net185),
    .B1(net121),
    .B2(net682),
    .X(_0000_));
 sky130_fd_sc_hd__o22a_1 _3048_ (.A1(net259),
    .A2(_1743_),
    .B1(_1745_),
    .B2(net500),
    .X(_0001_));
 sky130_fd_sc_hd__o22a_1 _3049_ (.A1(net258),
    .A2(_1743_),
    .B1(_1745_),
    .B2(net384),
    .X(_0002_));
 sky130_fd_sc_hd__a22o_1 _3050_ (.A1(net256),
    .A2(net185),
    .B1(net121),
    .B2(net1990),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _3051_ (.A1(net254),
    .A2(net184),
    .B1(net120),
    .B2(net2310),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _3052_ (.A1(net252),
    .A2(net184),
    .B1(net120),
    .B2(net2182),
    .X(_0005_));
 sky130_fd_sc_hd__a22o_1 _3053_ (.A1(net250),
    .A2(net184),
    .B1(net120),
    .B2(net782),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _3054_ (.A1(net226),
    .A2(net185),
    .B1(net121),
    .B2(net1834),
    .X(_0007_));
 sky130_fd_sc_hd__a22o_1 _3055_ (.A1(net364),
    .A2(net184),
    .B1(net120),
    .B2(net2374),
    .X(_0008_));
 sky130_fd_sc_hd__a22o_1 _3056_ (.A1(net362),
    .A2(net185),
    .B1(net121),
    .B2(net1554),
    .X(_0009_));
 sky130_fd_sc_hd__a22o_1 _3057_ (.A1(net360),
    .A2(net184),
    .B1(net120),
    .B2(net2262),
    .X(_0010_));
 sky130_fd_sc_hd__a22o_1 _3058_ (.A1(net358),
    .A2(net185),
    .B1(net121),
    .B2(net1030),
    .X(_0011_));
 sky130_fd_sc_hd__a22o_1 _3059_ (.A1(net356),
    .A2(net184),
    .B1(net120),
    .B2(net1002),
    .X(_0012_));
 sky130_fd_sc_hd__a22o_1 _3060_ (.A1(net354),
    .A2(net185),
    .B1(net121),
    .B2(net2196),
    .X(_0013_));
 sky130_fd_sc_hd__a22o_1 _3061_ (.A1(net352),
    .A2(net185),
    .B1(net121),
    .B2(net950),
    .X(_0014_));
 sky130_fd_sc_hd__a22o_1 _3062_ (.A1(net350),
    .A2(net184),
    .B1(net120),
    .B2(net1876),
    .X(_0015_));
 sky130_fd_sc_hd__a22o_1 _3063_ (.A1(net348),
    .A2(net185),
    .B1(net121),
    .B2(net876),
    .X(_0016_));
 sky130_fd_sc_hd__a22o_1 _3064_ (.A1(net317),
    .A2(net185),
    .B1(net121),
    .B2(net1580),
    .X(_0017_));
 sky130_fd_sc_hd__a22o_1 _3065_ (.A1(net315),
    .A2(net184),
    .B1(net120),
    .B2(net1154),
    .X(_0018_));
 sky130_fd_sc_hd__a22o_1 _3066_ (.A1(net313),
    .A2(net184),
    .B1(net120),
    .B2(net1194),
    .X(_0019_));
 sky130_fd_sc_hd__a22o_1 _3067_ (.A1(net311),
    .A2(net184),
    .B1(net120),
    .B2(net1916),
    .X(_0020_));
 sky130_fd_sc_hd__a22o_1 _3068_ (.A1(net309),
    .A2(net184),
    .B1(net120),
    .B2(net2344),
    .X(_0021_));
 sky130_fd_sc_hd__a22o_1 _3069_ (.A1(net307),
    .A2(net185),
    .B1(net121),
    .B2(net2062),
    .X(_0022_));
 sky130_fd_sc_hd__a22o_1 _3070_ (.A1(net303),
    .A2(net184),
    .B1(net120),
    .B2(net1890),
    .X(_0023_));
 sky130_fd_sc_hd__a22o_1 _3071_ (.A1(net302),
    .A2(net185),
    .B1(net121),
    .B2(net1792),
    .X(_0024_));
 sky130_fd_sc_hd__a22o_1 _3072_ (.A1(net300),
    .A2(net184),
    .B1(net120),
    .B2(net1320),
    .X(_0025_));
 sky130_fd_sc_hd__a22o_1 _3073_ (.A1(net298),
    .A2(net184),
    .B1(net120),
    .B2(net2194),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_1 _3074_ (.A1(net267),
    .A2(net184),
    .B1(net120),
    .B2(net894),
    .X(_0027_));
 sky130_fd_sc_hd__a22o_1 _3075_ (.A1(net264),
    .A2(net185),
    .B1(net121),
    .B2(net1294),
    .X(_0028_));
 sky130_fd_sc_hd__and4_2 _3076_ (.A(net293),
    .B(net341),
    .C(net216),
    .D(_1732_),
    .X(_1746_));
 sky130_fd_sc_hd__nand2_2 _3077_ (.A(_1687_),
    .B(_1732_),
    .Y(_1747_));
 sky130_fd_sc_hd__nor2_2 _3078_ (.A(net368),
    .B(net183),
    .Y(_1748_));
 sky130_fd_sc_hd__or2_2 _3079_ (.A(net368),
    .B(net183),
    .X(_1749_));
 sky130_fd_sc_hd__o22a_1 _3080_ (.A1(net227),
    .A2(_1747_),
    .B1(_1749_),
    .B2(net556),
    .X(_0029_));
 sky130_fd_sc_hd__o22a_1 _3081_ (.A1(net346),
    .A2(_1747_),
    .B1(_1749_),
    .B2(net606),
    .X(_0030_));
 sky130_fd_sc_hd__a22o_1 _3082_ (.A1(net269),
    .A2(net182),
    .B1(net118),
    .B2(net1546),
    .X(_0031_));
 sky130_fd_sc_hd__a22o_1 _3083_ (.A1(net261),
    .A2(net183),
    .B1(net119),
    .B2(net736),
    .X(_0032_));
 sky130_fd_sc_hd__o22a_1 _3084_ (.A1(net259),
    .A2(_1747_),
    .B1(_1749_),
    .B2(net524),
    .X(_0033_));
 sky130_fd_sc_hd__o22a_1 _3085_ (.A1(net258),
    .A2(_1747_),
    .B1(_1749_),
    .B2(net536),
    .X(_0034_));
 sky130_fd_sc_hd__a22o_1 _3086_ (.A1(net256),
    .A2(net183),
    .B1(net119),
    .B2(net1542),
    .X(_0035_));
 sky130_fd_sc_hd__a22o_1 _3087_ (.A1(net254),
    .A2(net182),
    .B1(net118),
    .B2(net664),
    .X(_0036_));
 sky130_fd_sc_hd__a22o_1 _3088_ (.A1(net252),
    .A2(net183),
    .B1(net118),
    .B2(net1026),
    .X(_0037_));
 sky130_fd_sc_hd__a22o_1 _3089_ (.A1(net250),
    .A2(net182),
    .B1(net118),
    .B2(net1738),
    .X(_0038_));
 sky130_fd_sc_hd__a22o_1 _3090_ (.A1(net226),
    .A2(net183),
    .B1(net119),
    .B2(net1058),
    .X(_0039_));
 sky130_fd_sc_hd__a22o_1 _3091_ (.A1(net364),
    .A2(net182),
    .B1(net118),
    .B2(net2290),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _3092_ (.A1(net362),
    .A2(net183),
    .B1(net119),
    .B2(net712),
    .X(_0041_));
 sky130_fd_sc_hd__a22o_1 _3093_ (.A1(net360),
    .A2(net182),
    .B1(net118),
    .B2(net1956),
    .X(_0042_));
 sky130_fd_sc_hd__a22o_1 _3094_ (.A1(net358),
    .A2(net183),
    .B1(net119),
    .B2(net2266),
    .X(_0043_));
 sky130_fd_sc_hd__a22o_1 _3095_ (.A1(net356),
    .A2(net182),
    .B1(net118),
    .B2(net1156),
    .X(_0044_));
 sky130_fd_sc_hd__a22o_1 _3096_ (.A1(net354),
    .A2(net183),
    .B1(net119),
    .B2(net1322),
    .X(_0045_));
 sky130_fd_sc_hd__a22o_1 _3097_ (.A1(net352),
    .A2(net183),
    .B1(net119),
    .B2(net1470),
    .X(_0046_));
 sky130_fd_sc_hd__a22o_1 _3098_ (.A1(net350),
    .A2(net182),
    .B1(net118),
    .B2(net1688),
    .X(_0047_));
 sky130_fd_sc_hd__a22o_1 _3099_ (.A1(net348),
    .A2(net183),
    .B1(net119),
    .B2(net1650),
    .X(_0048_));
 sky130_fd_sc_hd__a22o_1 _3100_ (.A1(net317),
    .A2(net183),
    .B1(net119),
    .B2(net1912),
    .X(_0049_));
 sky130_fd_sc_hd__a22o_1 _3101_ (.A1(net315),
    .A2(net182),
    .B1(net118),
    .B2(net1434),
    .X(_0050_));
 sky130_fd_sc_hd__a22o_1 _3102_ (.A1(net313),
    .A2(net182),
    .B1(net118),
    .B2(net2276),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_1 _3103_ (.A1(net311),
    .A2(net182),
    .B1(net118),
    .B2(net1258),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _3104_ (.A1(net309),
    .A2(net182),
    .B1(net118),
    .B2(net1856),
    .X(_0053_));
 sky130_fd_sc_hd__a22o_1 _3105_ (.A1(net307),
    .A2(net182),
    .B1(net118),
    .B2(net1810),
    .X(_0054_));
 sky130_fd_sc_hd__a22o_1 _3106_ (.A1(net303),
    .A2(net182),
    .B1(net119),
    .B2(net2074),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _3107_ (.A1(net302),
    .A2(net183),
    .B1(net119),
    .B2(net1404),
    .X(_0056_));
 sky130_fd_sc_hd__a22o_1 _3108_ (.A1(net300),
    .A2(net182),
    .B1(net118),
    .B2(net1416),
    .X(_0057_));
 sky130_fd_sc_hd__a22o_1 _3109_ (.A1(net298),
    .A2(net182),
    .B1(net118),
    .B2(net1700),
    .X(_0058_));
 sky130_fd_sc_hd__a22o_1 _3110_ (.A1(net267),
    .A2(net182),
    .B1(net118),
    .B2(net920),
    .X(_0059_));
 sky130_fd_sc_hd__a22o_1 _3111_ (.A1(net264),
    .A2(net183),
    .B1(net119),
    .B2(net660),
    .X(_0060_));
 sky130_fd_sc_hd__and3_1 _3112_ (.A(net217),
    .B(_1675_),
    .C(_1692_),
    .X(_1750_));
 sky130_fd_sc_hd__nand2_2 _3113_ (.A(_1676_),
    .B(_1692_),
    .Y(_1751_));
 sky130_fd_sc_hd__nor2_1 _3114_ (.A(net365),
    .B(net181),
    .Y(_1752_));
 sky130_fd_sc_hd__or2_2 _3115_ (.A(net365),
    .B(net180),
    .X(_1753_));
 sky130_fd_sc_hd__o22a_1 _3116_ (.A1(net228),
    .A2(_1751_),
    .B1(_1753_),
    .B2(net1762),
    .X(_0061_));
 sky130_fd_sc_hd__o22a_1 _3117_ (.A1(net345),
    .A2(_1751_),
    .B1(_1753_),
    .B2(net400),
    .X(_0062_));
 sky130_fd_sc_hd__a22o_1 _3118_ (.A1(net268),
    .A2(net180),
    .B1(net116),
    .B2(net1088),
    .X(_0063_));
 sky130_fd_sc_hd__a22o_1 _3119_ (.A1(net261),
    .A2(net181),
    .B1(net116),
    .B2(net2240),
    .X(_0064_));
 sky130_fd_sc_hd__o22a_1 _3120_ (.A1(net260),
    .A2(_1751_),
    .B1(_1753_),
    .B2(net598),
    .X(_0065_));
 sky130_fd_sc_hd__o22a_1 _3121_ (.A1(net257),
    .A2(_1751_),
    .B1(_1753_),
    .B2(net652),
    .X(_0066_));
 sky130_fd_sc_hd__a22o_1 _3122_ (.A1(net255),
    .A2(net181),
    .B1(net117),
    .B2(net1098),
    .X(_0067_));
 sky130_fd_sc_hd__a22o_1 _3123_ (.A1(net253),
    .A2(net180),
    .B1(net116),
    .B2(net1572),
    .X(_0068_));
 sky130_fd_sc_hd__a22o_1 _3124_ (.A1(net251),
    .A2(net181),
    .B1(net116),
    .B2(net2354),
    .X(_0069_));
 sky130_fd_sc_hd__a22o_1 _3125_ (.A1(net249),
    .A2(net180),
    .B1(net116),
    .B2(net2008),
    .X(_0070_));
 sky130_fd_sc_hd__a22o_1 _3126_ (.A1(net225),
    .A2(net181),
    .B1(net117),
    .B2(net836),
    .X(_0071_));
 sky130_fd_sc_hd__a22o_1 _3127_ (.A1(net363),
    .A2(net180),
    .B1(net116),
    .B2(net1756),
    .X(_0072_));
 sky130_fd_sc_hd__a22o_1 _3128_ (.A1(net361),
    .A2(net181),
    .B1(net117),
    .B2(net710),
    .X(_0073_));
 sky130_fd_sc_hd__a22o_1 _3129_ (.A1(net359),
    .A2(net180),
    .B1(net117),
    .B2(net1666),
    .X(_0074_));
 sky130_fd_sc_hd__a22o_1 _3130_ (.A1(net357),
    .A2(net181),
    .B1(net117),
    .B2(net1888),
    .X(_0075_));
 sky130_fd_sc_hd__a22o_1 _3131_ (.A1(net355),
    .A2(net181),
    .B1(net117),
    .B2(net1004),
    .X(_0076_));
 sky130_fd_sc_hd__a22o_1 _3132_ (.A1(net353),
    .A2(net181),
    .B1(net117),
    .B2(net1748),
    .X(_0077_));
 sky130_fd_sc_hd__a22o_1 _3133_ (.A1(net351),
    .A2(net180),
    .B1(net117),
    .B2(net1150),
    .X(_0078_));
 sky130_fd_sc_hd__a22o_1 _3134_ (.A1(net349),
    .A2(net180),
    .B1(net116),
    .B2(net1826),
    .X(_0079_));
 sky130_fd_sc_hd__a22o_1 _3135_ (.A1(net347),
    .A2(net181),
    .B1(net117),
    .B2(net936),
    .X(_0080_));
 sky130_fd_sc_hd__a22o_1 _3136_ (.A1(net316),
    .A2(net181),
    .B1(net117),
    .B2(net1944),
    .X(_0081_));
 sky130_fd_sc_hd__a22o_1 _3137_ (.A1(net314),
    .A2(net180),
    .B1(net116),
    .B2(net910),
    .X(_0082_));
 sky130_fd_sc_hd__a22o_1 _3138_ (.A1(net312),
    .A2(net180),
    .B1(net116),
    .B2(net1718),
    .X(_0083_));
 sky130_fd_sc_hd__a22o_1 _3139_ (.A1(net310),
    .A2(net180),
    .B1(net116),
    .B2(net1522),
    .X(_0084_));
 sky130_fd_sc_hd__a22o_1 _3140_ (.A1(net308),
    .A2(net180),
    .B1(net116),
    .B2(net1564),
    .X(_0085_));
 sky130_fd_sc_hd__a22o_1 _3141_ (.A1(net306),
    .A2(net180),
    .B1(net116),
    .B2(net2244),
    .X(_0086_));
 sky130_fd_sc_hd__a22o_1 _3142_ (.A1(net304),
    .A2(net180),
    .B1(net116),
    .B2(net1900),
    .X(_0087_));
 sky130_fd_sc_hd__a22o_1 _3143_ (.A1(net301),
    .A2(net181),
    .B1(net117),
    .B2(net932),
    .X(_0088_));
 sky130_fd_sc_hd__a22o_1 _3144_ (.A1(net299),
    .A2(net181),
    .B1(net116),
    .B2(net1102),
    .X(_0089_));
 sky130_fd_sc_hd__a22o_1 _3145_ (.A1(net297),
    .A2(net180),
    .B1(net116),
    .B2(net1218),
    .X(_0090_));
 sky130_fd_sc_hd__a22o_1 _3146_ (.A1(net266),
    .A2(net180),
    .B1(net116),
    .B2(net1120),
    .X(_0091_));
 sky130_fd_sc_hd__a22o_1 _3147_ (.A1(net265),
    .A2(net181),
    .B1(net117),
    .B2(net1838),
    .X(_0092_));
 sky130_fd_sc_hd__and4b_1 _3148_ (.A_N(net292),
    .B(net340),
    .C(net216),
    .D(_1741_),
    .X(_1754_));
 sky130_fd_sc_hd__nand2_2 _3149_ (.A(_1670_),
    .B(_1741_),
    .Y(_1755_));
 sky130_fd_sc_hd__nor2_1 _3150_ (.A(net368),
    .B(net179),
    .Y(_1756_));
 sky130_fd_sc_hd__or2_2 _3151_ (.A(net366),
    .B(net179),
    .X(_1757_));
 sky130_fd_sc_hd__o22a_1 _3152_ (.A1(net227),
    .A2(_1755_),
    .B1(_1757_),
    .B2(net494),
    .X(_0093_));
 sky130_fd_sc_hd__o22a_1 _3153_ (.A1(net346),
    .A2(_1755_),
    .B1(_1757_),
    .B2(net374),
    .X(_0094_));
 sky130_fd_sc_hd__a22o_1 _3154_ (.A1(net269),
    .A2(net178),
    .B1(net114),
    .B2(net1282),
    .X(_0095_));
 sky130_fd_sc_hd__a22o_1 _3155_ (.A1(net261),
    .A2(net179),
    .B1(net115),
    .B2(net1182),
    .X(_0096_));
 sky130_fd_sc_hd__o22a_1 _3156_ (.A1(net259),
    .A2(_1755_),
    .B1(_1757_),
    .B2(net386),
    .X(_0097_));
 sky130_fd_sc_hd__o22a_1 _3157_ (.A1(net258),
    .A2(_1755_),
    .B1(_1757_),
    .B2(net780),
    .X(_0098_));
 sky130_fd_sc_hd__a22o_1 _3158_ (.A1(net256),
    .A2(net179),
    .B1(net115),
    .B2(net1146),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _3159_ (.A1(net254),
    .A2(net178),
    .B1(net114),
    .B2(net760),
    .X(_0100_));
 sky130_fd_sc_hd__a22o_1 _3160_ (.A1(net252),
    .A2(net178),
    .B1(net114),
    .B2(net1210),
    .X(_0101_));
 sky130_fd_sc_hd__a22o_1 _3161_ (.A1(net250),
    .A2(net178),
    .B1(net114),
    .B2(net960),
    .X(_0102_));
 sky130_fd_sc_hd__a22o_1 _3162_ (.A1(net226),
    .A2(net179),
    .B1(net115),
    .B2(net756),
    .X(_0103_));
 sky130_fd_sc_hd__a22o_1 _3163_ (.A1(net364),
    .A2(net178),
    .B1(net114),
    .B2(net1978),
    .X(_0104_));
 sky130_fd_sc_hd__a22o_1 _3164_ (.A1(net362),
    .A2(net179),
    .B1(net115),
    .B2(net844),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _3165_ (.A1(net360),
    .A2(net178),
    .B1(net114),
    .B2(net1226),
    .X(_0106_));
 sky130_fd_sc_hd__a22o_1 _3166_ (.A1(net358),
    .A2(net179),
    .B1(net115),
    .B2(net1482),
    .X(_0107_));
 sky130_fd_sc_hd__a22o_1 _3167_ (.A1(net356),
    .A2(net178),
    .B1(net114),
    .B2(net748),
    .X(_0108_));
 sky130_fd_sc_hd__a22o_1 _3168_ (.A1(net354),
    .A2(net179),
    .B1(net115),
    .B2(net1206),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _3169_ (.A1(net352),
    .A2(net179),
    .B1(net115),
    .B2(net1374),
    .X(_0110_));
 sky130_fd_sc_hd__a22o_1 _3170_ (.A1(net350),
    .A2(net178),
    .B1(net114),
    .B2(net1998),
    .X(_0111_));
 sky130_fd_sc_hd__a22o_1 _3171_ (.A1(net348),
    .A2(net179),
    .B1(net115),
    .B2(net1066),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _3172_ (.A1(net317),
    .A2(net179),
    .B1(net115),
    .B2(net2190),
    .X(_0113_));
 sky130_fd_sc_hd__a22o_1 _3173_ (.A1(net315),
    .A2(net178),
    .B1(net114),
    .B2(net1440),
    .X(_0114_));
 sky130_fd_sc_hd__a22o_1 _3174_ (.A1(net313),
    .A2(net178),
    .B1(net114),
    .B2(net1732),
    .X(_0115_));
 sky130_fd_sc_hd__a22o_1 _3175_ (.A1(net311),
    .A2(net178),
    .B1(net114),
    .B2(net1064),
    .X(_0116_));
 sky130_fd_sc_hd__a22o_1 _3176_ (.A1(net309),
    .A2(net178),
    .B1(net114),
    .B2(net676),
    .X(_0117_));
 sky130_fd_sc_hd__a22o_1 _3177_ (.A1(net307),
    .A2(net179),
    .B1(net115),
    .B2(net1032),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_1 _3178_ (.A1(net303),
    .A2(net178),
    .B1(net114),
    .B2(net1854),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _3179_ (.A1(net302),
    .A2(net179),
    .B1(net115),
    .B2(net834),
    .X(_0120_));
 sky130_fd_sc_hd__a22o_1 _3180_ (.A1(net300),
    .A2(net178),
    .B1(net114),
    .B2(net754),
    .X(_0121_));
 sky130_fd_sc_hd__a22o_1 _3181_ (.A1(net298),
    .A2(net178),
    .B1(net114),
    .B2(net1192),
    .X(_0122_));
 sky130_fd_sc_hd__a22o_1 _3182_ (.A1(net267),
    .A2(net178),
    .B1(net114),
    .B2(net788),
    .X(_0123_));
 sky130_fd_sc_hd__a22o_1 _3183_ (.A1(net264),
    .A2(net179),
    .B1(net115),
    .B2(net1312),
    .X(_0124_));
 sky130_fd_sc_hd__and3_1 _3184_ (.A(net216),
    .B(_1686_),
    .C(_1693_),
    .X(_1758_));
 sky130_fd_sc_hd__nand2_1 _3185_ (.A(_1686_),
    .B(_1694_),
    .Y(_1759_));
 sky130_fd_sc_hd__nor2_1 _3186_ (.A(net369),
    .B(net176),
    .Y(_1760_));
 sky130_fd_sc_hd__or2_2 _3187_ (.A(net368),
    .B(net176),
    .X(_1761_));
 sky130_fd_sc_hd__o22a_1 _3188_ (.A1(net227),
    .A2(_1759_),
    .B1(_1761_),
    .B2(net574),
    .X(_0125_));
 sky130_fd_sc_hd__o22a_1 _3189_ (.A1(net346),
    .A2(_1759_),
    .B1(_1761_),
    .B2(net540),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _3190_ (.A1(net269),
    .A2(net177),
    .B1(net112),
    .B2(net1444),
    .X(_0127_));
 sky130_fd_sc_hd__a22o_1 _3191_ (.A1(net261),
    .A2(net176),
    .B1(net113),
    .B2(net946),
    .X(_0128_));
 sky130_fd_sc_hd__o22a_1 _3192_ (.A1(net259),
    .A2(_1759_),
    .B1(_1761_),
    .B2(net470),
    .X(_0129_));
 sky130_fd_sc_hd__o22a_1 _3193_ (.A1(net258),
    .A2(_1759_),
    .B1(_1761_),
    .B2(net554),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _3194_ (.A1(net256),
    .A2(net176),
    .B1(net113),
    .B2(net2172),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _3195_ (.A1(net254),
    .A2(net177),
    .B1(net112),
    .B2(net2044),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _3196_ (.A1(net252),
    .A2(net176),
    .B1(net112),
    .B2(net2048),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _3197_ (.A1(net250),
    .A2(net177),
    .B1(net112),
    .B2(net1388),
    .X(_0134_));
 sky130_fd_sc_hd__a22o_1 _3198_ (.A1(net226),
    .A2(net176),
    .B1(net113),
    .B2(net1630),
    .X(_0135_));
 sky130_fd_sc_hd__a22o_1 _3199_ (.A1(net364),
    .A2(net177),
    .B1(net112),
    .B2(net1508),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _3200_ (.A1(net362),
    .A2(net176),
    .B1(net113),
    .B2(net1036),
    .X(_0137_));
 sky130_fd_sc_hd__a22o_1 _3201_ (.A1(net360),
    .A2(net177),
    .B1(net112),
    .B2(net1236),
    .X(_0138_));
 sky130_fd_sc_hd__a22o_1 _3202_ (.A1(net358),
    .A2(net176),
    .B1(net113),
    .B2(net1018),
    .X(_0139_));
 sky130_fd_sc_hd__a22o_1 _3203_ (.A1(net356),
    .A2(net176),
    .B1(net113),
    .B2(net694),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _3204_ (.A1(net354),
    .A2(net177),
    .B1(net113),
    .B2(net1846),
    .X(_0141_));
 sky130_fd_sc_hd__a22o_1 _3205_ (.A1(net352),
    .A2(net176),
    .B1(net113),
    .B2(net940),
    .X(_0142_));
 sky130_fd_sc_hd__a22o_1 _3206_ (.A1(net350),
    .A2(net177),
    .B1(net112),
    .B2(net2148),
    .X(_0143_));
 sky130_fd_sc_hd__a22o_1 _3207_ (.A1(net348),
    .A2(net176),
    .B1(net113),
    .B2(net878),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_1 _3208_ (.A1(net317),
    .A2(net176),
    .B1(net113),
    .B2(net1250),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _3209_ (.A1(net315),
    .A2(net176),
    .B1(net112),
    .B2(net1506),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _3210_ (.A1(net313),
    .A2(net177),
    .B1(net112),
    .B2(net1326),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_1 _3211_ (.A1(net311),
    .A2(net177),
    .B1(net112),
    .B2(net1196),
    .X(_0148_));
 sky130_fd_sc_hd__a22o_1 _3212_ (.A1(net309),
    .A2(net177),
    .B1(net112),
    .B2(net2156),
    .X(_0149_));
 sky130_fd_sc_hd__a22o_1 _3213_ (.A1(net307),
    .A2(net177),
    .B1(net112),
    .B2(net2272),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_1 _3214_ (.A1(net303),
    .A2(net176),
    .B1(net112),
    .B2(net1136),
    .X(_0151_));
 sky130_fd_sc_hd__a22o_1 _3215_ (.A1(net302),
    .A2(net176),
    .B1(net113),
    .B2(net1462),
    .X(_0152_));
 sky130_fd_sc_hd__a22o_1 _3216_ (.A1(net300),
    .A2(net177),
    .B1(net112),
    .B2(net608),
    .X(_0153_));
 sky130_fd_sc_hd__a22o_1 _3217_ (.A1(net298),
    .A2(net177),
    .B1(net112),
    .B2(net2066),
    .X(_0154_));
 sky130_fd_sc_hd__a22o_1 _3218_ (.A1(net267),
    .A2(net177),
    .B1(net112),
    .B2(net1380),
    .X(_0155_));
 sky130_fd_sc_hd__a22o_1 _3219_ (.A1(net264),
    .A2(net176),
    .B1(net113),
    .B2(net670),
    .X(_0156_));
 sky130_fd_sc_hd__and4_1 _3220_ (.A(net283),
    .B(net331),
    .C(_1028_),
    .D(net217),
    .X(_1762_));
 sky130_fd_sc_hd__nand2_1 _3221_ (.A(_1028_),
    .B(_1687_),
    .Y(_1763_));
 sky130_fd_sc_hd__nor2_1 _3222_ (.A(net365),
    .B(net175),
    .Y(_1764_));
 sky130_fd_sc_hd__or2_2 _3223_ (.A(net365),
    .B(net175),
    .X(_1765_));
 sky130_fd_sc_hd__o22a_1 _3224_ (.A1(net228),
    .A2(_1763_),
    .B1(_1765_),
    .B2(net430),
    .X(_0157_));
 sky130_fd_sc_hd__o22a_1 _3225_ (.A1(net345),
    .A2(_1763_),
    .B1(_1765_),
    .B2(net408),
    .X(_0158_));
 sky130_fd_sc_hd__a22o_1 _3226_ (.A1(net268),
    .A2(net174),
    .B1(net110),
    .B2(net642),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _3227_ (.A1(net263),
    .A2(net175),
    .B1(net111),
    .B2(net848),
    .X(_0160_));
 sky130_fd_sc_hd__o22a_1 _3228_ (.A1(net260),
    .A2(_1763_),
    .B1(_1765_),
    .B2(net450),
    .X(_0161_));
 sky130_fd_sc_hd__o22a_1 _3229_ (.A1(net257),
    .A2(_1763_),
    .B1(_1765_),
    .B2(net530),
    .X(_0162_));
 sky130_fd_sc_hd__a22o_1 _3230_ (.A1(net255),
    .A2(net175),
    .B1(net111),
    .B2(net734),
    .X(_0163_));
 sky130_fd_sc_hd__a22o_1 _3231_ (.A1(net253),
    .A2(net174),
    .B1(net110),
    .B2(net808),
    .X(_0164_));
 sky130_fd_sc_hd__a22o_1 _3232_ (.A1(net251),
    .A2(net175),
    .B1(net110),
    .B2(net2242),
    .X(_0165_));
 sky130_fd_sc_hd__a22o_1 _3233_ (.A1(net249),
    .A2(net174),
    .B1(net110),
    .B2(net750),
    .X(_0166_));
 sky130_fd_sc_hd__a22o_1 _3234_ (.A1(net225),
    .A2(net175),
    .B1(net111),
    .B2(net966),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _3235_ (.A1(net363),
    .A2(net174),
    .B1(net110),
    .B2(net1794),
    .X(_0168_));
 sky130_fd_sc_hd__a22o_1 _3236_ (.A1(net361),
    .A2(net175),
    .B1(net111),
    .B2(net1318),
    .X(_0169_));
 sky130_fd_sc_hd__a22o_1 _3237_ (.A1(net359),
    .A2(net174),
    .B1(net110),
    .B2(net2340),
    .X(_0170_));
 sky130_fd_sc_hd__a22o_1 _3238_ (.A1(net357),
    .A2(net175),
    .B1(net111),
    .B2(net1472),
    .X(_0171_));
 sky130_fd_sc_hd__a22o_1 _3239_ (.A1(net355),
    .A2(net174),
    .B1(net110),
    .B2(net1204),
    .X(_0172_));
 sky130_fd_sc_hd__a22o_1 _3240_ (.A1(net353),
    .A2(net175),
    .B1(net111),
    .B2(net816),
    .X(_0173_));
 sky130_fd_sc_hd__a22o_1 _3241_ (.A1(net351),
    .A2(net175),
    .B1(net111),
    .B2(net2408),
    .X(_0174_));
 sky130_fd_sc_hd__a22o_1 _3242_ (.A1(net349),
    .A2(net174),
    .B1(net111),
    .B2(net1418),
    .X(_0175_));
 sky130_fd_sc_hd__a22o_1 _3243_ (.A1(net347),
    .A2(net175),
    .B1(net111),
    .B2(net800),
    .X(_0176_));
 sky130_fd_sc_hd__a22o_1 _3244_ (.A1(net316),
    .A2(net175),
    .B1(net111),
    .B2(net2296),
    .X(_0177_));
 sky130_fd_sc_hd__a22o_1 _3245_ (.A1(net314),
    .A2(net174),
    .B1(net110),
    .B2(net1260),
    .X(_0178_));
 sky130_fd_sc_hd__a22o_1 _3246_ (.A1(net312),
    .A2(net174),
    .B1(net110),
    .B2(net1248),
    .X(_0179_));
 sky130_fd_sc_hd__a22o_1 _3247_ (.A1(net310),
    .A2(net174),
    .B1(net110),
    .B2(net1722),
    .X(_0180_));
 sky130_fd_sc_hd__a22o_1 _3248_ (.A1(net308),
    .A2(net174),
    .B1(net110),
    .B2(net888),
    .X(_0181_));
 sky130_fd_sc_hd__a22o_1 _3249_ (.A1(net306),
    .A2(net174),
    .B1(net110),
    .B2(net1686),
    .X(_0182_));
 sky130_fd_sc_hd__a22o_1 _3250_ (.A1(net305),
    .A2(net174),
    .B1(net110),
    .B2(net1520),
    .X(_0183_));
 sky130_fd_sc_hd__a22o_1 _3251_ (.A1(net301),
    .A2(net175),
    .B1(net111),
    .B2(net1056),
    .X(_0184_));
 sky130_fd_sc_hd__a22o_1 _3252_ (.A1(net299),
    .A2(net174),
    .B1(net110),
    .B2(net1576),
    .X(_0185_));
 sky130_fd_sc_hd__a22o_1 _3253_ (.A1(net297),
    .A2(net174),
    .B1(net110),
    .B2(net2134),
    .X(_0186_));
 sky130_fd_sc_hd__a22o_1 _3254_ (.A1(net266),
    .A2(net174),
    .B1(net110),
    .B2(net872),
    .X(_0187_));
 sky130_fd_sc_hd__a22o_1 _3255_ (.A1(net265),
    .A2(net175),
    .B1(net111),
    .B2(net718),
    .X(_0188_));
 sky130_fd_sc_hd__and4_1 _3256_ (.A(net292),
    .B(net340),
    .C(net216),
    .D(_1741_),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_2 _3257_ (.A(_1687_),
    .B(_1741_),
    .Y(_1767_));
 sky130_fd_sc_hd__nor2_1 _3258_ (.A(net368),
    .B(net173),
    .Y(_1768_));
 sky130_fd_sc_hd__or2_2 _3259_ (.A(net366),
    .B(net173),
    .X(_1769_));
 sky130_fd_sc_hd__o22a_1 _3260_ (.A1(net227),
    .A2(_1767_),
    .B1(_1769_),
    .B2(net884),
    .X(_0189_));
 sky130_fd_sc_hd__o22a_1 _3261_ (.A1(net346),
    .A2(_1767_),
    .B1(_1769_),
    .B2(net426),
    .X(_0190_));
 sky130_fd_sc_hd__a22o_1 _3262_ (.A1(net269),
    .A2(net172),
    .B1(net108),
    .B2(net1922),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _3263_ (.A1(net262),
    .A2(net173),
    .B1(net109),
    .B2(net648),
    .X(_0192_));
 sky130_fd_sc_hd__o22a_1 _3264_ (.A1(net259),
    .A2(_1767_),
    .B1(_1769_),
    .B2(net462),
    .X(_0193_));
 sky130_fd_sc_hd__o22a_1 _3265_ (.A1(net258),
    .A2(_1767_),
    .B1(_1769_),
    .B2(net406),
    .X(_0194_));
 sky130_fd_sc_hd__a22o_1 _3266_ (.A1(net256),
    .A2(net173),
    .B1(net109),
    .B2(net990),
    .X(_0195_));
 sky130_fd_sc_hd__a22o_1 _3267_ (.A1(net254),
    .A2(net172),
    .B1(net108),
    .B2(net1620),
    .X(_0196_));
 sky130_fd_sc_hd__a22o_1 _3268_ (.A1(net252),
    .A2(net172),
    .B1(net108),
    .B2(net1122),
    .X(_0197_));
 sky130_fd_sc_hd__a22o_1 _3269_ (.A1(net250),
    .A2(net172),
    .B1(net108),
    .B2(net1314),
    .X(_0198_));
 sky130_fd_sc_hd__a22o_1 _3270_ (.A1(net226),
    .A2(net173),
    .B1(net109),
    .B2(net2058),
    .X(_0199_));
 sky130_fd_sc_hd__a22o_1 _3271_ (.A1(net364),
    .A2(net172),
    .B1(net108),
    .B2(net1914),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _3272_ (.A1(net362),
    .A2(net173),
    .B1(net109),
    .B2(net1586),
    .X(_0201_));
 sky130_fd_sc_hd__a22o_1 _3273_ (.A1(net360),
    .A2(net172),
    .B1(net108),
    .B2(net672),
    .X(_0202_));
 sky130_fd_sc_hd__a22o_1 _3274_ (.A1(net358),
    .A2(net173),
    .B1(net109),
    .B2(net942),
    .X(_0203_));
 sky130_fd_sc_hd__a22o_1 _3275_ (.A1(net356),
    .A2(net172),
    .B1(net108),
    .B2(net908),
    .X(_0204_));
 sky130_fd_sc_hd__a22o_1 _3276_ (.A1(net354),
    .A2(net173),
    .B1(net109),
    .B2(net1456),
    .X(_0205_));
 sky130_fd_sc_hd__a22o_1 _3277_ (.A1(net352),
    .A2(net173),
    .B1(net109),
    .B2(net2178),
    .X(_0206_));
 sky130_fd_sc_hd__a22o_1 _3278_ (.A1(net350),
    .A2(net172),
    .B1(net108),
    .B2(net1770),
    .X(_0207_));
 sky130_fd_sc_hd__a22o_1 _3279_ (.A1(net348),
    .A2(net173),
    .B1(net109),
    .B2(net1988),
    .X(_0208_));
 sky130_fd_sc_hd__a22o_1 _3280_ (.A1(net317),
    .A2(net173),
    .B1(net109),
    .B2(net952),
    .X(_0209_));
 sky130_fd_sc_hd__a22o_1 _3281_ (.A1(net315),
    .A2(net172),
    .B1(net108),
    .B2(net1096),
    .X(_0210_));
 sky130_fd_sc_hd__a22o_1 _3282_ (.A1(net313),
    .A2(net172),
    .B1(net108),
    .B2(net1606),
    .X(_0211_));
 sky130_fd_sc_hd__a22o_1 _3283_ (.A1(net311),
    .A2(net172),
    .B1(net108),
    .B2(net2336),
    .X(_0212_));
 sky130_fd_sc_hd__a22o_1 _3284_ (.A1(net309),
    .A2(net172),
    .B1(net108),
    .B2(net906),
    .X(_0213_));
 sky130_fd_sc_hd__a22o_1 _3285_ (.A1(net307),
    .A2(net173),
    .B1(net109),
    .B2(net1106),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_1 _3286_ (.A1(net303),
    .A2(net172),
    .B1(net108),
    .B2(net1172),
    .X(_0215_));
 sky130_fd_sc_hd__a22o_1 _3287_ (.A1(net302),
    .A2(net173),
    .B1(net109),
    .B2(net592),
    .X(_0216_));
 sky130_fd_sc_hd__a22o_1 _3288_ (.A1(net300),
    .A2(net172),
    .B1(net108),
    .B2(net1094),
    .X(_0217_));
 sky130_fd_sc_hd__a22o_1 _3289_ (.A1(net298),
    .A2(net172),
    .B1(net108),
    .B2(net1844),
    .X(_0218_));
 sky130_fd_sc_hd__a22o_1 _3290_ (.A1(net267),
    .A2(net172),
    .B1(net108),
    .B2(net1870),
    .X(_0219_));
 sky130_fd_sc_hd__a22o_1 _3291_ (.A1(net264),
    .A2(net173),
    .B1(net109),
    .B2(net1142),
    .X(_0220_));
 sky130_fd_sc_hd__and3_1 _3292_ (.A(_1027_),
    .B(net217),
    .C(_1675_),
    .X(_1770_));
 sky130_fd_sc_hd__nand2_1 _3293_ (.A(_1027_),
    .B(_1676_),
    .Y(_1771_));
 sky130_fd_sc_hd__nor2_1 _3294_ (.A(net367),
    .B(net171),
    .Y(_1772_));
 sky130_fd_sc_hd__or2_2 _3295_ (.A(net366),
    .B(net171),
    .X(_1773_));
 sky130_fd_sc_hd__o22a_1 _3296_ (.A1(net228),
    .A2(_1771_),
    .B1(_1773_),
    .B2(net498),
    .X(_0221_));
 sky130_fd_sc_hd__o22a_1 _3297_ (.A1(net345),
    .A2(_1771_),
    .B1(_1773_),
    .B2(net432),
    .X(_0222_));
 sky130_fd_sc_hd__a22o_1 _3298_ (.A1(net268),
    .A2(net170),
    .B1(net106),
    .B2(net1822),
    .X(_0223_));
 sky130_fd_sc_hd__a22o_1 _3299_ (.A1(net263),
    .A2(net171),
    .B1(net107),
    .B2(net1304),
    .X(_0224_));
 sky130_fd_sc_hd__o22a_1 _3300_ (.A1(net260),
    .A2(_1771_),
    .B1(_1773_),
    .B2(net434),
    .X(_0225_));
 sky130_fd_sc_hd__o22a_1 _3301_ (.A1(net257),
    .A2(_1771_),
    .B1(_1773_),
    .B2(net514),
    .X(_0226_));
 sky130_fd_sc_hd__a22o_1 _3302_ (.A1(net255),
    .A2(net171),
    .B1(net107),
    .B2(net798),
    .X(_0227_));
 sky130_fd_sc_hd__a22o_1 _3303_ (.A1(net253),
    .A2(net170),
    .B1(net106),
    .B2(net1166),
    .X(_0228_));
 sky130_fd_sc_hd__a22o_1 _3304_ (.A1(net251),
    .A2(net171),
    .B1(net107),
    .B2(net2384),
    .X(_0229_));
 sky130_fd_sc_hd__a22o_1 _3305_ (.A1(net249),
    .A2(net170),
    .B1(net106),
    .B2(net1828),
    .X(_0230_));
 sky130_fd_sc_hd__a22o_1 _3306_ (.A1(net225),
    .A2(net171),
    .B1(net107),
    .B2(net2164),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _3307_ (.A1(net363),
    .A2(net170),
    .B1(net106),
    .B2(net1514),
    .X(_0232_));
 sky130_fd_sc_hd__a22o_1 _3308_ (.A1(net361),
    .A2(net171),
    .B1(net107),
    .B2(net2316),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _3309_ (.A1(net359),
    .A2(net170),
    .B1(net106),
    .B2(net2092),
    .X(_0234_));
 sky130_fd_sc_hd__a22o_1 _3310_ (.A1(net357),
    .A2(net171),
    .B1(net107),
    .B2(net2128),
    .X(_0235_));
 sky130_fd_sc_hd__a22o_1 _3311_ (.A1(net355),
    .A2(net170),
    .B1(net106),
    .B2(net1238),
    .X(_0236_));
 sky130_fd_sc_hd__a22o_1 _3312_ (.A1(net353),
    .A2(net171),
    .B1(net107),
    .B2(net1276),
    .X(_0237_));
 sky130_fd_sc_hd__a22o_1 _3313_ (.A1(net351),
    .A2(net171),
    .B1(net107),
    .B2(net698),
    .X(_0238_));
 sky130_fd_sc_hd__a22o_1 _3314_ (.A1(net349),
    .A2(net170),
    .B1(net106),
    .B2(net822),
    .X(_0239_));
 sky130_fd_sc_hd__a22o_1 _3315_ (.A1(net347),
    .A2(net171),
    .B1(net107),
    .B2(net1636),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _3316_ (.A1(net316),
    .A2(net171),
    .B1(net107),
    .B2(net1758),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_1 _3317_ (.A1(net314),
    .A2(net170),
    .B1(net106),
    .B2(net826),
    .X(_0242_));
 sky130_fd_sc_hd__a22o_1 _3318_ (.A1(net312),
    .A2(net170),
    .B1(net106),
    .B2(net1816),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _3319_ (.A1(net310),
    .A2(net170),
    .B1(net106),
    .B2(net1164),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _3320_ (.A1(net308),
    .A2(net170),
    .B1(net106),
    .B2(net2388),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _3321_ (.A1(net306),
    .A2(net170),
    .B1(net106),
    .B2(net2174),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_1 _3322_ (.A1(net305),
    .A2(net170),
    .B1(net106),
    .B2(net2026),
    .X(_0247_));
 sky130_fd_sc_hd__a22o_1 _3323_ (.A1(net301),
    .A2(net171),
    .B1(net107),
    .B2(net1766),
    .X(_0248_));
 sky130_fd_sc_hd__a22o_1 _3324_ (.A1(net299),
    .A2(net170),
    .B1(net106),
    .B2(net1976),
    .X(_0249_));
 sky130_fd_sc_hd__a22o_1 _3325_ (.A1(net297),
    .A2(net170),
    .B1(net106),
    .B2(net2284),
    .X(_0250_));
 sky130_fd_sc_hd__a22o_1 _3326_ (.A1(net266),
    .A2(net170),
    .B1(net106),
    .B2(net1588),
    .X(_0251_));
 sky130_fd_sc_hd__a22o_1 _3327_ (.A1(net265),
    .A2(net171),
    .B1(net107),
    .B2(net2346),
    .X(_0252_));
 sky130_fd_sc_hd__and3_1 _3328_ (.A(_1669_),
    .B(_1693_),
    .C(_1711_),
    .X(_1774_));
 sky130_fd_sc_hd__nand2_1 _3329_ (.A(_1694_),
    .B(_1711_),
    .Y(_1775_));
 sky130_fd_sc_hd__nor2_1 _3330_ (.A(net369),
    .B(net169),
    .Y(_1776_));
 sky130_fd_sc_hd__or2_2 _3331_ (.A(net368),
    .B(net169),
    .X(_1777_));
 sky130_fd_sc_hd__o22a_1 _3332_ (.A1(net227),
    .A2(_1775_),
    .B1(_1777_),
    .B2(net382),
    .X(_0253_));
 sky130_fd_sc_hd__o22a_1 _3333_ (.A1(net346),
    .A2(_1775_),
    .B1(_1777_),
    .B2(net768),
    .X(_0254_));
 sky130_fd_sc_hd__a22o_1 _3334_ (.A1(net269),
    .A2(net168),
    .B1(net104),
    .B2(net644),
    .X(_0255_));
 sky130_fd_sc_hd__a22o_1 _3335_ (.A1(net262),
    .A2(net169),
    .B1(net105),
    .B2(net1368),
    .X(_0256_));
 sky130_fd_sc_hd__o22a_1 _3336_ (.A1(net259),
    .A2(_1775_),
    .B1(_1777_),
    .B2(net370),
    .X(_0257_));
 sky130_fd_sc_hd__o22a_1 _3337_ (.A1(net258),
    .A2(_1775_),
    .B1(_1777_),
    .B2(net562),
    .X(_0258_));
 sky130_fd_sc_hd__a22o_1 _3338_ (.A1(net256),
    .A2(net169),
    .B1(net105),
    .B2(net1538),
    .X(_0259_));
 sky130_fd_sc_hd__a22o_1 _3339_ (.A1(net254),
    .A2(net168),
    .B1(net104),
    .B2(net1040),
    .X(_0260_));
 sky130_fd_sc_hd__a22o_1 _3340_ (.A1(net252),
    .A2(net168),
    .B1(net104),
    .B2(net1924),
    .X(_0261_));
 sky130_fd_sc_hd__a22o_1 _3341_ (.A1(net250),
    .A2(net168),
    .B1(net104),
    .B2(net1006),
    .X(_0262_));
 sky130_fd_sc_hd__a22o_1 _3342_ (.A1(net226),
    .A2(net169),
    .B1(net105),
    .B2(net1640),
    .X(_0263_));
 sky130_fd_sc_hd__a22o_1 _3343_ (.A1(net364),
    .A2(net168),
    .B1(net104),
    .B2(net1494),
    .X(_0264_));
 sky130_fd_sc_hd__a22o_1 _3344_ (.A1(net362),
    .A2(net169),
    .B1(net105),
    .B2(net1706),
    .X(_0265_));
 sky130_fd_sc_hd__a22o_1 _3345_ (.A1(net360),
    .A2(net169),
    .B1(net104),
    .B2(net830),
    .X(_0266_));
 sky130_fd_sc_hd__a22o_1 _3346_ (.A1(net358),
    .A2(net169),
    .B1(net105),
    .B2(net2230),
    .X(_0267_));
 sky130_fd_sc_hd__a22o_1 _3347_ (.A1(net356),
    .A2(net168),
    .B1(net105),
    .B2(net978),
    .X(_0268_));
 sky130_fd_sc_hd__a22o_1 _3348_ (.A1(net354),
    .A2(net169),
    .B1(net105),
    .B2(net1452),
    .X(_0269_));
 sky130_fd_sc_hd__a22o_1 _3349_ (.A1(net352),
    .A2(net169),
    .B1(net105),
    .B2(net1768),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_1 _3350_ (.A1(net350),
    .A2(net168),
    .B1(net104),
    .B2(net1216),
    .X(_0271_));
 sky130_fd_sc_hd__a22o_1 _3351_ (.A1(net348),
    .A2(net169),
    .B1(net105),
    .B2(net1632),
    .X(_0272_));
 sky130_fd_sc_hd__a22o_1 _3352_ (.A1(net317),
    .A2(net169),
    .B1(net105),
    .B2(net1232),
    .X(_0273_));
 sky130_fd_sc_hd__a22o_1 _3353_ (.A1(net315),
    .A2(net168),
    .B1(net104),
    .B2(net974),
    .X(_0274_));
 sky130_fd_sc_hd__a22o_1 _3354_ (.A1(net313),
    .A2(net168),
    .B1(net104),
    .B2(net2210),
    .X(_0275_));
 sky130_fd_sc_hd__a22o_1 _3355_ (.A1(net311),
    .A2(net168),
    .B1(net104),
    .B2(net934),
    .X(_0276_));
 sky130_fd_sc_hd__a22o_1 _3356_ (.A1(net309),
    .A2(net168),
    .B1(net104),
    .B2(net1830),
    .X(_0277_));
 sky130_fd_sc_hd__a22o_1 _3357_ (.A1(net307),
    .A2(net168),
    .B1(net104),
    .B2(net2146),
    .X(_0278_));
 sky130_fd_sc_hd__a22o_1 _3358_ (.A1(net303),
    .A2(net168),
    .B1(net104),
    .B2(net1014),
    .X(_0279_));
 sky130_fd_sc_hd__a22o_1 _3359_ (.A1(net302),
    .A2(net169),
    .B1(net105),
    .B2(net1264),
    .X(_0280_));
 sky130_fd_sc_hd__a22o_1 _3360_ (.A1(net300),
    .A2(net168),
    .B1(net104),
    .B2(net2030),
    .X(_0281_));
 sky130_fd_sc_hd__a22o_1 _3361_ (.A1(net298),
    .A2(net168),
    .B1(net104),
    .B2(net2132),
    .X(_0282_));
 sky130_fd_sc_hd__a22o_1 _3362_ (.A1(net267),
    .A2(net168),
    .B1(net104),
    .B2(net922),
    .X(_0283_));
 sky130_fd_sc_hd__a22o_1 _3363_ (.A1(net264),
    .A2(net169),
    .B1(net105),
    .B2(net1034),
    .X(_0284_));
 sky130_fd_sc_hd__and4b_1 _3364_ (.A_N(net294),
    .B(net342),
    .C(_1669_),
    .D(_1711_),
    .X(_1778_));
 sky130_fd_sc_hd__nand2_2 _3365_ (.A(_1670_),
    .B(_1711_),
    .Y(_1779_));
 sky130_fd_sc_hd__nor2_1 _3366_ (.A(net369),
    .B(net166),
    .Y(_1780_));
 sky130_fd_sc_hd__or2_2 _3367_ (.A(net368),
    .B(net167),
    .X(_1781_));
 sky130_fd_sc_hd__o22a_1 _3368_ (.A1(net227),
    .A2(_1779_),
    .B1(_1781_),
    .B2(net378),
    .X(_0285_));
 sky130_fd_sc_hd__o22a_1 _3369_ (.A1(net346),
    .A2(_1779_),
    .B1(_1781_),
    .B2(net504),
    .X(_0286_));
 sky130_fd_sc_hd__a22o_1 _3370_ (.A1(net269),
    .A2(net166),
    .B1(net102),
    .B2(net2246),
    .X(_0287_));
 sky130_fd_sc_hd__a22o_1 _3371_ (.A1(net262),
    .A2(net167),
    .B1(net102),
    .B2(net1400),
    .X(_0288_));
 sky130_fd_sc_hd__o22a_1 _3372_ (.A1(net259),
    .A2(_1779_),
    .B1(_1781_),
    .B2(net436),
    .X(_0289_));
 sky130_fd_sc_hd__o22a_1 _3373_ (.A1(net258),
    .A2(_1779_),
    .B1(_1781_),
    .B2(net394),
    .X(_0290_));
 sky130_fd_sc_hd__a22o_1 _3374_ (.A1(net256),
    .A2(net167),
    .B1(net103),
    .B2(net1886),
    .X(_0291_));
 sky130_fd_sc_hd__a22o_1 _3375_ (.A1(net254),
    .A2(net166),
    .B1(net102),
    .B2(net1608),
    .X(_0292_));
 sky130_fd_sc_hd__a22o_1 _3376_ (.A1(net252),
    .A2(net166),
    .B1(net102),
    .B2(net1176),
    .X(_0293_));
 sky130_fd_sc_hd__a22o_1 _3377_ (.A1(net250),
    .A2(net166),
    .B1(net102),
    .B2(net584),
    .X(_0294_));
 sky130_fd_sc_hd__a22o_1 _3378_ (.A1(net226),
    .A2(net167),
    .B1(net103),
    .B2(net998),
    .X(_0295_));
 sky130_fd_sc_hd__a22o_1 _3379_ (.A1(net364),
    .A2(net166),
    .B1(net102),
    .B2(net1198),
    .X(_0296_));
 sky130_fd_sc_hd__a22o_1 _3380_ (.A1(net362),
    .A2(net167),
    .B1(net103),
    .B2(net1160),
    .X(_0297_));
 sky130_fd_sc_hd__a22o_1 _3381_ (.A1(net360),
    .A2(net167),
    .B1(net102),
    .B2(net784),
    .X(_0298_));
 sky130_fd_sc_hd__a22o_1 _3382_ (.A1(net358),
    .A2(net167),
    .B1(net103),
    .B2(net2176),
    .X(_0299_));
 sky130_fd_sc_hd__a22o_1 _3383_ (.A1(net356),
    .A2(net166),
    .B1(net103),
    .B2(net1028),
    .X(_0300_));
 sky130_fd_sc_hd__a22o_1 _3384_ (.A1(net354),
    .A2(net167),
    .B1(net103),
    .B2(net902),
    .X(_0301_));
 sky130_fd_sc_hd__a22o_1 _3385_ (.A1(net352),
    .A2(net167),
    .B1(net103),
    .B2(net2064),
    .X(_0302_));
 sky130_fd_sc_hd__a22o_1 _3386_ (.A1(net350),
    .A2(net166),
    .B1(net102),
    .B2(net776),
    .X(_0303_));
 sky130_fd_sc_hd__a22o_1 _3387_ (.A1(net348),
    .A2(net167),
    .B1(net103),
    .B2(net1780),
    .X(_0304_));
 sky130_fd_sc_hd__a22o_1 _3388_ (.A1(net317),
    .A2(net167),
    .B1(net103),
    .B2(net926),
    .X(_0305_));
 sky130_fd_sc_hd__a22o_1 _3389_ (.A1(net315),
    .A2(net166),
    .B1(net102),
    .B2(net1188),
    .X(_0306_));
 sky130_fd_sc_hd__a22o_1 _3390_ (.A1(net313),
    .A2(net167),
    .B1(net102),
    .B2(net1372),
    .X(_0307_));
 sky130_fd_sc_hd__a22o_1 _3391_ (.A1(net311),
    .A2(net166),
    .B1(net102),
    .B2(net2080),
    .X(_0308_));
 sky130_fd_sc_hd__a22o_1 _3392_ (.A1(net309),
    .A2(net166),
    .B1(net102),
    .B2(net1786),
    .X(_0309_));
 sky130_fd_sc_hd__a22o_1 _3393_ (.A1(net307),
    .A2(net166),
    .B1(net102),
    .B2(net1358),
    .X(_0310_));
 sky130_fd_sc_hd__a22o_1 _3394_ (.A1(net303),
    .A2(net166),
    .B1(net103),
    .B2(net1798),
    .X(_0311_));
 sky130_fd_sc_hd__a22o_1 _3395_ (.A1(net302),
    .A2(net167),
    .B1(net103),
    .B2(net988),
    .X(_0312_));
 sky130_fd_sc_hd__a22o_1 _3396_ (.A1(net300),
    .A2(net166),
    .B1(net102),
    .B2(net1712),
    .X(_0313_));
 sky130_fd_sc_hd__a22o_1 _3397_ (.A1(net298),
    .A2(net166),
    .B1(net102),
    .B2(net772),
    .X(_0314_));
 sky130_fd_sc_hd__a22o_1 _3398_ (.A1(net267),
    .A2(net166),
    .B1(net102),
    .B2(net1430),
    .X(_0315_));
 sky130_fd_sc_hd__a22o_1 _3399_ (.A1(net32),
    .A2(net167),
    .B1(net103),
    .B2(net1436),
    .X(_0316_));
 sky130_fd_sc_hd__and3_1 _3400_ (.A(net216),
    .B(_1693_),
    .C(_1732_),
    .X(_1782_));
 sky130_fd_sc_hd__nand2_2 _3401_ (.A(_1694_),
    .B(_1732_),
    .Y(_1783_));
 sky130_fd_sc_hd__nor2_2 _3402_ (.A(net368),
    .B(net165),
    .Y(_1784_));
 sky130_fd_sc_hd__or2_2 _3403_ (.A(net368),
    .B(net165),
    .X(_1785_));
 sky130_fd_sc_hd__o22a_1 _3404_ (.A1(net227),
    .A2(_1783_),
    .B1(_1785_),
    .B2(net1740),
    .X(_0317_));
 sky130_fd_sc_hd__o22a_1 _3405_ (.A1(net346),
    .A2(_1783_),
    .B1(_1785_),
    .B2(net512),
    .X(_0318_));
 sky130_fd_sc_hd__a22o_1 _3406_ (.A1(net269),
    .A2(net164),
    .B1(net100),
    .B2(net1806),
    .X(_0319_));
 sky130_fd_sc_hd__a22o_1 _3407_ (.A1(net262),
    .A2(net165),
    .B1(net101),
    .B2(net1228),
    .X(_0320_));
 sky130_fd_sc_hd__o22a_1 _3408_ (.A1(net259),
    .A2(_1783_),
    .B1(_1785_),
    .B2(net596),
    .X(_0321_));
 sky130_fd_sc_hd__o22a_1 _3409_ (.A1(net258),
    .A2(_1783_),
    .B1(_1785_),
    .B2(net696),
    .X(_0322_));
 sky130_fd_sc_hd__a22o_1 _3410_ (.A1(net256),
    .A2(net165),
    .B1(net101),
    .B2(net1730),
    .X(_0323_));
 sky130_fd_sc_hd__a22o_1 _3411_ (.A1(net254),
    .A2(net164),
    .B1(net100),
    .B2(net1734),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _3412_ (.A1(net252),
    .A2(net165),
    .B1(net100),
    .B2(net1190),
    .X(_0325_));
 sky130_fd_sc_hd__a22o_1 _3413_ (.A1(net250),
    .A2(net164),
    .B1(net100),
    .B2(net706),
    .X(_0326_));
 sky130_fd_sc_hd__a22o_1 _3414_ (.A1(net226),
    .A2(net165),
    .B1(net101),
    .B2(net1132),
    .X(_0327_));
 sky130_fd_sc_hd__a22o_1 _3415_ (.A1(net364),
    .A2(net164),
    .B1(net100),
    .B2(net2056),
    .X(_0328_));
 sky130_fd_sc_hd__a22o_1 _3416_ (.A1(net362),
    .A2(net165),
    .B1(net101),
    .B2(net1964),
    .X(_0329_));
 sky130_fd_sc_hd__a22o_1 _3417_ (.A1(net360),
    .A2(net164),
    .B1(net100),
    .B2(net1054),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _3418_ (.A1(net358),
    .A2(net165),
    .B1(net101),
    .B2(net1906),
    .X(_0331_));
 sky130_fd_sc_hd__a22o_1 _3419_ (.A1(net356),
    .A2(net164),
    .B1(net100),
    .B2(net1800),
    .X(_0332_));
 sky130_fd_sc_hd__a22o_1 _3420_ (.A1(net354),
    .A2(net165),
    .B1(net101),
    .B2(net1396),
    .X(_0333_));
 sky130_fd_sc_hd__a22o_1 _3421_ (.A1(net352),
    .A2(net165),
    .B1(net101),
    .B2(net1590),
    .X(_0334_));
 sky130_fd_sc_hd__a22o_1 _3422_ (.A1(net350),
    .A2(net164),
    .B1(net100),
    .B2(net1488),
    .X(_0335_));
 sky130_fd_sc_hd__a22o_1 _3423_ (.A1(net348),
    .A2(net165),
    .B1(net101),
    .B2(net1548),
    .X(_0336_));
 sky130_fd_sc_hd__a22o_1 _3424_ (.A1(net317),
    .A2(net165),
    .B1(net101),
    .B2(net1350),
    .X(_0337_));
 sky130_fd_sc_hd__a22o_1 _3425_ (.A1(net315),
    .A2(net164),
    .B1(net100),
    .B2(net1908),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _3426_ (.A1(net313),
    .A2(net164),
    .B1(net100),
    .B2(net2004),
    .X(_0339_));
 sky130_fd_sc_hd__a22o_1 _3427_ (.A1(net311),
    .A2(net164),
    .B1(net100),
    .B2(net890),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _3428_ (.A1(net309),
    .A2(net164),
    .B1(net100),
    .B2(net2192),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _3429_ (.A1(net307),
    .A2(net164),
    .B1(net100),
    .B2(net2082),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _3430_ (.A1(net303),
    .A2(net164),
    .B1(net101),
    .B2(net1696),
    .X(_0343_));
 sky130_fd_sc_hd__a22o_1 _3431_ (.A1(net302),
    .A2(net165),
    .B1(net101),
    .B2(net1038),
    .X(_0344_));
 sky130_fd_sc_hd__a22o_1 _3432_ (.A1(net300),
    .A2(net164),
    .B1(net100),
    .B2(net1980),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_1 _3433_ (.A1(net298),
    .A2(net164),
    .B1(net100),
    .B2(net1938),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _3434_ (.A1(net267),
    .A2(net164),
    .B1(net100),
    .B2(net1492),
    .X(_0347_));
 sky130_fd_sc_hd__a22o_1 _3435_ (.A1(net265),
    .A2(net165),
    .B1(net101),
    .B2(net716),
    .X(_0348_));
 sky130_fd_sc_hd__and3_1 _3436_ (.A(_1027_),
    .B(net217),
    .C(_1693_),
    .X(_1786_));
 sky130_fd_sc_hd__nand2_1 _3437_ (.A(_1027_),
    .B(_1694_),
    .Y(_1787_));
 sky130_fd_sc_hd__nor2_1 _3438_ (.A(net367),
    .B(net163),
    .Y(_1788_));
 sky130_fd_sc_hd__or2_1 _3439_ (.A(net366),
    .B(net163),
    .X(_1789_));
 sky130_fd_sc_hd__o22a_1 _3440_ (.A1(net228),
    .A2(_1787_),
    .B1(_1789_),
    .B2(net414),
    .X(_0349_));
 sky130_fd_sc_hd__o22a_1 _3441_ (.A1(net345),
    .A2(_1787_),
    .B1(_1789_),
    .B2(net376),
    .X(_0350_));
 sky130_fd_sc_hd__a22o_1 _3442_ (.A1(net268),
    .A2(net162),
    .B1(net98),
    .B2(net2052),
    .X(_0351_));
 sky130_fd_sc_hd__a22o_1 _3443_ (.A1(net263),
    .A2(net163),
    .B1(net99),
    .B2(net1242),
    .X(_0352_));
 sky130_fd_sc_hd__o22a_1 _3444_ (.A1(net260),
    .A2(_1787_),
    .B1(_1789_),
    .B2(net474),
    .X(_0353_));
 sky130_fd_sc_hd__o22a_1 _3445_ (.A1(net257),
    .A2(_1787_),
    .B1(_1789_),
    .B2(net568),
    .X(_0354_));
 sky130_fd_sc_hd__a22o_1 _3446_ (.A1(net255),
    .A2(net163),
    .B1(net99),
    .B2(net1848),
    .X(_0355_));
 sky130_fd_sc_hd__a22o_1 _3447_ (.A1(net253),
    .A2(net162),
    .B1(net98),
    .B2(net2206),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _3448_ (.A1(net251),
    .A2(net162),
    .B1(net98),
    .B2(net2250),
    .X(_0357_));
 sky130_fd_sc_hd__a22o_1 _3449_ (.A1(net249),
    .A2(net162),
    .B1(net98),
    .B2(net2168),
    .X(_0358_));
 sky130_fd_sc_hd__a22o_1 _3450_ (.A1(net225),
    .A2(net162),
    .B1(net98),
    .B2(net2288),
    .X(_0359_));
 sky130_fd_sc_hd__a22o_1 _3451_ (.A1(net363),
    .A2(net162),
    .B1(net98),
    .B2(net2202),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _3452_ (.A1(net361),
    .A2(net163),
    .B1(net99),
    .B2(net1048),
    .X(_0361_));
 sky130_fd_sc_hd__a22o_1 _3453_ (.A1(net359),
    .A2(net163),
    .B1(net98),
    .B2(net2096),
    .X(_0362_));
 sky130_fd_sc_hd__a22o_1 _3454_ (.A1(net357),
    .A2(net163),
    .B1(net99),
    .B2(net764),
    .X(_0363_));
 sky130_fd_sc_hd__a22o_1 _3455_ (.A1(net355),
    .A2(net162),
    .B1(net98),
    .B2(net1532),
    .X(_0364_));
 sky130_fd_sc_hd__a22o_1 _3456_ (.A1(net353),
    .A2(net163),
    .B1(net99),
    .B2(net1678),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _3457_ (.A1(net351),
    .A2(net163),
    .B1(net99),
    .B2(net1340),
    .X(_0366_));
 sky130_fd_sc_hd__a22o_1 _3458_ (.A1(net349),
    .A2(net162),
    .B1(net99),
    .B2(net1968),
    .X(_0367_));
 sky130_fd_sc_hd__a22o_1 _3459_ (.A1(net347),
    .A2(net163),
    .B1(net99),
    .B2(net904),
    .X(_0368_));
 sky130_fd_sc_hd__a22o_1 _3460_ (.A1(net316),
    .A2(net163),
    .B1(net99),
    .B2(net2118),
    .X(_0369_));
 sky130_fd_sc_hd__a22o_1 _3461_ (.A1(net314),
    .A2(net163),
    .B1(net99),
    .B2(net2018),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _3462_ (.A1(net312),
    .A2(net162),
    .B1(net98),
    .B2(net1708),
    .X(_0371_));
 sky130_fd_sc_hd__a22o_1 _3463_ (.A1(net310),
    .A2(net162),
    .B1(net98),
    .B2(net1344),
    .X(_0372_));
 sky130_fd_sc_hd__a22o_1 _3464_ (.A1(net308),
    .A2(net162),
    .B1(net98),
    .B2(net1896),
    .X(_0373_));
 sky130_fd_sc_hd__a22o_1 _3465_ (.A1(net306),
    .A2(net162),
    .B1(net98),
    .B2(net1946),
    .X(_0374_));
 sky130_fd_sc_hd__a22o_1 _3466_ (.A1(net305),
    .A2(net162),
    .B1(net98),
    .B2(net1366),
    .X(_0375_));
 sky130_fd_sc_hd__a22o_1 _3467_ (.A1(net301),
    .A2(net163),
    .B1(net99),
    .B2(net1348),
    .X(_0376_));
 sky130_fd_sc_hd__a22o_1 _3468_ (.A1(net299),
    .A2(net162),
    .B1(net98),
    .B2(net1584),
    .X(_0377_));
 sky130_fd_sc_hd__a22o_1 _3469_ (.A1(net297),
    .A2(net162),
    .B1(net98),
    .B2(net1698),
    .X(_0378_));
 sky130_fd_sc_hd__a22o_1 _3470_ (.A1(net266),
    .A2(net162),
    .B1(net98),
    .B2(net1466),
    .X(_0379_));
 sky130_fd_sc_hd__a22o_1 _3471_ (.A1(net265),
    .A2(net163),
    .B1(net99),
    .B2(net1804),
    .X(_0380_));
 sky130_fd_sc_hd__and3_1 _3472_ (.A(_1028_),
    .B(net217),
    .C(_1693_),
    .X(_1790_));
 sky130_fd_sc_hd__nand2_2 _3473_ (.A(_1028_),
    .B(_1694_),
    .Y(_1791_));
 sky130_fd_sc_hd__nor2_1 _3474_ (.A(net366),
    .B(net161),
    .Y(_1792_));
 sky130_fd_sc_hd__or2_2 _3475_ (.A(net366),
    .B(net161),
    .X(_1793_));
 sky130_fd_sc_hd__o22a_1 _3476_ (.A1(net228),
    .A2(_1791_),
    .B1(_1793_),
    .B2(net492),
    .X(_0381_));
 sky130_fd_sc_hd__o22a_1 _3477_ (.A1(net345),
    .A2(_1791_),
    .B1(_1793_),
    .B2(net456),
    .X(_0382_));
 sky130_fd_sc_hd__a22o_1 _3478_ (.A1(net268),
    .A2(net160),
    .B1(net96),
    .B2(net824),
    .X(_0383_));
 sky130_fd_sc_hd__a22o_1 _3479_ (.A1(net263),
    .A2(net161),
    .B1(net97),
    .B2(net1596),
    .X(_0384_));
 sky130_fd_sc_hd__o22a_1 _3480_ (.A1(net260),
    .A2(_1791_),
    .B1(_1793_),
    .B2(net520),
    .X(_0385_));
 sky130_fd_sc_hd__o22a_1 _3481_ (.A1(net257),
    .A2(_1791_),
    .B1(_1793_),
    .B2(net1266),
    .X(_0386_));
 sky130_fd_sc_hd__a22o_1 _3482_ (.A1(net255),
    .A2(net161),
    .B1(net97),
    .B2(net1052),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _3483_ (.A1(net253),
    .A2(net160),
    .B1(net96),
    .B2(net914),
    .X(_0388_));
 sky130_fd_sc_hd__a22o_1 _3484_ (.A1(net251),
    .A2(net160),
    .B1(net96),
    .B2(net2258),
    .X(_0389_));
 sky130_fd_sc_hd__a22o_1 _3485_ (.A1(net249),
    .A2(net160),
    .B1(net96),
    .B2(net2318),
    .X(_0390_));
 sky130_fd_sc_hd__a22o_1 _3486_ (.A1(net225),
    .A2(net161),
    .B1(net97),
    .B2(net1566),
    .X(_0391_));
 sky130_fd_sc_hd__a22o_1 _3487_ (.A1(net363),
    .A2(net160),
    .B1(net96),
    .B2(net1858),
    .X(_0392_));
 sky130_fd_sc_hd__a22o_1 _3488_ (.A1(net361),
    .A2(net161),
    .B1(net97),
    .B2(net1186),
    .X(_0393_));
 sky130_fd_sc_hd__a22o_1 _3489_ (.A1(net359),
    .A2(net160),
    .B1(net96),
    .B2(net2208),
    .X(_0394_));
 sky130_fd_sc_hd__a22o_1 _3490_ (.A1(net357),
    .A2(net161),
    .B1(net97),
    .B2(net1342),
    .X(_0395_));
 sky130_fd_sc_hd__a22o_1 _3491_ (.A1(net355),
    .A2(net160),
    .B1(net96),
    .B2(net948),
    .X(_0396_));
 sky130_fd_sc_hd__a22o_1 _3492_ (.A1(net353),
    .A2(net161),
    .B1(net97),
    .B2(net924),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _3493_ (.A1(net351),
    .A2(net161),
    .B1(net97),
    .B2(net1426),
    .X(_0398_));
 sky130_fd_sc_hd__a22o_1 _3494_ (.A1(net349),
    .A2(net160),
    .B1(net97),
    .B2(net2268),
    .X(_0399_));
 sky130_fd_sc_hd__a22o_1 _3495_ (.A1(net347),
    .A2(net161),
    .B1(net97),
    .B2(net886),
    .X(_0400_));
 sky130_fd_sc_hd__a22o_1 _3496_ (.A1(net316),
    .A2(net161),
    .B1(net97),
    .B2(net2016),
    .X(_0401_));
 sky130_fd_sc_hd__a22o_1 _3497_ (.A1(net314),
    .A2(net160),
    .B1(net96),
    .B2(net1432),
    .X(_0402_));
 sky130_fd_sc_hd__a22o_1 _3498_ (.A1(net312),
    .A2(net160),
    .B1(net96),
    .B2(net2024),
    .X(_0403_));
 sky130_fd_sc_hd__a22o_1 _3499_ (.A1(net310),
    .A2(net161),
    .B1(net96),
    .B2(net1868),
    .X(_0404_));
 sky130_fd_sc_hd__a22o_1 _3500_ (.A1(net308),
    .A2(net160),
    .B1(net96),
    .B2(net2322),
    .X(_0405_));
 sky130_fd_sc_hd__a22o_1 _3501_ (.A1(net306),
    .A2(net160),
    .B1(net96),
    .B2(net846),
    .X(_0406_));
 sky130_fd_sc_hd__a22o_1 _3502_ (.A1(net305),
    .A2(net160),
    .B1(net96),
    .B2(net954),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _3503_ (.A1(net301),
    .A2(net161),
    .B1(net97),
    .B2(net1948),
    .X(_0408_));
 sky130_fd_sc_hd__a22o_1 _3504_ (.A1(net299),
    .A2(net160),
    .B1(net96),
    .B2(net1162),
    .X(_0409_));
 sky130_fd_sc_hd__a22o_1 _3505_ (.A1(net297),
    .A2(net160),
    .B1(net96),
    .B2(net1308),
    .X(_0410_));
 sky130_fd_sc_hd__a22o_1 _3506_ (.A1(net266),
    .A2(net160),
    .B1(net96),
    .B2(net656),
    .X(_0411_));
 sky130_fd_sc_hd__a22o_1 _3507_ (.A1(net265),
    .A2(net161),
    .B1(net97),
    .B2(net658),
    .X(_0412_));
 sky130_fd_sc_hd__and3_1 _3508_ (.A(net216),
    .B(_1675_),
    .C(_1741_),
    .X(_1794_));
 sky130_fd_sc_hd__nand2_1 _3509_ (.A(_1676_),
    .B(_1741_),
    .Y(_1795_));
 sky130_fd_sc_hd__nor2_1 _3510_ (.A(net368),
    .B(net159),
    .Y(_1796_));
 sky130_fd_sc_hd__or2_2 _3511_ (.A(net366),
    .B(net159),
    .X(_1797_));
 sky130_fd_sc_hd__o22a_1 _3512_ (.A1(net227),
    .A2(_1795_),
    .B1(_1797_),
    .B2(net544),
    .X(_0413_));
 sky130_fd_sc_hd__o22a_1 _3513_ (.A1(net346),
    .A2(_1795_),
    .B1(_1797_),
    .B2(net438),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _3514_ (.A1(net269),
    .A2(net158),
    .B1(net94),
    .B2(net996),
    .X(_0415_));
 sky130_fd_sc_hd__a22o_1 _3515_ (.A1(net262),
    .A2(net159),
    .B1(net95),
    .B2(net864),
    .X(_0416_));
 sky130_fd_sc_hd__o22a_1 _3516_ (.A1(net259),
    .A2(_1795_),
    .B1(_1797_),
    .B2(net552),
    .X(_0417_));
 sky130_fd_sc_hd__o22a_1 _3517_ (.A1(net258),
    .A2(_1795_),
    .B1(_1797_),
    .B2(net518),
    .X(_0418_));
 sky130_fd_sc_hd__a22o_1 _3518_ (.A1(net256),
    .A2(net159),
    .B1(net95),
    .B2(net1562),
    .X(_0419_));
 sky130_fd_sc_hd__a22o_1 _3519_ (.A1(net254),
    .A2(net158),
    .B1(net94),
    .B2(net778),
    .X(_0420_));
 sky130_fd_sc_hd__a22o_1 _3520_ (.A1(net252),
    .A2(net158),
    .B1(net94),
    .B2(net1764),
    .X(_0421_));
 sky130_fd_sc_hd__a22o_1 _3521_ (.A1(net250),
    .A2(net158),
    .B1(net94),
    .B2(net1046),
    .X(_0422_));
 sky130_fd_sc_hd__a22o_1 _3522_ (.A1(net226),
    .A2(net159),
    .B1(net95),
    .B2(net1328),
    .X(_0423_));
 sky130_fd_sc_hd__a22o_1 _3523_ (.A1(net364),
    .A2(net158),
    .B1(net94),
    .B2(net2010),
    .X(_0424_));
 sky130_fd_sc_hd__a22o_1 _3524_ (.A1(net362),
    .A2(net159),
    .B1(net95),
    .B2(net1424),
    .X(_0425_));
 sky130_fd_sc_hd__a22o_1 _3525_ (.A1(net360),
    .A2(net158),
    .B1(net94),
    .B2(net1604),
    .X(_0426_));
 sky130_fd_sc_hd__a22o_1 _3526_ (.A1(net358),
    .A2(net159),
    .B1(net95),
    .B2(net976),
    .X(_0427_));
 sky130_fd_sc_hd__a22o_1 _3527_ (.A1(net356),
    .A2(net158),
    .B1(net94),
    .B2(net1378),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_1 _3528_ (.A1(net354),
    .A2(net159),
    .B1(net95),
    .B2(net720),
    .X(_0429_));
 sky130_fd_sc_hd__a22o_1 _3529_ (.A1(net352),
    .A2(net159),
    .B1(net95),
    .B2(net1104),
    .X(_0430_));
 sky130_fd_sc_hd__a22o_1 _3530_ (.A1(net350),
    .A2(net158),
    .B1(net94),
    .B2(net1288),
    .X(_0431_));
 sky130_fd_sc_hd__a22o_1 _3531_ (.A1(net348),
    .A2(net159),
    .B1(net95),
    .B2(net1170),
    .X(_0432_));
 sky130_fd_sc_hd__a22o_1 _3532_ (.A1(net317),
    .A2(net159),
    .B1(net95),
    .B2(net1704),
    .X(_0433_));
 sky130_fd_sc_hd__a22o_1 _3533_ (.A1(net315),
    .A2(net158),
    .B1(net94),
    .B2(net1084),
    .X(_0434_));
 sky130_fd_sc_hd__a22o_1 _3534_ (.A1(net313),
    .A2(net158),
    .B1(net94),
    .B2(net1668),
    .X(_0435_));
 sky130_fd_sc_hd__a22o_1 _3535_ (.A1(net311),
    .A2(net158),
    .B1(net94),
    .B2(net1790),
    .X(_0436_));
 sky130_fd_sc_hd__a22o_1 _3536_ (.A1(net309),
    .A2(net158),
    .B1(net94),
    .B2(net1338),
    .X(_0437_));
 sky130_fd_sc_hd__a22o_1 _3537_ (.A1(net307),
    .A2(net159),
    .B1(net95),
    .B2(net2140),
    .X(_0438_));
 sky130_fd_sc_hd__a22o_1 _3538_ (.A1(net303),
    .A2(net158),
    .B1(net94),
    .B2(net1144),
    .X(_0439_));
 sky130_fd_sc_hd__a22o_1 _3539_ (.A1(net302),
    .A2(net159),
    .B1(net95),
    .B2(net944),
    .X(_0440_));
 sky130_fd_sc_hd__a22o_1 _3540_ (.A1(net300),
    .A2(net158),
    .B1(net94),
    .B2(net668),
    .X(_0441_));
 sky130_fd_sc_hd__a22o_1 _3541_ (.A1(net298),
    .A2(net158),
    .B1(net94),
    .B2(net1060),
    .X(_0442_));
 sky130_fd_sc_hd__a22o_1 _3542_ (.A1(net267),
    .A2(net158),
    .B1(net94),
    .B2(net1082),
    .X(_0443_));
 sky130_fd_sc_hd__a22o_1 _3543_ (.A1(net265),
    .A2(net159),
    .B1(net95),
    .B2(net1230),
    .X(_0444_));
 sky130_fd_sc_hd__and3_1 _3544_ (.A(net216),
    .B(_1675_),
    .C(_1686_),
    .X(_1798_));
 sky130_fd_sc_hd__nand2_1 _3545_ (.A(_1676_),
    .B(_1686_),
    .Y(_1799_));
 sky130_fd_sc_hd__nor2_1 _3546_ (.A(net369),
    .B(net156),
    .Y(_1800_));
 sky130_fd_sc_hd__or2_2 _3547_ (.A(net366),
    .B(net156),
    .X(_1801_));
 sky130_fd_sc_hd__o22a_1 _3548_ (.A1(net227),
    .A2(_1799_),
    .B1(_1801_),
    .B2(net546),
    .X(_0445_));
 sky130_fd_sc_hd__o22a_1 _3549_ (.A1(net346),
    .A2(_1799_),
    .B1(_1801_),
    .B2(net472),
    .X(_0446_));
 sky130_fd_sc_hd__a22o_1 _3550_ (.A1(net269),
    .A2(net157),
    .B1(net92),
    .B2(net1928),
    .X(_0447_));
 sky130_fd_sc_hd__a22o_1 _3551_ (.A1(net262),
    .A2(net156),
    .B1(net93),
    .B2(net832),
    .X(_0448_));
 sky130_fd_sc_hd__o22a_1 _3552_ (.A1(net259),
    .A2(_1799_),
    .B1(_1801_),
    .B2(net488),
    .X(_0449_));
 sky130_fd_sc_hd__o22a_1 _3553_ (.A1(net258),
    .A2(_1799_),
    .B1(_1801_),
    .B2(net440),
    .X(_0450_));
 sky130_fd_sc_hd__a22o_1 _3554_ (.A1(net256),
    .A2(net156),
    .B1(net93),
    .B2(net1634),
    .X(_0451_));
 sky130_fd_sc_hd__a22o_1 _3555_ (.A1(net254),
    .A2(net157),
    .B1(net92),
    .B2(net2260),
    .X(_0452_));
 sky130_fd_sc_hd__a22o_1 _3556_ (.A1(net252),
    .A2(net156),
    .B1(net92),
    .B2(net1200),
    .X(_0453_));
 sky130_fd_sc_hd__a22o_1 _3557_ (.A1(net250),
    .A2(net157),
    .B1(net92),
    .B2(net1776),
    .X(_0454_));
 sky130_fd_sc_hd__a22o_1 _3558_ (.A1(net226),
    .A2(net156),
    .B1(net93),
    .B2(net1086),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _3559_ (.A1(net364),
    .A2(net157),
    .B1(net92),
    .B2(net1782),
    .X(_0456_));
 sky130_fd_sc_hd__a22o_1 _3560_ (.A1(net362),
    .A2(net156),
    .B1(net93),
    .B2(net1202),
    .X(_0457_));
 sky130_fd_sc_hd__a22o_1 _3561_ (.A1(net360),
    .A2(net157),
    .B1(net92),
    .B2(net1108),
    .X(_0458_));
 sky130_fd_sc_hd__a22o_1 _3562_ (.A1(net358),
    .A2(net156),
    .B1(net93),
    .B2(net1528),
    .X(_0459_));
 sky130_fd_sc_hd__a22o_1 _3563_ (.A1(net356),
    .A2(net156),
    .B1(net93),
    .B2(net702),
    .X(_0460_));
 sky130_fd_sc_hd__a22o_1 _3564_ (.A1(net354),
    .A2(net156),
    .B1(net93),
    .B2(net994),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _3565_ (.A1(net352),
    .A2(net156),
    .B1(net93),
    .B2(net1252),
    .X(_0462_));
 sky130_fd_sc_hd__a22o_1 _3566_ (.A1(net350),
    .A2(net157),
    .B1(net92),
    .B2(net964),
    .X(_0463_));
 sky130_fd_sc_hd__a22o_1 _3567_ (.A1(net348),
    .A2(net157),
    .B1(net93),
    .B2(net620),
    .X(_0464_));
 sky130_fd_sc_hd__a22o_1 _3568_ (.A1(net317),
    .A2(net156),
    .B1(net93),
    .B2(net1516),
    .X(_0465_));
 sky130_fd_sc_hd__a22o_1 _3569_ (.A1(net315),
    .A2(net156),
    .B1(net92),
    .B2(net1714),
    .X(_0466_));
 sky130_fd_sc_hd__a22o_1 _3570_ (.A1(net313),
    .A2(net157),
    .B1(net92),
    .B2(net1496),
    .X(_0467_));
 sky130_fd_sc_hd__a22o_1 _3571_ (.A1(net311),
    .A2(net157),
    .B1(net92),
    .B2(net1574),
    .X(_0468_));
 sky130_fd_sc_hd__a22o_1 _3572_ (.A1(net309),
    .A2(net157),
    .B1(net92),
    .B2(net1918),
    .X(_0469_));
 sky130_fd_sc_hd__a22o_1 _3573_ (.A1(net307),
    .A2(net157),
    .B1(net92),
    .B2(net2102),
    .X(_0470_));
 sky130_fd_sc_hd__a22o_1 _3574_ (.A1(net303),
    .A2(net156),
    .B1(net92),
    .B2(net724),
    .X(_0471_));
 sky130_fd_sc_hd__a22o_1 _3575_ (.A1(net302),
    .A2(net156),
    .B1(net93),
    .B2(net1022),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _3576_ (.A1(net300),
    .A2(net157),
    .B1(net92),
    .B2(net628),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _3577_ (.A1(net298),
    .A2(net157),
    .B1(net92),
    .B2(net812),
    .X(_0474_));
 sky130_fd_sc_hd__a22o_1 _3578_ (.A1(net267),
    .A2(net157),
    .B1(net92),
    .B2(net704),
    .X(_0475_));
 sky130_fd_sc_hd__a22o_1 _3579_ (.A1(net265),
    .A2(net156),
    .B1(net93),
    .B2(net1842),
    .X(_0476_));
 sky130_fd_sc_hd__and4b_1 _3580_ (.A_N(net291),
    .B(net339),
    .C(_1669_),
    .D(_1686_),
    .X(_1802_));
 sky130_fd_sc_hd__nand2_1 _3581_ (.A(_1670_),
    .B(_1686_),
    .Y(_1803_));
 sky130_fd_sc_hd__nor2_1 _3582_ (.A(net368),
    .B(net154),
    .Y(_1804_));
 sky130_fd_sc_hd__or2_2 _3583_ (.A(net367),
    .B(net154),
    .X(_1805_));
 sky130_fd_sc_hd__o22a_1 _3584_ (.A1(net8),
    .A2(_1803_),
    .B1(_1805_),
    .B2(net428),
    .X(_0477_));
 sky130_fd_sc_hd__o22a_1 _3585_ (.A1(net346),
    .A2(_1803_),
    .B1(_1805_),
    .B2(net398),
    .X(_0478_));
 sky130_fd_sc_hd__a22o_1 _3586_ (.A1(net269),
    .A2(net155),
    .B1(net90),
    .B2(net1074),
    .X(_0479_));
 sky130_fd_sc_hd__a22o_1 _3587_ (.A1(net262),
    .A2(net154),
    .B1(net90),
    .B2(net796),
    .X(_0480_));
 sky130_fd_sc_hd__o22a_1 _3588_ (.A1(net259),
    .A2(_1803_),
    .B1(_1805_),
    .B2(net418),
    .X(_0481_));
 sky130_fd_sc_hd__o22a_1 _3589_ (.A1(net258),
    .A2(_1803_),
    .B1(_1805_),
    .B2(net392),
    .X(_0482_));
 sky130_fd_sc_hd__a22o_1 _3590_ (.A1(net256),
    .A2(net154),
    .B1(net91),
    .B2(net1670),
    .X(_0483_));
 sky130_fd_sc_hd__a22o_1 _3591_ (.A1(net254),
    .A2(net155),
    .B1(net90),
    .B2(net1784),
    .X(_0484_));
 sky130_fd_sc_hd__a22o_1 _3592_ (.A1(net252),
    .A2(net154),
    .B1(net91),
    .B2(net1044),
    .X(_0485_));
 sky130_fd_sc_hd__a22o_1 _3593_ (.A1(net250),
    .A2(net155),
    .B1(net90),
    .B2(net1592),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_1 _3594_ (.A1(net226),
    .A2(net154),
    .B1(net91),
    .B2(net762),
    .X(_0487_));
 sky130_fd_sc_hd__a22o_1 _3595_ (.A1(net364),
    .A2(net155),
    .B1(net90),
    .B2(net1244),
    .X(_0488_));
 sky130_fd_sc_hd__a22o_1 _3596_ (.A1(net362),
    .A2(net154),
    .B1(net91),
    .B2(net688),
    .X(_0489_));
 sky130_fd_sc_hd__a22o_1 _3597_ (.A1(net360),
    .A2(net155),
    .B1(net90),
    .B2(net838),
    .X(_0490_));
 sky130_fd_sc_hd__a22o_1 _3598_ (.A1(net358),
    .A2(net154),
    .B1(net91),
    .B2(net1398),
    .X(_0491_));
 sky130_fd_sc_hd__a22o_1 _3599_ (.A1(net356),
    .A2(net154),
    .B1(net91),
    .B2(net774),
    .X(_0492_));
 sky130_fd_sc_hd__a22o_1 _3600_ (.A1(net354),
    .A2(net155),
    .B1(net91),
    .B2(net1062),
    .X(_0493_));
 sky130_fd_sc_hd__a22o_1 _3601_ (.A1(net352),
    .A2(net154),
    .B1(net91),
    .B2(net814),
    .X(_0494_));
 sky130_fd_sc_hd__a22o_1 _3602_ (.A1(net350),
    .A2(net155),
    .B1(net90),
    .B2(net1112),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _3603_ (.A1(net348),
    .A2(net154),
    .B1(net91),
    .B2(net1126),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _3604_ (.A1(net317),
    .A2(net154),
    .B1(net91),
    .B2(net1628),
    .X(_0497_));
 sky130_fd_sc_hd__a22o_1 _3605_ (.A1(net315),
    .A2(net154),
    .B1(net90),
    .B2(net1254),
    .X(_0498_));
 sky130_fd_sc_hd__a22o_1 _3606_ (.A1(net313),
    .A2(net155),
    .B1(net90),
    .B2(net1124),
    .X(_0499_));
 sky130_fd_sc_hd__a22o_1 _3607_ (.A1(net311),
    .A2(net155),
    .B1(net90),
    .B2(net962),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _3608_ (.A1(net309),
    .A2(net155),
    .B1(net90),
    .B2(net2020),
    .X(_0501_));
 sky130_fd_sc_hd__a22o_1 _3609_ (.A1(net307),
    .A2(net155),
    .B1(net90),
    .B2(net1892),
    .X(_0502_));
 sky130_fd_sc_hd__a22o_1 _3610_ (.A1(net304),
    .A2(net154),
    .B1(net90),
    .B2(net1300),
    .X(_0503_));
 sky130_fd_sc_hd__a22o_1 _3611_ (.A1(net302),
    .A2(net154),
    .B1(net91),
    .B2(net980),
    .X(_0504_));
 sky130_fd_sc_hd__a22o_1 _3612_ (.A1(net300),
    .A2(net155),
    .B1(net90),
    .B2(net930),
    .X(_0505_));
 sky130_fd_sc_hd__a22o_1 _3613_ (.A1(net298),
    .A2(net155),
    .B1(net90),
    .B2(net790),
    .X(_0506_));
 sky130_fd_sc_hd__a22o_1 _3614_ (.A1(net267),
    .A2(net155),
    .B1(net90),
    .B2(net1760),
    .X(_0507_));
 sky130_fd_sc_hd__a22o_1 _3615_ (.A1(net265),
    .A2(net154),
    .B1(net91),
    .B2(net862),
    .X(_0508_));
 sky130_fd_sc_hd__and4b_2 _3616_ (.A_N(net293),
    .B(net341),
    .C(_1669_),
    .D(_1732_),
    .X(_1806_));
 sky130_fd_sc_hd__nand2_2 _3617_ (.A(_1670_),
    .B(_1732_),
    .Y(_1807_));
 sky130_fd_sc_hd__nor2_1 _3618_ (.A(net369),
    .B(net153),
    .Y(_1808_));
 sky130_fd_sc_hd__or2_2 _3619_ (.A(net368),
    .B(net153),
    .X(_1809_));
 sky130_fd_sc_hd__o22a_1 _3620_ (.A1(net228),
    .A2(_1807_),
    .B1(_1809_),
    .B2(net538),
    .X(_0509_));
 sky130_fd_sc_hd__o22a_1 _3621_ (.A1(net346),
    .A2(_1807_),
    .B1(_1809_),
    .B2(net570),
    .X(_0510_));
 sky130_fd_sc_hd__a22o_1 _3622_ (.A1(net269),
    .A2(net152),
    .B1(net88),
    .B2(net1818),
    .X(_0511_));
 sky130_fd_sc_hd__a22o_1 _3623_ (.A1(net262),
    .A2(net153),
    .B1(net89),
    .B2(net1092),
    .X(_0512_));
 sky130_fd_sc_hd__o22a_1 _3624_ (.A1(net34),
    .A2(_1807_),
    .B1(_1809_),
    .B2(net548),
    .X(_0513_));
 sky130_fd_sc_hd__o22a_1 _3625_ (.A1(net258),
    .A2(_1807_),
    .B1(_1809_),
    .B2(net600),
    .X(_0514_));
 sky130_fd_sc_hd__a22o_1 _3626_ (.A1(net256),
    .A2(net153),
    .B1(net88),
    .B2(net1184),
    .X(_0515_));
 sky130_fd_sc_hd__a22o_1 _3627_ (.A1(net254),
    .A2(net152),
    .B1(net88),
    .B2(net2104),
    .X(_0516_));
 sky130_fd_sc_hd__a22o_1 _3628_ (.A1(net252),
    .A2(net153),
    .B1(net88),
    .B2(net1334),
    .X(_0517_));
 sky130_fd_sc_hd__a22o_1 _3629_ (.A1(net250),
    .A2(net152),
    .B1(net88),
    .B2(net870),
    .X(_0518_));
 sky130_fd_sc_hd__a22o_1 _3630_ (.A1(net226),
    .A2(net153),
    .B1(net89),
    .B2(net1480),
    .X(_0519_));
 sky130_fd_sc_hd__a22o_1 _3631_ (.A1(net364),
    .A2(net152),
    .B1(net88),
    .B2(net2222),
    .X(_0520_));
 sky130_fd_sc_hd__a22o_1 _3632_ (.A1(net362),
    .A2(net153),
    .B1(net89),
    .B2(net840),
    .X(_0521_));
 sky130_fd_sc_hd__a22o_1 _3633_ (.A1(net360),
    .A2(net152),
    .B1(net88),
    .B2(net1420),
    .X(_0522_));
 sky130_fd_sc_hd__a22o_1 _3634_ (.A1(net358),
    .A2(net153),
    .B1(net89),
    .B2(net1510),
    .X(_0523_));
 sky130_fd_sc_hd__a22o_1 _3635_ (.A1(net356),
    .A2(net152),
    .B1(net89),
    .B2(net2124),
    .X(_0524_));
 sky130_fd_sc_hd__a22o_1 _3636_ (.A1(net354),
    .A2(net153),
    .B1(net89),
    .B2(net742),
    .X(_0525_));
 sky130_fd_sc_hd__a22o_1 _3637_ (.A1(net352),
    .A2(net153),
    .B1(net89),
    .B2(net1208),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _3638_ (.A1(net350),
    .A2(net152),
    .B1(net88),
    .B2(net1402),
    .X(_0527_));
 sky130_fd_sc_hd__a22o_1 _3639_ (.A1(net348),
    .A2(net153),
    .B1(net89),
    .B2(net1280),
    .X(_0528_));
 sky130_fd_sc_hd__a22o_1 _3640_ (.A1(net317),
    .A2(net153),
    .B1(net89),
    .B2(net1412),
    .X(_0529_));
 sky130_fd_sc_hd__a22o_1 _3641_ (.A1(net315),
    .A2(net152),
    .B1(net88),
    .B2(net1754),
    .X(_0530_));
 sky130_fd_sc_hd__a22o_1 _3642_ (.A1(net313),
    .A2(net152),
    .B1(net88),
    .B2(net730),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_1 _3643_ (.A1(net311),
    .A2(net152),
    .B1(net88),
    .B2(net506),
    .X(_0532_));
 sky130_fd_sc_hd__a22o_1 _3644_ (.A1(net309),
    .A2(net152),
    .B1(net88),
    .B2(net2410),
    .X(_0533_));
 sky130_fd_sc_hd__a22o_1 _3645_ (.A1(net307),
    .A2(net152),
    .B1(net88),
    .B2(net1728),
    .X(_0534_));
 sky130_fd_sc_hd__a22o_1 _3646_ (.A1(net304),
    .A2(net152),
    .B1(net89),
    .B2(net1836),
    .X(_0535_));
 sky130_fd_sc_hd__a22o_1 _3647_ (.A1(net302),
    .A2(net153),
    .B1(net89),
    .B2(net2228),
    .X(_0536_));
 sky130_fd_sc_hd__a22o_1 _3648_ (.A1(net300),
    .A2(net152),
    .B1(net88),
    .B2(net594),
    .X(_0537_));
 sky130_fd_sc_hd__a22o_1 _3649_ (.A1(net298),
    .A2(net152),
    .B1(net88),
    .B2(net810),
    .X(_0538_));
 sky130_fd_sc_hd__a22o_1 _3650_ (.A1(net267),
    .A2(net152),
    .B1(net88),
    .B2(net854),
    .X(_0539_));
 sky130_fd_sc_hd__a22o_1 _3651_ (.A1(net265),
    .A2(net153),
    .B1(net89),
    .B2(net2362),
    .X(_0540_));
 sky130_fd_sc_hd__dfxtp_1 _3652_ (.CLK(clknet_leaf_22_clk),
    .D(net477),
    .Q(\mem[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3653_ (.CLK(clknet_leaf_23_clk),
    .D(net389),
    .Q(\mem[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3654_ (.CLK(clknet_leaf_93_clk),
    .D(net619),
    .Q(\mem[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3655_ (.CLK(clknet_leaf_17_clk),
    .D(net875),
    .Q(\mem[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3656_ (.CLK(clknet_leaf_24_clk),
    .D(net449),
    .Q(\mem[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3657_ (.CLK(clknet_leaf_24_clk),
    .D(net529),
    .Q(\mem[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3658_ (.CLK(clknet_leaf_19_clk),
    .D(net1429),
    .Q(\mem[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3659_ (.CLK(clknet_leaf_3_clk),
    .D(net1331),
    .Q(\mem[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3660_ (.CLK(clknet_leaf_9_clk),
    .D(net2395),
    .Q(\mem[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3661_ (.CLK(clknet_leaf_90_clk),
    .D(net1285),
    .Q(\mem[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3662_ (.CLK(clknet_leaf_15_clk),
    .D(net615),
    .Q(\mem[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3663_ (.CLK(clknet_leaf_83_clk),
    .D(net1639),
    .Q(\mem[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3664_ (.CLK(clknet_leaf_17_clk),
    .D(net1661),
    .Q(\mem[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3665_ (.CLK(clknet_leaf_9_clk),
    .D(net2397),
    .Q(\mem[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3666_ (.CLK(clknet_leaf_18_clk),
    .D(net1451),
    .Q(\mem[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3667_ (.CLK(clknet_leaf_4_clk),
    .D(net2087),
    .Q(\mem[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3668_ (.CLK(clknet_leaf_18_clk),
    .D(net2221),
    .Q(\mem[21][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3669_ (.CLK(clknet_leaf_30_clk),
    .D(net767),
    .Q(\mem[21][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3670_ (.CLK(clknet_leaf_9_clk),
    .D(net1867),
    .Q(\mem[21][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3671_ (.CLK(clknet_leaf_11_clk),
    .D(net1665),
    .Q(\mem[21][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3672_ (.CLK(clknet_leaf_20_clk),
    .D(net2327),
    .Q(\mem[21][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3673_ (.CLK(clknet_leaf_7_clk),
    .D(net939),
    .Q(\mem[21][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3674_ (.CLK(clknet_leaf_84_clk),
    .D(net2007),
    .Q(\mem[21][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3675_ (.CLK(clknet_leaf_83_clk),
    .D(net985),
    .Q(\mem[21][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3676_ (.CLK(clknet_leaf_0_clk),
    .D(net2117),
    .Q(\mem[21][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3677_ (.CLK(clknet_leaf_83_clk),
    .D(net1559),
    .Q(\mem[21][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3678_ (.CLK(clknet_leaf_3_clk),
    .D(net859),
    .Q(\mem[21][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3679_ (.CLK(clknet_leaf_19_clk),
    .D(net679),
    .Q(\mem[21][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3680_ (.CLK(clknet_leaf_4_clk),
    .D(net913),
    .Q(\mem[21][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3681_ (.CLK(clknet_leaf_1_clk),
    .D(net843),
    .Q(\mem[21][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3682_ (.CLK(clknet_leaf_3_clk),
    .D(net1503),
    .Q(\mem[21][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3683_ (.CLK(clknet_leaf_15_clk),
    .D(net1073),
    .Q(\mem[21][31] ));
 sky130_fd_sc_hd__dfxtp_2 _3684_ (.CLK(clknet_leaf_59_clk),
    .D(_0573_),
    .Q(net42));
 sky130_fd_sc_hd__dfxtp_1 _3685_ (.CLK(clknet_leaf_22_clk),
    .D(net567),
    .Q(\mem[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3686_ (.CLK(clknet_leaf_23_clk),
    .D(net443),
    .Q(\mem[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3687_ (.CLK(clknet_leaf_93_clk),
    .D(net857),
    .Q(\mem[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3688_ (.CLK(clknet_leaf_17_clk),
    .D(net1875),
    .Q(\mem[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3689_ (.CLK(clknet_leaf_24_clk),
    .D(net587),
    .Q(\mem[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3690_ (.CLK(clknet_leaf_24_clk),
    .D(net897),
    .Q(\mem[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3691_ (.CLK(clknet_leaf_21_clk),
    .D(net853),
    .Q(\mem[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3692_ (.CLK(clknet_leaf_3_clk),
    .D(net1461),
    .Q(\mem[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3693_ (.CLK(clknet_leaf_9_clk),
    .D(net2305),
    .Q(\mem[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3694_ (.CLK(clknet_leaf_90_clk),
    .D(net1627),
    .Q(\mem[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3695_ (.CLK(clknet_leaf_16_clk),
    .D(net1181),
    .Q(\mem[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3696_ (.CLK(clknet_leaf_8_clk),
    .D(net1135),
    .Q(\mem[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3697_ (.CLK(clknet_leaf_17_clk),
    .D(net1743),
    .Q(\mem[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3698_ (.CLK(clknet_leaf_9_clk),
    .D(net2181),
    .Q(\mem[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3699_ (.CLK(clknet_leaf_18_clk),
    .D(net1931),
    .Q(\mem[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3700_ (.CLK(clknet_leaf_4_clk),
    .D(net1603),
    .Q(\mem[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3701_ (.CLK(clknet_leaf_17_clk),
    .D(net1257),
    .Q(\mem[22][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3702_ (.CLK(clknet_leaf_30_clk),
    .D(net1499),
    .Q(\mem[22][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3703_ (.CLK(clknet_leaf_8_clk),
    .D(net1599),
    .Q(\mem[22][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3704_ (.CLK(clknet_leaf_11_clk),
    .D(net2095),
    .Q(\mem[22][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3705_ (.CLK(clknet_leaf_20_clk),
    .D(net1955),
    .Q(\mem[22][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3706_ (.CLK(clknet_leaf_1_clk),
    .D(net2249),
    .Q(\mem[22][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3707_ (.CLK(clknet_leaf_84_clk),
    .D(net1747),
    .Q(\mem[22][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3708_ (.CLK(clknet_leaf_83_clk),
    .D(net1223),
    .Q(\mem[22][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3709_ (.CLK(clknet_leaf_93_clk),
    .D(net647),
    .Q(\mem[22][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3710_ (.CLK(clknet_leaf_83_clk),
    .D(net2111),
    .Q(\mem[22][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3711_ (.CLK(clknet_leaf_3_clk),
    .D(net1803),
    .Q(\mem[22][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3712_ (.CLK(clknet_leaf_18_clk),
    .D(net1525),
    .Q(\mem[22][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3713_ (.CLK(clknet_leaf_4_clk),
    .D(net2199),
    .Q(\mem[22][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3714_ (.CLK(clknet_leaf_1_clk),
    .D(net1873),
    .Q(\mem[22][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3715_ (.CLK(clknet_leaf_3_clk),
    .D(net901),
    .Q(\mem[22][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3716_ (.CLK(clknet_leaf_16_clk),
    .D(net1583),
    .Q(\mem[22][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3717_ (.CLK(clknet_leaf_28_clk),
    .D(net445),
    .Q(\mem[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3718_ (.CLK(clknet_leaf_28_clk),
    .D(net453),
    .Q(\mem[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3719_ (.CLK(clknet_leaf_90_clk),
    .D(net709),
    .Q(\mem[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3720_ (.CLK(clknet_leaf_10_clk),
    .D(net2079),
    .Q(\mem[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3721_ (.CLK(clknet_leaf_28_clk),
    .D(net417),
    .Q(\mem[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3722_ (.CLK(clknet_leaf_27_clk),
    .D(net469),
    .Q(\mem[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3723_ (.CLK(clknet_leaf_30_clk),
    .D(net733),
    .Q(\mem[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3724_ (.CLK(clknet_leaf_1_clk),
    .D(net1333),
    .Q(\mem[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3725_ (.CLK(clknet_leaf_10_clk),
    .D(net2353),
    .Q(\mem[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3726_ (.CLK(clknet_leaf_89_clk),
    .D(net1653),
    .Q(\mem[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3727_ (.CLK(clknet_leaf_6_clk),
    .D(net1297),
    .Q(\mem[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3728_ (.CLK(clknet_leaf_86_clk),
    .D(net1455),
    .Q(\mem[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3729_ (.CLK(clknet_leaf_11_clk),
    .D(net2139),
    .Q(\mem[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3730_ (.CLK(clknet_leaf_81_clk),
    .D(net1971),
    .Q(\mem[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3731_ (.CLK(clknet_leaf_12_clk),
    .D(net1303),
    .Q(\mem[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3732_ (.CLK(clknet_leaf_9_clk),
    .D(net2279),
    .Q(\mem[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3733_ (.CLK(clknet_leaf_14_clk),
    .D(net1797),
    .Q(\mem[30][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3734_ (.CLK(clknet_leaf_32_clk),
    .D(net1021),
    .Q(\mem[30][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3735_ (.CLK(clknet_leaf_82_clk),
    .D(net1691),
    .Q(\mem[30][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3736_ (.CLK(clknet_leaf_32_clk),
    .D(net1043),
    .Q(\mem[30][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3737_ (.CLK(clknet_leaf_22_clk),
    .D(net1377),
    .Q(\mem[30][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3738_ (.CLK(clknet_leaf_8_clk),
    .D(net1449),
    .Q(\mem[30][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3739_ (.CLK(clknet_leaf_82_clk),
    .D(net1773),
    .Q(\mem[30][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3740_ (.CLK(clknet_leaf_86_clk),
    .D(net681),
    .Q(\mem[30][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3741_ (.CLK(clknet_leaf_86_clk),
    .D(net2001),
    .Q(\mem[30][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3742_ (.CLK(clknet_leaf_85_clk),
    .D(net1129),
    .Q(\mem[30][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3743_ (.CLK(clknet_leaf_85_clk),
    .D(net753),
    .Q(\mem[30][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3744_ (.CLK(clknet_leaf_12_clk),
    .D(net1683),
    .Q(\mem[30][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3745_ (.CLK(clknet_leaf_7_clk),
    .D(net2061),
    .Q(\mem[30][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3746_ (.CLK(clknet_leaf_91_clk),
    .D(net969),
    .Q(\mem[30][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3747_ (.CLK(clknet_leaf_90_clk),
    .D(net1561),
    .Q(\mem[30][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3748_ (.CLK(clknet_leaf_33_clk),
    .D(net611),
    .Q(\mem[30][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3749_ (.CLK(clknet_leaf_42_clk),
    .D(net481),
    .Q(\mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3750_ (.CLK(clknet_leaf_41_clk),
    .D(net421),
    .Q(\mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3751_ (.CLK(clknet_leaf_73_clk),
    .D(net1179),
    .Q(\mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3752_ (.CLK(clknet_leaf_55_clk),
    .D(net1363),
    .Q(\mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3753_ (.CLK(clknet_leaf_41_clk),
    .D(net423),
    .Q(\mem[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3754_ (.CLK(clknet_leaf_42_clk),
    .D(net627),
    .Q(\mem[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3755_ (.CLK(clknet_leaf_51_clk),
    .D(net1353),
    .Q(\mem[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3756_ (.CLK(clknet_leaf_71_clk),
    .D(net1647),
    .Q(\mem[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3757_ (.CLK(clknet_leaf_57_clk),
    .D(net1141),
    .Q(\mem[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3758_ (.CLK(clknet_leaf_70_clk),
    .D(net1655),
    .Q(\mem[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3759_ (.CLK(clknet_leaf_50_clk),
    .D(net1235),
    .Q(\mem[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3760_ (.CLK(clknet_leaf_72_clk),
    .D(net2325),
    .Q(\mem[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3761_ (.CLK(clknet_leaf_36_clk),
    .D(net1119),
    .Q(\mem[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3762_ (.CLK(clknet_leaf_60_clk),
    .D(net745),
    .Q(\mem[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3763_ (.CLK(clknet_leaf_51_clk),
    .D(net2255),
    .Q(\mem[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3764_ (.CLK(clknet_leaf_61_clk),
    .D(net2023),
    .Q(\mem[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3765_ (.CLK(clknet_leaf_34_clk),
    .D(net1619),
    .Q(\mem[15][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3766_ (.CLK(clknet_leaf_46_clk),
    .D(net919),
    .Q(\mem[15][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3767_ (.CLK(clknet_leaf_58_clk),
    .D(net2137),
    .Q(\mem[15][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3768_ (.CLK(clknet_leaf_50_clk),
    .D(net1311),
    .Q(\mem[15][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3769_ (.CLK(clknet_leaf_38_clk),
    .D(net851),
    .Q(\mem[15][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3770_ (.CLK(clknet_leaf_60_clk),
    .D(net1273),
    .Q(\mem[15][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3771_ (.CLK(clknet_leaf_70_clk),
    .D(net2287),
    .Q(\mem[15][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3772_ (.CLK(clknet_leaf_69_clk),
    .D(net829),
    .Q(\mem[15][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3773_ (.CLK(clknet_leaf_72_clk),
    .D(net1411),
    .Q(\mem[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3774_ (.CLK(clknet_leaf_72_clk),
    .D(net1279),
    .Q(\mem[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3775_ (.CLK(clknet_leaf_56_clk),
    .D(net1325),
    .Q(\mem[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3776_ (.CLK(clknet_leaf_37_clk),
    .D(net631),
    .Q(\mem[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3777_ (.CLK(clknet_leaf_78_clk),
    .D(net1293),
    .Q(\mem[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3778_ (.CLK(clknet_leaf_72_clk),
    .D(net1519),
    .Q(\mem[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3779_ (.CLK(clknet_leaf_73_clk),
    .D(net993),
    .Q(\mem[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3780_ (.CLK(clknet_leaf_53_clk),
    .D(net1001),
    .Q(\mem[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3781_ (.CLK(clknet_leaf_26_clk),
    .D(net543),
    .Q(\mem[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3782_ (.CLK(clknet_leaf_26_clk),
    .D(net497),
    .Q(\mem[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3783_ (.CLK(clknet_leaf_92_clk),
    .D(net1569),
    .Q(\mem[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3784_ (.CLK(clknet_leaf_10_clk),
    .D(net2205),
    .Q(\mem[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3785_ (.CLK(clknet_leaf_26_clk),
    .D(net485),
    .Q(\mem[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3786_ (.CLK(clknet_leaf_26_clk),
    .D(net535),
    .Q(\mem[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3787_ (.CLK(clknet_leaf_30_clk),
    .D(net651),
    .Q(\mem[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3788_ (.CLK(clknet_leaf_90_clk),
    .D(net1247),
    .Q(\mem[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3789_ (.CLK(clknet_leaf_81_clk),
    .D(net1505),
    .Q(\mem[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3790_ (.CLK(clknet_leaf_88_clk),
    .D(net2003),
    .Q(\mem[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3791_ (.CLK(clknet_leaf_15_clk),
    .D(net883),
    .Q(\mem[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3792_ (.CLK(clknet_leaf_86_clk),
    .D(net1951),
    .Q(\mem[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3793_ (.CLK(clknet_leaf_11_clk),
    .D(net2051),
    .Q(\mem[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3794_ (.CLK(clknet_leaf_81_clk),
    .D(net1861),
    .Q(\mem[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3795_ (.CLK(clknet_leaf_11_clk),
    .D(net1393),
    .Q(\mem[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3796_ (.CLK(clknet_leaf_9_clk),
    .D(net2321),
    .Q(\mem[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3797_ (.CLK(clknet_leaf_14_clk),
    .D(net1117),
    .Q(\mem[24][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3798_ (.CLK(clknet_leaf_31_clk),
    .D(net1269),
    .Q(\mem[24][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3799_ (.CLK(clknet_leaf_81_clk),
    .D(net2281),
    .Q(\mem[24][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3800_ (.CLK(clknet_leaf_33_clk),
    .D(net1675),
    .Q(\mem[24][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3801_ (.CLK(clknet_leaf_13_clk),
    .D(net589),
    .Q(\mem[24][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3802_ (.CLK(clknet_leaf_8_clk),
    .D(net983),
    .Q(\mem[24][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3803_ (.CLK(clknet_leaf_85_clk),
    .D(net1287),
    .Q(\mem[24][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3804_ (.CLK(clknet_leaf_87_clk),
    .D(net641),
    .Q(\mem[24][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3805_ (.CLK(clknet_leaf_88_clk),
    .D(net1643),
    .Q(\mem[24][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3806_ (.CLK(clknet_leaf_87_clk),
    .D(net2107),
    .Q(\mem[24][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3807_ (.CLK(clknet_leaf_85_clk),
    .D(net1711),
    .Q(\mem[24][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3808_ (.CLK(clknet_leaf_13_clk),
    .D(net805),
    .Q(\mem[24][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3809_ (.CLK(clknet_leaf_7_clk),
    .D(net1275),
    .Q(\mem[24][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3810_ (.CLK(clknet_leaf_88_clk),
    .D(net1973),
    .Q(\mem[24][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3811_ (.CLK(clknet_leaf_91_clk),
    .D(net623),
    .Q(\mem[24][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3812_ (.CLK(clknet_leaf_33_clk),
    .D(net1317),
    .Q(\mem[24][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3813_ (.CLK(clknet_leaf_27_clk),
    .D(net447),
    .Q(\mem[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3814_ (.CLK(clknet_leaf_28_clk),
    .D(net637),
    .Q(\mem[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3815_ (.CLK(clknet_leaf_89_clk),
    .D(net2405),
    .Q(\mem[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3816_ (.CLK(clknet_leaf_10_clk),
    .D(net2381),
    .Q(\mem[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3817_ (.CLK(clknet_leaf_40_clk),
    .D(net579),
    .Q(\mem[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3818_ (.CLK(clknet_leaf_27_clk),
    .D(net491),
    .Q(\mem[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3819_ (.CLK(clknet_leaf_30_clk),
    .D(net1595),
    .Q(\mem[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3820_ (.CLK(clknet_leaf_8_clk),
    .D(net1657),
    .Q(\mem[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3821_ (.CLK(clknet_leaf_10_clk),
    .D(net2309),
    .Q(\mem[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3822_ (.CLK(clknet_leaf_89_clk),
    .D(net2033),
    .Q(\mem[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3823_ (.CLK(clknet_leaf_6_clk),
    .D(net1825),
    .Q(\mem[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3824_ (.CLK(clknet_leaf_86_clk),
    .D(net1995),
    .Q(\mem[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3825_ (.CLK(clknet_leaf_11_clk),
    .D(net2127),
    .Q(\mem[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3826_ (.CLK(clknet_leaf_81_clk),
    .D(net2343),
    .Q(\mem[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3827_ (.CLK(clknet_leaf_12_clk),
    .D(net2371),
    .Q(\mem[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3828_ (.CLK(clknet_leaf_9_clk),
    .D(net2329),
    .Q(\mem[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3829_ (.CLK(clknet_leaf_13_clk),
    .D(net1307),
    .Q(\mem[31][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3830_ (.CLK(clknet_leaf_32_clk),
    .D(net2253),
    .Q(\mem[31][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3831_ (.CLK(clknet_leaf_81_clk),
    .D(net2151),
    .Q(\mem[31][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3832_ (.CLK(clknet_leaf_32_clk),
    .D(net1703),
    .Q(\mem[31][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3833_ (.CLK(clknet_leaf_20_clk),
    .D(net2351),
    .Q(\mem[31][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3834_ (.CLK(clknet_leaf_8_clk),
    .D(net1775),
    .Q(\mem[31][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3835_ (.CLK(clknet_leaf_82_clk),
    .D(net1551),
    .Q(\mem[31][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3836_ (.CLK(clknet_leaf_86_clk),
    .D(net1779),
    .Q(\mem[31][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3837_ (.CLK(clknet_leaf_89_clk),
    .D(net2187),
    .Q(\mem[31][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3838_ (.CLK(clknet_leaf_85_clk),
    .D(net1693),
    .Q(\mem[31][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3839_ (.CLK(clknet_leaf_85_clk),
    .D(net2101),
    .Q(\mem[31][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3840_ (.CLK(clknet_leaf_13_clk),
    .D(net1299),
    .Q(\mem[31][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3841_ (.CLK(clknet_leaf_7_clk),
    .D(net2161),
    .Q(\mem[31][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3842_ (.CLK(clknet_leaf_89_clk),
    .D(net1987),
    .Q(\mem[31][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3843_ (.CLK(clknet_leaf_91_clk),
    .D(net2387),
    .Q(\mem[31][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3844_ (.CLK(clknet_leaf_33_clk),
    .D(net1921),
    .Q(\mem[31][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3845_ (.CLK(clknet_leaf_25_clk),
    .D(net425),
    .Q(\mem[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3846_ (.CLK(clknet_leaf_26_clk),
    .D(net397),
    .Q(\mem[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3847_ (.CLK(clknet_leaf_92_clk),
    .D(net795),
    .Q(\mem[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3848_ (.CLK(clknet_leaf_10_clk),
    .D(net2219),
    .Q(\mem[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3849_ (.CLK(clknet_leaf_26_clk),
    .D(net413),
    .Q(\mem[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3850_ (.CLK(clknet_leaf_25_clk),
    .D(net403),
    .Q(\mem[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3851_ (.CLK(clknet_leaf_12_clk),
    .D(net957),
    .Q(\mem[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3852_ (.CLK(clknet_leaf_90_clk),
    .D(net1159),
    .Q(\mem[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3853_ (.CLK(clknet_leaf_81_clk),
    .D(net2055),
    .Q(\mem[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3854_ (.CLK(clknet_leaf_88_clk),
    .D(net1415),
    .Q(\mem[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3855_ (.CLK(clknet_leaf_14_clk),
    .D(net1225),
    .Q(\mem[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3856_ (.CLK(clknet_leaf_86_clk),
    .D(net1091),
    .Q(\mem[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3857_ (.CLK(clknet_leaf_11_clk),
    .D(net1395),
    .Q(\mem[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3858_ (.CLK(clknet_leaf_81_clk),
    .D(net2109),
    .Q(\mem[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3859_ (.CLK(clknet_leaf_11_clk),
    .D(net2225),
    .Q(\mem[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3860_ (.CLK(clknet_leaf_6_clk),
    .D(net1081),
    .Q(\mem[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3861_ (.CLK(clknet_leaf_14_clk),
    .D(net2167),
    .Q(\mem[25][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3862_ (.CLK(clknet_leaf_32_clk),
    .D(net929),
    .Q(\mem[25][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3863_ (.CLK(clknet_leaf_81_clk),
    .D(net1943),
    .Q(\mem[25][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3864_ (.CLK(clknet_leaf_32_clk),
    .D(net687),
    .Q(\mem[25][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3865_ (.CLK(clknet_leaf_20_clk),
    .D(net1541),
    .Q(\mem[25][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3866_ (.CLK(clknet_leaf_8_clk),
    .D(net701),
    .Q(\mem[25][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3867_ (.CLK(clknet_leaf_85_clk),
    .D(net639),
    .Q(\mem[25][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3868_ (.CLK(clknet_leaf_87_clk),
    .D(net1079),
    .Q(\mem[25][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3869_ (.CLK(clknet_leaf_88_clk),
    .D(net1865),
    .Q(\mem[25][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3870_ (.CLK(clknet_leaf_86_clk),
    .D(net1011),
    .Q(\mem[25][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3871_ (.CLK(clknet_leaf_84_clk),
    .D(net1131),
    .Q(\mem[25][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3872_ (.CLK(clknet_leaf_12_clk),
    .D(net2043),
    .Q(\mem[25][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3873_ (.CLK(clknet_leaf_7_clk),
    .D(net2037),
    .Q(\mem[25][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3874_ (.CLK(clknet_leaf_88_clk),
    .D(net1937),
    .Q(\mem[25][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3875_ (.CLK(clknet_leaf_91_clk),
    .D(net1361),
    .Q(\mem[25][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3876_ (.CLK(clknet_leaf_33_clk),
    .D(net1153),
    .Q(\mem[25][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3877_ (.CLK(clknet_leaf_25_clk),
    .D(net533),
    .Q(\mem[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3878_ (.CLK(clknet_leaf_27_clk),
    .D(net381),
    .Q(\mem[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3879_ (.CLK(clknet_leaf_92_clk),
    .D(net917),
    .Q(\mem[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3880_ (.CLK(clknet_leaf_10_clk),
    .D(net1975),
    .Q(\mem[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3881_ (.CLK(clknet_leaf_25_clk),
    .D(net405),
    .Q(\mem[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3882_ (.CLK(clknet_leaf_25_clk),
    .D(net577),
    .Q(\mem[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3883_ (.CLK(clknet_leaf_30_clk),
    .D(net807),
    .Q(\mem[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3884_ (.CLK(clknet_leaf_0_clk),
    .D(net1215),
    .Q(\mem[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3885_ (.CLK(clknet_leaf_10_clk),
    .D(net1853),
    .Q(\mem[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3886_ (.CLK(clknet_leaf_88_clk),
    .D(net1365),
    .Q(\mem[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3887_ (.CLK(clknet_leaf_15_clk),
    .D(net625),
    .Q(\mem[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3888_ (.CLK(clknet_leaf_87_clk),
    .D(net1385),
    .Q(\mem[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3889_ (.CLK(clknet_leaf_14_clk),
    .D(net1271),
    .Q(\mem[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3890_ (.CLK(clknet_leaf_81_clk),
    .D(net2331),
    .Q(\mem[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3891_ (.CLK(clknet_leaf_11_clk),
    .D(net2015),
    .Q(\mem[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3892_ (.CLK(clknet_leaf_6_clk),
    .D(net893),
    .Q(\mem[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3893_ (.CLK(clknet_leaf_14_clk),
    .D(net715),
    .Q(\mem[27][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3894_ (.CLK(clknet_leaf_31_clk),
    .D(net1725),
    .Q(\mem[27][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3895_ (.CLK(clknet_leaf_81_clk),
    .D(net1993),
    .Q(\mem[27][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3896_ (.CLK(clknet_leaf_33_clk),
    .D(net1025),
    .Q(\mem[27][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3897_ (.CLK(clknet_leaf_20_clk),
    .D(net1409),
    .Q(\mem[27][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3898_ (.CLK(clknet_leaf_7_clk),
    .D(net1545),
    .Q(\mem[27][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3899_ (.CLK(clknet_leaf_86_clk),
    .D(net1579),
    .Q(\mem[27][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3900_ (.CLK(clknet_leaf_88_clk),
    .D(net1149),
    .Q(\mem[27][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3901_ (.CLK(clknet_leaf_88_clk),
    .D(net2089),
    .Q(\mem[27][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3902_ (.CLK(clknet_leaf_87_clk),
    .D(net1649),
    .Q(\mem[27][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3903_ (.CLK(clknet_leaf_84_clk),
    .D(net2233),
    .Q(\mem[27][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3904_ (.CLK(clknet_leaf_13_clk),
    .D(net633),
    .Q(\mem[27][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3905_ (.CLK(clknet_leaf_5_clk),
    .D(net1213),
    .Q(\mem[27][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3906_ (.CLK(clknet_leaf_92_clk),
    .D(net667),
    .Q(\mem[27][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3907_ (.CLK(clknet_leaf_92_clk),
    .D(net663),
    .Q(\mem[27][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3908_ (.CLK(clknet_leaf_10_clk),
    .D(net2153),
    .Q(\mem[27][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3909_ (.CLK(clknet_leaf_39_clk),
    .D(net411),
    .Q(\mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3910_ (.CLK(clknet_leaf_40_clk),
    .D(net373),
    .Q(\mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3911_ (.CLK(clknet_leaf_78_clk),
    .D(net1841),
    .Q(\mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3912_ (.CLK(clknet_leaf_55_clk),
    .D(net693),
    .Q(\mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3913_ (.CLK(clknet_leaf_39_clk),
    .D(net461),
    .Q(\mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3914_ (.CLK(clknet_leaf_39_clk),
    .D(net459),
    .Q(\mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3915_ (.CLK(clknet_leaf_47_clk),
    .D(net1659),
    .Q(\mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3916_ (.CLK(clknet_leaf_65_clk),
    .D(net1695),
    .Q(\mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3917_ (.CLK(clknet_leaf_57_clk),
    .D(net1645),
    .Q(\mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3918_ (.CLK(clknet_leaf_64_clk),
    .D(net759),
    .Q(\mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3919_ (.CLK(clknet_leaf_48_clk),
    .D(net861),
    .Q(\mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3920_ (.CLK(clknet_leaf_77_clk),
    .D(net869),
    .Q(\mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3921_ (.CLK(clknet_leaf_37_clk),
    .D(net1101),
    .Q(\mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3922_ (.CLK(clknet_leaf_64_clk),
    .D(net1487),
    .Q(\mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3923_ (.CLK(clknet_leaf_47_clk),
    .D(net2113),
    .Q(\mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3924_ (.CLK(clknet_leaf_62_clk),
    .D(net1013),
    .Q(\mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3925_ (.CLK(clknet_leaf_55_clk),
    .D(net723),
    .Q(\mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3926_ (.CLK(clknet_leaf_47_clk),
    .D(net1753),
    .Q(\mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3927_ (.CLK(clknet_leaf_59_clk),
    .D(net1469),
    .Q(\mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3928_ (.CLK(clknet_leaf_47_clk),
    .D(net1663),
    .Q(\mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3929_ (.CLK(clknet_leaf_52_clk),
    .D(net1997),
    .Q(\mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3930_ (.CLK(clknet_leaf_63_clk),
    .D(net771),
    .Q(\mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3931_ (.CLK(clknet_leaf_59_clk),
    .D(net2121),
    .Q(\mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3932_ (.CLK(clknet_leaf_65_clk),
    .D(net1953),
    .Q(\mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3933_ (.CLK(clknet_leaf_76_clk),
    .D(net2085),
    .Q(\mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3934_ (.CLK(clknet_leaf_77_clk),
    .D(net1391),
    .Q(\mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3935_ (.CLK(clknet_leaf_56_clk),
    .D(net1111),
    .Q(\mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3936_ (.CLK(clknet_leaf_52_clk),
    .D(net1899),
    .Q(\mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3937_ (.CLK(clknet_leaf_58_clk),
    .D(net1911),
    .Q(\mem[3][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3938_ (.CLK(clknet_leaf_78_clk),
    .D(net1169),
    .Q(\mem[3][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3939_ (.CLK(clknet_leaf_78_clk),
    .D(net1615),
    .Q(\mem[3][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3940_ (.CLK(clknet_leaf_54_clk),
    .D(net2163),
    .Q(\mem[3][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3941_ (.CLK(clknet_leaf_28_clk),
    .D(net559),
    .Q(\mem[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3942_ (.CLK(clknet_leaf_28_clk),
    .D(net465),
    .Q(\mem[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3943_ (.CLK(clknet_leaf_91_clk),
    .D(net691),
    .Q(\mem[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3944_ (.CLK(clknet_leaf_10_clk),
    .D(net2407),
    .Q(\mem[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3945_ (.CLK(clknet_leaf_27_clk),
    .D(net565),
    .Q(\mem[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3946_ (.CLK(clknet_leaf_28_clk),
    .D(net561),
    .Q(\mem[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3947_ (.CLK(clknet_leaf_22_clk),
    .D(net1383),
    .Q(\mem[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3948_ (.CLK(clknet_leaf_0_clk),
    .D(net2099),
    .Q(\mem[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3949_ (.CLK(clknet_leaf_10_clk),
    .D(net2357),
    .Q(\mem[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3950_ (.CLK(clknet_leaf_88_clk),
    .D(net2115),
    .Q(\mem[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3951_ (.CLK(clknet_leaf_5_clk),
    .D(net1527),
    .Q(\mem[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3952_ (.CLK(clknet_leaf_87_clk),
    .D(net1601),
    .Q(\mem[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3953_ (.CLK(clknet_leaf_6_clk),
    .D(net1371),
    .Q(\mem[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3954_ (.CLK(clknet_leaf_81_clk),
    .D(net2013),
    .Q(\mem[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3955_ (.CLK(clknet_leaf_12_clk),
    .D(net1985),
    .Q(\mem[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3956_ (.CLK(clknet_leaf_9_clk),
    .D(net2299),
    .Q(\mem[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3957_ (.CLK(clknet_leaf_14_clk),
    .D(net1851),
    .Q(\mem[28][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3958_ (.CLK(clknet_leaf_32_clk),
    .D(net1139),
    .Q(\mem[28][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3959_ (.CLK(clknet_leaf_81_clk),
    .D(net2265),
    .Q(\mem[28][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3960_ (.CLK(clknet_leaf_35_clk),
    .D(net1465),
    .Q(\mem[28][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3961_ (.CLK(clknet_leaf_22_clk),
    .D(net2035),
    .Q(\mem[28][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3962_ (.CLK(clknet_leaf_8_clk),
    .D(net2271),
    .Q(\mem[28][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3963_ (.CLK(clknet_leaf_79_clk),
    .D(net2069),
    .Q(\mem[28][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3964_ (.CLK(clknet_leaf_87_clk),
    .D(net1513),
    .Q(\mem[28][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3965_ (.CLK(clknet_leaf_89_clk),
    .D(net1537),
    .Q(\mem[28][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3966_ (.CLK(clknet_leaf_73_clk),
    .D(net2041),
    .Q(\mem[28][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3967_ (.CLK(clknet_leaf_74_clk),
    .D(net1941),
    .Q(\mem[28][26] ));
 sky130_fd_sc_hd__dfxtp_1 _3968_ (.CLK(clknet_leaf_20_clk),
    .D(net1885),
    .Q(\mem[28][27] ));
 sky130_fd_sc_hd__dfxtp_1 _3969_ (.CLK(clknet_leaf_7_clk),
    .D(net793),
    .Q(\mem[28][28] ));
 sky130_fd_sc_hd__dfxtp_1 _3970_ (.CLK(clknet_leaf_88_clk),
    .D(net2213),
    .Q(\mem[28][29] ));
 sky130_fd_sc_hd__dfxtp_1 _3971_ (.CLK(clknet_leaf_92_clk),
    .D(net1557),
    .Q(\mem[28][30] ));
 sky130_fd_sc_hd__dfxtp_1 _3972_ (.CLK(clknet_leaf_34_clk),
    .D(net1263),
    .Q(\mem[28][31] ));
 sky130_fd_sc_hd__dfxtp_1 _3973_ (.CLK(clknet_leaf_39_clk),
    .D(net511),
    .Q(\mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _3974_ (.CLK(clknet_leaf_40_clk),
    .D(net391),
    .Q(\mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _3975_ (.CLK(clknet_leaf_75_clk),
    .D(net635),
    .Q(\mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _3976_ (.CLK(clknet_leaf_55_clk),
    .D(net987),
    .Q(\mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _3977_ (.CLK(clknet_leaf_39_clk),
    .D(net591),
    .Q(\mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _3978_ (.CLK(clknet_leaf_40_clk),
    .D(net551),
    .Q(\mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _3979_ (.CLK(clknet_leaf_47_clk),
    .D(net1531),
    .Q(\mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _3980_ (.CLK(clknet_leaf_65_clk),
    .D(net1905),
    .Q(\mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _3981_ (.CLK(clknet_leaf_57_clk),
    .D(net729),
    .Q(\mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _3982_ (.CLK(clknet_leaf_67_clk),
    .D(net613),
    .Q(\mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _3983_ (.CLK(clknet_leaf_62_clk),
    .D(net1745),
    .Q(\mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _3984_ (.CLK(clknet_leaf_77_clk),
    .D(net1355),
    .Q(\mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _3985_ (.CLK(clknet_leaf_37_clk),
    .D(net655),
    .Q(\mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _3986_ (.CLK(clknet_leaf_64_clk),
    .D(net1115),
    .Q(\mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _3987_ (.CLK(clknet_leaf_47_clk),
    .D(net1833),
    .Q(\mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _3988_ (.CLK(clknet_leaf_62_clk),
    .D(net1241),
    .Q(\mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _3989_ (.CLK(clknet_leaf_35_clk),
    .D(net821),
    .Q(\mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 _3990_ (.CLK(clknet_leaf_47_clk),
    .D(net1477),
    .Q(\mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 _3991_ (.CLK(clknet_leaf_58_clk),
    .D(net1625),
    .Q(\mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 _3992_ (.CLK(clknet_leaf_48_clk),
    .D(net2257),
    .Q(\mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 _3993_ (.CLK(clknet_leaf_51_clk),
    .D(net1491),
    .Q(\mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 _3994_ (.CLK(clknet_leaf_63_clk),
    .D(net803),
    .Q(\mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 _3995_ (.CLK(clknet_leaf_59_clk),
    .D(net1895),
    .Q(\mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 _3996_ (.CLK(clknet_leaf_65_clk),
    .D(net1443),
    .Q(\mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 _3997_ (.CLK(clknet_leaf_76_clk),
    .D(net1337),
    .Q(\mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 _3998_ (.CLK(clknet_leaf_77_clk),
    .D(net1903),
    .Q(\mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 _3999_ (.CLK(clknet_leaf_56_clk),
    .D(net2071),
    .Q(\mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4000_ (.CLK(clknet_leaf_52_clk),
    .D(net1501),
    .Q(\mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4001_ (.CLK(clknet_leaf_78_clk),
    .D(net959),
    .Q(\mem[2][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4002_ (.CLK(clknet_leaf_78_clk),
    .D(net1017),
    .Q(\mem[2][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4003_ (.CLK(clknet_leaf_78_clk),
    .D(net1727),
    .Q(\mem[2][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4004_ (.CLK(clknet_leaf_54_clk),
    .D(net1721),
    .Q(\mem[2][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4005_ (.CLK(clknet_leaf_28_clk),
    .D(net483),
    .Q(\mem[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4006_ (.CLK(clknet_leaf_29_clk),
    .D(net503),
    .Q(\mem[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4007_ (.CLK(clknet_leaf_0_clk),
    .D(net2413),
    .Q(\mem[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4008_ (.CLK(clknet_leaf_5_clk),
    .D(net2303),
    .Q(\mem[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4009_ (.CLK(clknet_leaf_24_clk),
    .D(net573),
    .Q(\mem[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4010_ (.CLK(clknet_leaf_25_clk),
    .D(net455),
    .Q(\mem[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4011_ (.CLK(clknet_leaf_21_clk),
    .D(net1571),
    .Q(\mem[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4012_ (.CLK(clknet_leaf_2_clk),
    .D(net2295),
    .Q(\mem[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4013_ (.CLK(clknet_leaf_11_clk),
    .D(net1883),
    .Q(\mem[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4014_ (.CLK(clknet_leaf_89_clk),
    .D(net2379),
    .Q(\mem[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4015_ (.CLK(clknet_leaf_5_clk),
    .D(net1617),
    .Q(\mem[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4016_ (.CLK(clknet_leaf_89_clk),
    .D(net2393),
    .Q(\mem[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4017_ (.CLK(clknet_leaf_17_clk),
    .D(net1071),
    .Q(\mem[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4018_ (.CLK(clknet_leaf_9_clk),
    .D(net2377),
    .Q(\mem[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4019_ (.CLK(clknet_leaf_20_clk),
    .D(net2235),
    .Q(\mem[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4020_ (.CLK(clknet_leaf_5_clk),
    .D(net2369),
    .Q(\mem[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4021_ (.CLK(clknet_leaf_18_clk),
    .D(net1963),
    .Q(\mem[19][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4022_ (.CLK(clknet_leaf_30_clk),
    .D(net1613),
    .Q(\mem[19][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4023_ (.CLK(clknet_leaf_83_clk),
    .D(net2217),
    .Q(\mem[19][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4024_ (.CLK(clknet_leaf_11_clk),
    .D(net2307),
    .Q(\mem[19][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4025_ (.CLK(clknet_leaf_20_clk),
    .D(net2403),
    .Q(\mem[19][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4026_ (.CLK(clknet_leaf_6_clk),
    .D(net1813),
    .Q(\mem[19][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4027_ (.CLK(clknet_leaf_89_clk),
    .D(net2123),
    .Q(\mem[19][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4028_ (.CLK(clknet_leaf_83_clk),
    .D(net2201),
    .Q(\mem[19][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4029_ (.CLK(clknet_leaf_93_clk),
    .D(net973),
    .Q(\mem[19][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4030_ (.CLK(clknet_leaf_84_clk),
    .D(net2383),
    .Q(\mem[19][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4031_ (.CLK(clknet_leaf_3_clk),
    .D(net1051),
    .Q(\mem[19][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4032_ (.CLK(clknet_leaf_21_clk),
    .D(net867),
    .Q(\mem[19][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4033_ (.CLK(clknet_leaf_4_clk),
    .D(net1535),
    .Q(\mem[19][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4034_ (.CLK(clknet_leaf_0_clk),
    .D(net1737),
    .Q(\mem[19][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4035_ (.CLK(clknet_leaf_2_clk),
    .D(net1717),
    .Q(\mem[19][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4036_ (.CLK(clknet_leaf_11_clk),
    .D(net2339),
    .Q(\mem[19][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4037_ (.CLK(clknet_leaf_22_clk),
    .D(net1077),
    .Q(\mem[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4038_ (.CLK(clknet_leaf_29_clk),
    .D(net479),
    .Q(\mem[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4039_ (.CLK(clknet_leaf_0_clk),
    .D(net2155),
    .Q(\mem[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4040_ (.CLK(clknet_leaf_16_clk),
    .D(net2237),
    .Q(\mem[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4041_ (.CLK(clknet_leaf_22_clk),
    .D(net527),
    .Q(\mem[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4042_ (.CLK(clknet_leaf_22_clk),
    .D(net603),
    .Q(\mem[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4043_ (.CLK(clknet_leaf_20_clk),
    .D(net1879),
    .Q(\mem[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4044_ (.CLK(clknet_leaf_0_clk),
    .D(net2293),
    .Q(\mem[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4045_ (.CLK(clknet_leaf_9_clk),
    .D(net2401),
    .Q(\mem[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4046_ (.CLK(clknet_leaf_89_clk),
    .D(net2039),
    .Q(\mem[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4047_ (.CLK(clknet_leaf_5_clk),
    .D(net2091),
    .Q(\mem[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4048_ (.CLK(clknet_leaf_84_clk),
    .D(net1553),
    .Q(\mem[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4049_ (.CLK(clknet_leaf_16_clk),
    .D(net1681),
    .Q(\mem[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4050_ (.CLK(clknet_leaf_81_clk),
    .D(net2399),
    .Q(\mem[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4051_ (.CLK(clknet_leaf_19_clk),
    .D(net1935),
    .Q(\mem[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4052_ (.CLK(clknet_leaf_5_clk),
    .D(net2189),
    .Q(\mem[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4053_ (.CLK(clknet_leaf_14_clk),
    .D(net1927),
    .Q(\mem[17][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4054_ (.CLK(clknet_leaf_31_clk),
    .D(net1475),
    .Q(\mem[17][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4055_ (.CLK(clknet_leaf_81_clk),
    .D(net2185),
    .Q(\mem[17][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4056_ (.CLK(clknet_leaf_31_clk),
    .D(net2073),
    .Q(\mem[17][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4057_ (.CLK(clknet_leaf_20_clk),
    .D(net2275),
    .Q(\mem[17][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4058_ (.CLK(clknet_leaf_9_clk),
    .D(net2415),
    .Q(\mem[17][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4059_ (.CLK(clknet_leaf_84_clk),
    .D(net1809),
    .Q(\mem[17][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4060_ (.CLK(clknet_leaf_82_clk),
    .D(net1347),
    .Q(\mem[17][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4061_ (.CLK(clknet_leaf_0_clk),
    .D(net2131),
    .Q(\mem[17][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4062_ (.CLK(clknet_leaf_84_clk),
    .D(net2391),
    .Q(\mem[17][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4063_ (.CLK(clknet_leaf_2_clk),
    .D(net1439),
    .Q(\mem[17][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4064_ (.CLK(clknet_leaf_19_clk),
    .D(net899),
    .Q(\mem[17][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4065_ (.CLK(clknet_leaf_7_clk),
    .D(net1447),
    .Q(\mem[17][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4066_ (.CLK(clknet_leaf_1_clk),
    .D(net1815),
    .Q(\mem[17][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4067_ (.CLK(clknet_leaf_1_clk),
    .D(net1967),
    .Q(\mem[17][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4068_ (.CLK(clknet_leaf_11_clk),
    .D(net2373),
    .Q(\mem[17][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4069_ (.CLK(clknet_leaf_43_clk),
    .D(net881),
    .Q(\mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4070_ (.CLK(clknet_leaf_43_clk),
    .D(net581),
    .Q(\mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4071_ (.CLK(clknet_leaf_74_clk),
    .D(net971),
    .Q(\mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4072_ (.CLK(clknet_leaf_55_clk),
    .D(net1407),
    .Q(\mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4073_ (.CLK(clknet_leaf_43_clk),
    .D(net517),
    .Q(\mem[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4074_ (.CLK(clknet_leaf_43_clk),
    .D(net605),
    .Q(\mem[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4075_ (.CLK(clknet_leaf_45_clk),
    .D(net1961),
    .Q(\mem[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4076_ (.CLK(clknet_leaf_66_clk),
    .D(net685),
    .Q(\mem[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4077_ (.CLK(clknet_leaf_54_clk),
    .D(net747),
    .Q(\mem[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4078_ (.CLK(clknet_leaf_70_clk),
    .D(net1009),
    .Q(\mem[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4079_ (.CLK(clknet_leaf_48_clk),
    .D(net1751),
    .Q(\mem[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4080_ (.CLK(clknet_leaf_71_clk),
    .D(net1685),
    .Q(\mem[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4081_ (.CLK(clknet_leaf_36_clk),
    .D(net617),
    .Q(\mem[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4082_ (.CLK(clknet_leaf_65_clk),
    .D(net1291),
    .Q(\mem[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4083_ (.CLK(clknet_leaf_47_clk),
    .D(net2283),
    .Q(\mem[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4084_ (.CLK(clknet_leaf_62_clk),
    .D(net1423),
    .Q(\mem[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4085_ (.CLK(clknet_leaf_34_clk),
    .D(net675),
    .Q(\mem[6][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4086_ (.CLK(clknet_leaf_45_clk),
    .D(net1175),
    .Q(\mem[6][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4087_ (.CLK(clknet_leaf_58_clk),
    .D(net2359),
    .Q(\mem[6][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4088_ (.CLK(clknet_leaf_48_clk),
    .D(net1069),
    .Q(\mem[6][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4089_ (.CLK(clknet_leaf_44_clk),
    .D(net2047),
    .Q(\mem[6][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4090_ (.CLK(clknet_leaf_62_clk),
    .D(net1221),
    .Q(\mem[6][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4091_ (.CLK(clknet_leaf_71_clk),
    .D(net2029),
    .Q(\mem[6][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4092_ (.CLK(clknet_leaf_67_clk),
    .D(net1485),
    .Q(\mem[6][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4093_ (.CLK(clknet_leaf_72_clk),
    .D(net2313),
    .Q(\mem[6][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4094_ (.CLK(clknet_leaf_71_clk),
    .D(net2367),
    .Q(\mem[6][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4095_ (.CLK(clknet_leaf_56_clk),
    .D(net2171),
    .Q(\mem[6][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4096_ (.CLK(clknet_leaf_38_clk),
    .D(net741),
    .Q(\mem[6][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4097_ (.CLK(clknet_leaf_79_clk),
    .D(net739),
    .Q(\mem[6][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4098_ (.CLK(clknet_leaf_74_clk),
    .D(net2145),
    .Q(\mem[6][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4099_ (.CLK(clknet_leaf_79_clk),
    .D(net1623),
    .Q(\mem[6][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4100_ (.CLK(clknet_leaf_53_clk),
    .D(net787),
    .Q(\mem[6][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4101_ (.CLK(clknet_leaf_27_clk),
    .D(net509),
    .Q(\mem[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4102_ (.CLK(clknet_leaf_28_clk),
    .D(net467),
    .Q(\mem[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4103_ (.CLK(clknet_leaf_91_clk),
    .D(net1881),
    .Q(\mem[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4104_ (.CLK(clknet_leaf_10_clk),
    .D(net2227),
    .Q(\mem[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4105_ (.CLK(clknet_leaf_27_clk),
    .D(net583),
    .Q(\mem[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4106_ (.CLK(clknet_leaf_27_clk),
    .D(net727),
    .Q(\mem[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4107_ (.CLK(clknet_leaf_22_clk),
    .D(net2315),
    .Q(\mem[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4108_ (.CLK(clknet_leaf_0_clk),
    .D(net1959),
    .Q(\mem[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4109_ (.CLK(clknet_leaf_10_clk),
    .D(net2417),
    .Q(\mem[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4110_ (.CLK(clknet_leaf_88_clk),
    .D(net2143),
    .Q(\mem[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4111_ (.CLK(clknet_leaf_5_clk),
    .D(net1673),
    .Q(\mem[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4112_ (.CLK(clknet_leaf_73_clk),
    .D(net1611),
    .Q(\mem[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4113_ (.CLK(clknet_leaf_15_clk),
    .D(net1387),
    .Q(\mem[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4114_ (.CLK(clknet_leaf_81_clk),
    .D(net2349),
    .Q(\mem[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4115_ (.CLK(clknet_leaf_12_clk),
    .D(net2361),
    .Q(\mem[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4116_ (.CLK(clknet_leaf_9_clk),
    .D(net2333),
    .Q(\mem[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4117_ (.CLK(clknet_leaf_14_clk),
    .D(net1863),
    .Q(\mem[29][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4118_ (.CLK(clknet_leaf_32_clk),
    .D(net1983),
    .Q(\mem[29][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4119_ (.CLK(clknet_leaf_81_clk),
    .D(net2159),
    .Q(\mem[29][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4120_ (.CLK(clknet_leaf_32_clk),
    .D(net2077),
    .Q(\mem[29][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4121_ (.CLK(clknet_leaf_22_clk),
    .D(net2239),
    .Q(\mem[29][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4122_ (.CLK(clknet_leaf_8_clk),
    .D(net2301),
    .Q(\mem[29][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4123_ (.CLK(clknet_leaf_82_clk),
    .D(net819),
    .Q(\mem[29][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4124_ (.CLK(clknet_leaf_87_clk),
    .D(net1821),
    .Q(\mem[29][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4125_ (.CLK(clknet_leaf_88_clk),
    .D(net2335),
    .Q(\mem[29][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4126_ (.CLK(clknet_leaf_86_clk),
    .D(net1677),
    .Q(\mem[29][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4127_ (.CLK(clknet_leaf_85_clk),
    .D(net1459),
    .Q(\mem[29][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4128_ (.CLK(clknet_leaf_13_clk),
    .D(net1789),
    .Q(\mem[29][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4129_ (.CLK(clknet_leaf_7_clk),
    .D(net2215),
    .Q(\mem[29][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4130_ (.CLK(clknet_leaf_88_clk),
    .D(net1933),
    .Q(\mem[29][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4131_ (.CLK(clknet_leaf_92_clk),
    .D(net1479),
    .Q(\mem[29][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4132_ (.CLK(clknet_leaf_10_clk),
    .D(net2365),
    .Q(\mem[29][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4133_ (.CLK(clknet_leaf_41_clk),
    .D(net523),
    .Q(\mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4134_ (.CLK(clknet_leaf_40_clk),
    .D(net487),
    .Q(\mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4135_ (.CLK(clknet_leaf_74_clk),
    .D(net1357),
    .Q(\mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4136_ (.CLK(clknet_leaf_55_clk),
    .D(net683),
    .Q(\mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4137_ (.CLK(clknet_leaf_41_clk),
    .D(net501),
    .Q(\mem[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4138_ (.CLK(clknet_leaf_42_clk),
    .D(net385),
    .Q(\mem[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4139_ (.CLK(clknet_leaf_46_clk),
    .D(net1991),
    .Q(\mem[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4140_ (.CLK(clknet_leaf_65_clk),
    .D(net2311),
    .Q(\mem[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4141_ (.CLK(clknet_leaf_57_clk),
    .D(net2183),
    .Q(\mem[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4142_ (.CLK(clknet_leaf_67_clk),
    .D(net783),
    .Q(\mem[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4143_ (.CLK(clknet_leaf_49_clk),
    .D(net1835),
    .Q(\mem[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4144_ (.CLK(clknet_leaf_71_clk),
    .D(net2375),
    .Q(\mem[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4145_ (.CLK(clknet_leaf_35_clk),
    .D(net1555),
    .Q(\mem[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4146_ (.CLK(clknet_leaf_65_clk),
    .D(net2263),
    .Q(\mem[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4147_ (.CLK(clknet_leaf_51_clk),
    .D(net1031),
    .Q(\mem[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4148_ (.CLK(clknet_leaf_61_clk),
    .D(net1003),
    .Q(\mem[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4149_ (.CLK(clknet_leaf_35_clk),
    .D(net2197),
    .Q(\mem[8][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4150_ (.CLK(clknet_leaf_45_clk),
    .D(net951),
    .Q(\mem[8][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4151_ (.CLK(clknet_leaf_58_clk),
    .D(net1877),
    .Q(\mem[8][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4152_ (.CLK(clknet_leaf_49_clk),
    .D(net877),
    .Q(\mem[8][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4153_ (.CLK(clknet_leaf_45_clk),
    .D(net1581),
    .Q(\mem[8][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4154_ (.CLK(clknet_leaf_62_clk),
    .D(net1155),
    .Q(\mem[8][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4155_ (.CLK(clknet_leaf_65_clk),
    .D(net1195),
    .Q(\mem[8][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4156_ (.CLK(clknet_leaf_65_clk),
    .D(net1917),
    .Q(\mem[8][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4157_ (.CLK(clknet_leaf_71_clk),
    .D(net2345),
    .Q(\mem[8][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4158_ (.CLK(clknet_leaf_71_clk),
    .D(net2063),
    .Q(\mem[8][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4159_ (.CLK(clknet_leaf_56_clk),
    .D(net1891),
    .Q(\mem[8][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4160_ (.CLK(clknet_leaf_44_clk),
    .D(net1793),
    .Q(\mem[8][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4161_ (.CLK(clknet_leaf_80_clk),
    .D(net1321),
    .Q(\mem[8][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4162_ (.CLK(clknet_leaf_75_clk),
    .D(net2195),
    .Q(\mem[8][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4163_ (.CLK(clknet_leaf_75_clk),
    .D(net895),
    .Q(\mem[8][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4164_ (.CLK(clknet_leaf_53_clk),
    .D(net1295),
    .Q(\mem[8][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4165_ (.CLK(clknet_leaf_43_clk),
    .D(net557),
    .Q(\mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4166_ (.CLK(clknet_leaf_43_clk),
    .D(net607),
    .Q(\mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4167_ (.CLK(clknet_leaf_74_clk),
    .D(net1547),
    .Q(\mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4168_ (.CLK(clknet_leaf_55_clk),
    .D(net737),
    .Q(\mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4169_ (.CLK(clknet_leaf_43_clk),
    .D(net525),
    .Q(\mem[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4170_ (.CLK(clknet_leaf_43_clk),
    .D(net537),
    .Q(\mem[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4171_ (.CLK(clknet_leaf_45_clk),
    .D(net1543),
    .Q(\mem[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4172_ (.CLK(clknet_leaf_67_clk),
    .D(net665),
    .Q(\mem[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4173_ (.CLK(clknet_leaf_54_clk),
    .D(net1027),
    .Q(\mem[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4174_ (.CLK(clknet_leaf_69_clk),
    .D(net1739),
    .Q(\mem[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4175_ (.CLK(clknet_leaf_48_clk),
    .D(net1059),
    .Q(\mem[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4176_ (.CLK(clknet_leaf_71_clk),
    .D(net2291),
    .Q(\mem[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4177_ (.CLK(clknet_leaf_36_clk),
    .D(net713),
    .Q(\mem[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4178_ (.CLK(clknet_leaf_65_clk),
    .D(net1957),
    .Q(\mem[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4179_ (.CLK(clknet_leaf_47_clk),
    .D(net2267),
    .Q(\mem[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4180_ (.CLK(clknet_leaf_62_clk),
    .D(net1157),
    .Q(\mem[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4181_ (.CLK(clknet_leaf_34_clk),
    .D(net1323),
    .Q(\mem[7][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4182_ (.CLK(clknet_leaf_45_clk),
    .D(net1471),
    .Q(\mem[7][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4183_ (.CLK(clknet_leaf_58_clk),
    .D(net1689),
    .Q(\mem[7][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4184_ (.CLK(clknet_leaf_47_clk),
    .D(net1651),
    .Q(\mem[7][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4185_ (.CLK(clknet_leaf_44_clk),
    .D(net1913),
    .Q(\mem[7][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4186_ (.CLK(clknet_leaf_63_clk),
    .D(net1435),
    .Q(\mem[7][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4187_ (.CLK(clknet_leaf_71_clk),
    .D(net2277),
    .Q(\mem[7][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4188_ (.CLK(clknet_leaf_67_clk),
    .D(net1259),
    .Q(\mem[7][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4189_ (.CLK(clknet_leaf_72_clk),
    .D(net1857),
    .Q(\mem[7][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4190_ (.CLK(clknet_leaf_71_clk),
    .D(net1811),
    .Q(\mem[7][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4191_ (.CLK(clknet_leaf_56_clk),
    .D(net2075),
    .Q(\mem[7][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4192_ (.CLK(clknet_leaf_44_clk),
    .D(net1405),
    .Q(\mem[7][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4193_ (.CLK(clknet_leaf_79_clk),
    .D(net1417),
    .Q(\mem[7][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4194_ (.CLK(clknet_leaf_74_clk),
    .D(net1701),
    .Q(\mem[7][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4195_ (.CLK(clknet_leaf_79_clk),
    .D(net921),
    .Q(\mem[7][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4196_ (.CLK(clknet_leaf_53_clk),
    .D(net661),
    .Q(\mem[7][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4197_ (.CLK(clknet_leaf_24_clk),
    .D(net1763),
    .Q(\mem[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4198_ (.CLK(clknet_leaf_25_clk),
    .D(net401),
    .Q(\mem[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4199_ (.CLK(clknet_leaf_92_clk),
    .D(net1089),
    .Q(\mem[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4200_ (.CLK(clknet_leaf_10_clk),
    .D(net2241),
    .Q(\mem[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4201_ (.CLK(clknet_leaf_24_clk),
    .D(net599),
    .Q(\mem[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4202_ (.CLK(clknet_leaf_25_clk),
    .D(net653),
    .Q(\mem[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4203_ (.CLK(clknet_leaf_12_clk),
    .D(net1099),
    .Q(\mem[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4204_ (.CLK(clknet_leaf_0_clk),
    .D(net1573),
    .Q(\mem[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4205_ (.CLK(clknet_leaf_10_clk),
    .D(net2355),
    .Q(\mem[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4206_ (.CLK(clknet_leaf_88_clk),
    .D(net2009),
    .Q(\mem[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4207_ (.CLK(clknet_leaf_15_clk),
    .D(net837),
    .Q(\mem[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4208_ (.CLK(clknet_leaf_86_clk),
    .D(net1757),
    .Q(\mem[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4209_ (.CLK(clknet_leaf_14_clk),
    .D(net711),
    .Q(\mem[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4210_ (.CLK(clknet_leaf_81_clk),
    .D(net1667),
    .Q(\mem[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4211_ (.CLK(clknet_leaf_11_clk),
    .D(net1889),
    .Q(\mem[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4212_ (.CLK(clknet_leaf_6_clk),
    .D(net1005),
    .Q(\mem[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4213_ (.CLK(clknet_leaf_14_clk),
    .D(net1749),
    .Q(\mem[26][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4214_ (.CLK(clknet_leaf_31_clk),
    .D(net1151),
    .Q(\mem[26][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4215_ (.CLK(clknet_leaf_82_clk),
    .D(net1827),
    .Q(\mem[26][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4216_ (.CLK(clknet_leaf_33_clk),
    .D(net937),
    .Q(\mem[26][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4217_ (.CLK(clknet_leaf_20_clk),
    .D(net1945),
    .Q(\mem[26][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4218_ (.CLK(clknet_leaf_7_clk),
    .D(net911),
    .Q(\mem[26][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4219_ (.CLK(clknet_leaf_86_clk),
    .D(net1719),
    .Q(\mem[26][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4220_ (.CLK(clknet_leaf_88_clk),
    .D(net1523),
    .Q(\mem[26][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4221_ (.CLK(clknet_leaf_88_clk),
    .D(net1565),
    .Q(\mem[26][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4222_ (.CLK(clknet_leaf_87_clk),
    .D(net2245),
    .Q(\mem[26][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4223_ (.CLK(clknet_leaf_84_clk),
    .D(net1901),
    .Q(\mem[26][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4224_ (.CLK(clknet_leaf_13_clk),
    .D(net933),
    .Q(\mem[26][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4225_ (.CLK(clknet_leaf_5_clk),
    .D(net1103),
    .Q(\mem[26][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4226_ (.CLK(clknet_leaf_92_clk),
    .D(net1219),
    .Q(\mem[26][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4227_ (.CLK(clknet_leaf_92_clk),
    .D(net1121),
    .Q(\mem[26][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4228_ (.CLK(clknet_leaf_10_clk),
    .D(net1839),
    .Q(\mem[26][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4229_ (.CLK(clknet_leaf_42_clk),
    .D(net495),
    .Q(\mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4230_ (.CLK(clknet_leaf_40_clk),
    .D(net375),
    .Q(\mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4231_ (.CLK(clknet_leaf_74_clk),
    .D(net1283),
    .Q(\mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4232_ (.CLK(clknet_leaf_34_clk),
    .D(net1183),
    .Q(\mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4233_ (.CLK(clknet_leaf_41_clk),
    .D(net387),
    .Q(\mem[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4234_ (.CLK(clknet_leaf_42_clk),
    .D(net781),
    .Q(\mem[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4235_ (.CLK(clknet_leaf_46_clk),
    .D(net1147),
    .Q(\mem[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4236_ (.CLK(clknet_leaf_66_clk),
    .D(net761),
    .Q(\mem[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4237_ (.CLK(clknet_leaf_57_clk),
    .D(net1211),
    .Q(\mem[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4238_ (.CLK(clknet_leaf_66_clk),
    .D(net961),
    .Q(\mem[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4239_ (.CLK(clknet_leaf_49_clk),
    .D(net757),
    .Q(\mem[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4240_ (.CLK(clknet_leaf_71_clk),
    .D(net1979),
    .Q(\mem[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4241_ (.CLK(clknet_leaf_35_clk),
    .D(net845),
    .Q(\mem[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4242_ (.CLK(clknet_leaf_62_clk),
    .D(net1227),
    .Q(\mem[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4243_ (.CLK(clknet_leaf_49_clk),
    .D(net1483),
    .Q(\mem[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4244_ (.CLK(clknet_leaf_61_clk),
    .D(net749),
    .Q(\mem[9][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4245_ (.CLK(clknet_leaf_35_clk),
    .D(net1207),
    .Q(\mem[9][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4246_ (.CLK(clknet_leaf_45_clk),
    .D(net1375),
    .Q(\mem[9][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4247_ (.CLK(clknet_leaf_58_clk),
    .D(net1999),
    .Q(\mem[9][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4248_ (.CLK(clknet_leaf_49_clk),
    .D(net1067),
    .Q(\mem[9][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4249_ (.CLK(clknet_leaf_45_clk),
    .D(net2191),
    .Q(\mem[9][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4250_ (.CLK(clknet_leaf_61_clk),
    .D(net1441),
    .Q(\mem[9][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4251_ (.CLK(clknet_leaf_66_clk),
    .D(net1733),
    .Q(\mem[9][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4252_ (.CLK(clknet_leaf_65_clk),
    .D(net1065),
    .Q(\mem[9][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4253_ (.CLK(clknet_leaf_76_clk),
    .D(net677),
    .Q(\mem[9][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4254_ (.CLK(clknet_leaf_76_clk),
    .D(net1033),
    .Q(\mem[9][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4255_ (.CLK(clknet_leaf_80_clk),
    .D(net1855),
    .Q(\mem[9][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4256_ (.CLK(clknet_leaf_38_clk),
    .D(net835),
    .Q(\mem[9][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4257_ (.CLK(clknet_leaf_80_clk),
    .D(net755),
    .Q(\mem[9][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4258_ (.CLK(clknet_leaf_75_clk),
    .D(net1193),
    .Q(\mem[9][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4259_ (.CLK(clknet_leaf_75_clk),
    .D(net789),
    .Q(\mem[9][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4260_ (.CLK(clknet_leaf_53_clk),
    .D(net1313),
    .Q(\mem[9][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4261_ (.CLK(clknet_leaf_43_clk),
    .D(net575),
    .Q(\mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4262_ (.CLK(clknet_leaf_43_clk),
    .D(net541),
    .Q(\mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4263_ (.CLK(clknet_leaf_73_clk),
    .D(net1445),
    .Q(\mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4264_ (.CLK(clknet_leaf_54_clk),
    .D(net947),
    .Q(\mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4265_ (.CLK(clknet_leaf_43_clk),
    .D(net471),
    .Q(\mem[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4266_ (.CLK(clknet_leaf_43_clk),
    .D(net555),
    .Q(\mem[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4267_ (.CLK(clknet_leaf_46_clk),
    .D(net2173),
    .Q(\mem[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4268_ (.CLK(clknet_leaf_71_clk),
    .D(net2045),
    .Q(\mem[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4269_ (.CLK(clknet_leaf_57_clk),
    .D(net2049),
    .Q(\mem[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4270_ (.CLK(clknet_leaf_70_clk),
    .D(net1389),
    .Q(\mem[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4271_ (.CLK(clknet_leaf_49_clk),
    .D(net1631),
    .Q(\mem[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4272_ (.CLK(clknet_leaf_70_clk),
    .D(net1509),
    .Q(\mem[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4273_ (.CLK(clknet_leaf_36_clk),
    .D(net1037),
    .Q(\mem[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4274_ (.CLK(clknet_leaf_60_clk),
    .D(net1237),
    .Q(\mem[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4275_ (.CLK(clknet_leaf_51_clk),
    .D(net1019),
    .Q(\mem[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4276_ (.CLK(clknet_leaf_61_clk),
    .D(net695),
    .Q(\mem[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4277_ (.CLK(clknet_leaf_37_clk),
    .D(net1847),
    .Q(\mem[12][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4278_ (.CLK(clknet_leaf_46_clk),
    .D(net941),
    .Q(\mem[12][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4279_ (.CLK(clknet_leaf_58_clk),
    .D(net2149),
    .Q(\mem[12][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4280_ (.CLK(clknet_leaf_50_clk),
    .D(net879),
    .Q(\mem[12][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4281_ (.CLK(clknet_leaf_52_clk),
    .D(net1251),
    .Q(\mem[12][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4282_ (.CLK(clknet_leaf_60_clk),
    .D(net1507),
    .Q(\mem[12][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4283_ (.CLK(clknet_leaf_70_clk),
    .D(net1327),
    .Q(\mem[12][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4284_ (.CLK(clknet_leaf_69_clk),
    .D(net1197),
    .Q(\mem[12][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4285_ (.CLK(clknet_leaf_72_clk),
    .D(net2157),
    .Q(\mem[12][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4286_ (.CLK(clknet_leaf_72_clk),
    .D(net2273),
    .Q(\mem[12][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4287_ (.CLK(clknet_leaf_56_clk),
    .D(net1137),
    .Q(\mem[12][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4288_ (.CLK(clknet_leaf_52_clk),
    .D(net1463),
    .Q(\mem[12][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4289_ (.CLK(clknet_leaf_78_clk),
    .D(net609),
    .Q(\mem[12][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4290_ (.CLK(clknet_leaf_72_clk),
    .D(net2067),
    .Q(\mem[12][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4291_ (.CLK(clknet_leaf_72_clk),
    .D(net1381),
    .Q(\mem[12][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4292_ (.CLK(clknet_leaf_52_clk),
    .D(net671),
    .Q(\mem[12][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4293_ (.CLK(clknet_leaf_23_clk),
    .D(net431),
    .Q(\mem[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4294_ (.CLK(clknet_leaf_23_clk),
    .D(net409),
    .Q(\mem[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4295_ (.CLK(clknet_leaf_93_clk),
    .D(net643),
    .Q(\mem[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4296_ (.CLK(clknet_leaf_17_clk),
    .D(net849),
    .Q(\mem[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4297_ (.CLK(clknet_leaf_23_clk),
    .D(net451),
    .Q(\mem[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4298_ (.CLK(clknet_leaf_24_clk),
    .D(net531),
    .Q(\mem[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4299_ (.CLK(clknet_leaf_21_clk),
    .D(net735),
    .Q(\mem[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4300_ (.CLK(clknet_leaf_3_clk),
    .D(net809),
    .Q(\mem[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4301_ (.CLK(clknet_leaf_9_clk),
    .D(net2243),
    .Q(\mem[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4302_ (.CLK(clknet_leaf_90_clk),
    .D(net751),
    .Q(\mem[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4303_ (.CLK(clknet_leaf_16_clk),
    .D(net967),
    .Q(\mem[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4304_ (.CLK(clknet_leaf_8_clk),
    .D(net1795),
    .Q(\mem[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4305_ (.CLK(clknet_leaf_17_clk),
    .D(net1319),
    .Q(\mem[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4306_ (.CLK(clknet_leaf_9_clk),
    .D(net2341),
    .Q(\mem[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4307_ (.CLK(clknet_leaf_18_clk),
    .D(net1473),
    .Q(\mem[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4308_ (.CLK(clknet_leaf_4_clk),
    .D(net1205),
    .Q(\mem[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4309_ (.CLK(clknet_leaf_18_clk),
    .D(net817),
    .Q(\mem[23][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4310_ (.CLK(clknet_leaf_12_clk),
    .D(net2409),
    .Q(\mem[23][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4311_ (.CLK(clknet_leaf_8_clk),
    .D(net1419),
    .Q(\mem[23][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4312_ (.CLK(clknet_leaf_12_clk),
    .D(net801),
    .Q(\mem[23][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4313_ (.CLK(clknet_leaf_20_clk),
    .D(net2297),
    .Q(\mem[23][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4314_ (.CLK(clknet_leaf_1_clk),
    .D(net1261),
    .Q(\mem[23][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4315_ (.CLK(clknet_leaf_84_clk),
    .D(net1249),
    .Q(\mem[23][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4316_ (.CLK(clknet_leaf_8_clk),
    .D(net1723),
    .Q(\mem[23][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4317_ (.CLK(clknet_leaf_93_clk),
    .D(net889),
    .Q(\mem[23][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4318_ (.CLK(clknet_leaf_83_clk),
    .D(net1687),
    .Q(\mem[23][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4319_ (.CLK(clknet_leaf_4_clk),
    .D(net1521),
    .Q(\mem[23][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4320_ (.CLK(clknet_leaf_18_clk),
    .D(net1057),
    .Q(\mem[23][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4321_ (.CLK(clknet_leaf_4_clk),
    .D(net1577),
    .Q(\mem[23][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4322_ (.CLK(clknet_leaf_1_clk),
    .D(net2135),
    .Q(\mem[23][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4323_ (.CLK(clknet_leaf_3_clk),
    .D(net873),
    .Q(\mem[23][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4324_ (.CLK(clknet_leaf_16_clk),
    .D(net719),
    .Q(\mem[23][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4325_ (.CLK(clknet_leaf_26_clk),
    .D(net885),
    .Q(\mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4326_ (.CLK(clknet_leaf_27_clk),
    .D(net427),
    .Q(\mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4327_ (.CLK(clknet_leaf_74_clk),
    .D(net1923),
    .Q(\mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4328_ (.CLK(clknet_leaf_34_clk),
    .D(net649),
    .Q(\mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4329_ (.CLK(clknet_leaf_26_clk),
    .D(net463),
    .Q(\mem[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4330_ (.CLK(clknet_leaf_26_clk),
    .D(net407),
    .Q(\mem[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4331_ (.CLK(clknet_leaf_46_clk),
    .D(net991),
    .Q(\mem[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4332_ (.CLK(clknet_leaf_65_clk),
    .D(net1621),
    .Q(\mem[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4333_ (.CLK(clknet_leaf_56_clk),
    .D(net1123),
    .Q(\mem[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4334_ (.CLK(clknet_leaf_66_clk),
    .D(net1315),
    .Q(\mem[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4335_ (.CLK(clknet_leaf_49_clk),
    .D(net2059),
    .Q(\mem[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4336_ (.CLK(clknet_leaf_71_clk),
    .D(net1915),
    .Q(\mem[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4337_ (.CLK(clknet_leaf_35_clk),
    .D(net1587),
    .Q(\mem[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4338_ (.CLK(clknet_leaf_60_clk),
    .D(net673),
    .Q(\mem[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4339_ (.CLK(clknet_leaf_50_clk),
    .D(net943),
    .Q(\mem[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4340_ (.CLK(clknet_leaf_61_clk),
    .D(net909),
    .Q(\mem[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4341_ (.CLK(clknet_leaf_35_clk),
    .D(net1457),
    .Q(\mem[11][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4342_ (.CLK(clknet_leaf_45_clk),
    .D(net2179),
    .Q(\mem[11][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4343_ (.CLK(clknet_leaf_58_clk),
    .D(net1771),
    .Q(\mem[11][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4344_ (.CLK(clknet_leaf_49_clk),
    .D(net1989),
    .Q(\mem[11][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4345_ (.CLK(clknet_leaf_44_clk),
    .D(net953),
    .Q(\mem[11][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4346_ (.CLK(clknet_leaf_61_clk),
    .D(net1097),
    .Q(\mem[11][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4347_ (.CLK(clknet_leaf_59_clk),
    .D(net1607),
    .Q(\mem[11][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4348_ (.CLK(clknet_leaf_65_clk),
    .D(net2337),
    .Q(\mem[11][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4349_ (.CLK(clknet_leaf_76_clk),
    .D(net907),
    .Q(\mem[11][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4350_ (.CLK(clknet_leaf_76_clk),
    .D(net1107),
    .Q(\mem[11][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4351_ (.CLK(clknet_leaf_80_clk),
    .D(net1173),
    .Q(\mem[11][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4352_ (.CLK(clknet_leaf_38_clk),
    .D(net593),
    .Q(\mem[11][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4353_ (.CLK(clknet_leaf_80_clk),
    .D(net1095),
    .Q(\mem[11][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4354_ (.CLK(clknet_leaf_75_clk),
    .D(net1845),
    .Q(\mem[11][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4355_ (.CLK(clknet_leaf_75_clk),
    .D(net1871),
    .Q(\mem[11][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4356_ (.CLK(clknet_leaf_54_clk),
    .D(net1143),
    .Q(\mem[11][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4357_ (.CLK(clknet_leaf_28_clk),
    .D(net499),
    .Q(\mem[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4358_ (.CLK(clknet_leaf_29_clk),
    .D(net433),
    .Q(\mem[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4359_ (.CLK(clknet_leaf_0_clk),
    .D(net1823),
    .Q(\mem[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4360_ (.CLK(clknet_leaf_4_clk),
    .D(net1305),
    .Q(\mem[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4361_ (.CLK(clknet_leaf_23_clk),
    .D(net435),
    .Q(\mem[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4362_ (.CLK(clknet_leaf_29_clk),
    .D(net515),
    .Q(\mem[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4363_ (.CLK(clknet_leaf_21_clk),
    .D(net799),
    .Q(\mem[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4364_ (.CLK(clknet_leaf_2_clk),
    .D(net1167),
    .Q(\mem[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4365_ (.CLK(clknet_leaf_10_clk),
    .D(net2385),
    .Q(\mem[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4366_ (.CLK(clknet_leaf_89_clk),
    .D(net1829),
    .Q(\mem[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4367_ (.CLK(clknet_leaf_5_clk),
    .D(net2165),
    .Q(\mem[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4368_ (.CLK(clknet_leaf_89_clk),
    .D(net1515),
    .Q(\mem[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4369_ (.CLK(clknet_leaf_16_clk),
    .D(net2317),
    .Q(\mem[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4370_ (.CLK(clknet_leaf_9_clk),
    .D(net2093),
    .Q(\mem[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4371_ (.CLK(clknet_leaf_20_clk),
    .D(net2129),
    .Q(\mem[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4372_ (.CLK(clknet_leaf_5_clk),
    .D(net1239),
    .Q(\mem[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4373_ (.CLK(clknet_leaf_18_clk),
    .D(net1277),
    .Q(\mem[18][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4374_ (.CLK(clknet_leaf_30_clk),
    .D(net699),
    .Q(\mem[18][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4375_ (.CLK(clknet_leaf_83_clk),
    .D(net823),
    .Q(\mem[18][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4376_ (.CLK(clknet_leaf_11_clk),
    .D(net1637),
    .Q(\mem[18][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4377_ (.CLK(clknet_leaf_20_clk),
    .D(net1759),
    .Q(\mem[18][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4378_ (.CLK(clknet_leaf_6_clk),
    .D(net827),
    .Q(\mem[18][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4379_ (.CLK(clknet_leaf_89_clk),
    .D(net1817),
    .Q(\mem[18][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4380_ (.CLK(clknet_leaf_83_clk),
    .D(net1165),
    .Q(\mem[18][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4381_ (.CLK(clknet_leaf_0_clk),
    .D(net2389),
    .Q(\mem[18][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4382_ (.CLK(clknet_leaf_84_clk),
    .D(net2175),
    .Q(\mem[18][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4383_ (.CLK(clknet_leaf_2_clk),
    .D(net2027),
    .Q(\mem[18][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4384_ (.CLK(clknet_leaf_21_clk),
    .D(net1767),
    .Q(\mem[18][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4385_ (.CLK(clknet_leaf_5_clk),
    .D(net1977),
    .Q(\mem[18][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4386_ (.CLK(clknet_leaf_0_clk),
    .D(net2285),
    .Q(\mem[18][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4387_ (.CLK(clknet_leaf_2_clk),
    .D(net1589),
    .Q(\mem[18][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4388_ (.CLK(clknet_leaf_11_clk),
    .D(net2347),
    .Q(\mem[18][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4389_ (.CLK(clknet_leaf_38_clk),
    .D(net383),
    .Q(\mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4390_ (.CLK(clknet_leaf_44_clk),
    .D(net769),
    .Q(\mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4391_ (.CLK(clknet_leaf_76_clk),
    .D(net645),
    .Q(\mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4392_ (.CLK(clknet_leaf_54_clk),
    .D(net1369),
    .Q(\mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4393_ (.CLK(clknet_leaf_38_clk),
    .D(net371),
    .Q(\mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4394_ (.CLK(clknet_leaf_44_clk),
    .D(net563),
    .Q(\mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4395_ (.CLK(clknet_leaf_47_clk),
    .D(net1539),
    .Q(\mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4396_ (.CLK(clknet_leaf_64_clk),
    .D(net1041),
    .Q(\mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4397_ (.CLK(clknet_leaf_57_clk),
    .D(net1925),
    .Q(\mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4398_ (.CLK(clknet_leaf_64_clk),
    .D(net1007),
    .Q(\mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4399_ (.CLK(clknet_leaf_48_clk),
    .D(net1641),
    .Q(\mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4400_ (.CLK(clknet_leaf_66_clk),
    .D(net1495),
    .Q(\mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4401_ (.CLK(clknet_leaf_37_clk),
    .D(net1707),
    .Q(\mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4402_ (.CLK(clknet_leaf_64_clk),
    .D(net831),
    .Q(\mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4403_ (.CLK(clknet_leaf_47_clk),
    .D(net2231),
    .Q(\mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4404_ (.CLK(clknet_leaf_63_clk),
    .D(net979),
    .Q(\mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4405_ (.CLK(clknet_leaf_37_clk),
    .D(net1453),
    .Q(\mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4406_ (.CLK(clknet_leaf_47_clk),
    .D(net1769),
    .Q(\mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4407_ (.CLK(clknet_leaf_59_clk),
    .D(net1217),
    .Q(\mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4408_ (.CLK(clknet_leaf_48_clk),
    .D(net1633),
    .Q(\mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4409_ (.CLK(clknet_leaf_51_clk),
    .D(net1233),
    .Q(\mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4410_ (.CLK(clknet_leaf_63_clk),
    .D(net975),
    .Q(\mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4411_ (.CLK(clknet_leaf_59_clk),
    .D(net2211),
    .Q(\mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4412_ (.CLK(clknet_leaf_64_clk),
    .D(net935),
    .Q(\mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4413_ (.CLK(clknet_leaf_77_clk),
    .D(net1831),
    .Q(\mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4414_ (.CLK(clknet_leaf_58_clk),
    .D(net2147),
    .Q(\mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4415_ (.CLK(clknet_leaf_57_clk),
    .D(net1015),
    .Q(\mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4416_ (.CLK(clknet_leaf_52_clk),
    .D(net1265),
    .Q(\mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4417_ (.CLK(clknet_leaf_58_clk),
    .D(net2031),
    .Q(\mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4418_ (.CLK(clknet_leaf_77_clk),
    .D(net2133),
    .Q(\mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4419_ (.CLK(clknet_leaf_77_clk),
    .D(net923),
    .Q(\mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4420_ (.CLK(clknet_leaf_54_clk),
    .D(net1035),
    .Q(\mem[0][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4421_ (.CLK(clknet_leaf_39_clk),
    .D(net379),
    .Q(\mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4422_ (.CLK(clknet_leaf_39_clk),
    .D(net505),
    .Q(\mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4423_ (.CLK(clknet_leaf_75_clk),
    .D(net2247),
    .Q(\mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4424_ (.CLK(clknet_leaf_54_clk),
    .D(net1401),
    .Q(\mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4425_ (.CLK(clknet_leaf_39_clk),
    .D(net437),
    .Q(\mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4426_ (.CLK(clknet_leaf_39_clk),
    .D(net395),
    .Q(\mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4427_ (.CLK(clknet_leaf_47_clk),
    .D(net1887),
    .Q(\mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4428_ (.CLK(clknet_leaf_64_clk),
    .D(net1609),
    .Q(\mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4429_ (.CLK(clknet_leaf_57_clk),
    .D(net1177),
    .Q(\mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4430_ (.CLK(clknet_leaf_68_clk),
    .D(net585),
    .Q(\mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4431_ (.CLK(clknet_leaf_48_clk),
    .D(net999),
    .Q(\mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4432_ (.CLK(clknet_leaf_77_clk),
    .D(net1199),
    .Q(\mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4433_ (.CLK(clknet_leaf_37_clk),
    .D(net1161),
    .Q(\mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4434_ (.CLK(clknet_leaf_63_clk),
    .D(net785),
    .Q(\mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4435_ (.CLK(clknet_leaf_47_clk),
    .D(net2177),
    .Q(\mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4436_ (.CLK(clknet_leaf_63_clk),
    .D(net1029),
    .Q(\mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4437_ (.CLK(clknet_leaf_53_clk),
    .D(net903),
    .Q(\mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4438_ (.CLK(clknet_leaf_47_clk),
    .D(net2065),
    .Q(\mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4439_ (.CLK(clknet_leaf_59_clk),
    .D(net777),
    .Q(\mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4440_ (.CLK(clknet_leaf_48_clk),
    .D(net1781),
    .Q(\mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4441_ (.CLK(clknet_leaf_51_clk),
    .D(net927),
    .Q(\mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4442_ (.CLK(clknet_leaf_63_clk),
    .D(net1189),
    .Q(\mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4443_ (.CLK(clknet_leaf_59_clk),
    .D(net1373),
    .Q(\mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4444_ (.CLK(clknet_leaf_64_clk),
    .D(net2081),
    .Q(\mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4445_ (.CLK(clknet_leaf_76_clk),
    .D(net1787),
    .Q(\mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4446_ (.CLK(clknet_leaf_58_clk),
    .D(net1359),
    .Q(\mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4447_ (.CLK(clknet_leaf_57_clk),
    .D(net1799),
    .Q(\mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4448_ (.CLK(clknet_leaf_52_clk),
    .D(net989),
    .Q(\mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4449_ (.CLK(clknet_leaf_58_clk),
    .D(net1713),
    .Q(\mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4450_ (.CLK(clknet_leaf_77_clk),
    .D(net773),
    .Q(\mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4451_ (.CLK(clknet_leaf_77_clk),
    .D(net1431),
    .Q(\mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4452_ (.CLK(clknet_leaf_53_clk),
    .D(net1437),
    .Q(\mem[1][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4453_ (.CLK(clknet_leaf_43_clk),
    .D(net1741),
    .Q(\mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4454_ (.CLK(clknet_leaf_43_clk),
    .D(net513),
    .Q(\mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4455_ (.CLK(clknet_leaf_74_clk),
    .D(net1807),
    .Q(\mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4456_ (.CLK(clknet_leaf_55_clk),
    .D(net1229),
    .Q(\mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4457_ (.CLK(clknet_leaf_43_clk),
    .D(net597),
    .Q(\mem[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4458_ (.CLK(clknet_leaf_43_clk),
    .D(net697),
    .Q(\mem[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4459_ (.CLK(clknet_leaf_45_clk),
    .D(net1731),
    .Q(\mem[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4460_ (.CLK(clknet_leaf_67_clk),
    .D(net1735),
    .Q(\mem[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4461_ (.CLK(clknet_leaf_57_clk),
    .D(net1191),
    .Q(\mem[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4462_ (.CLK(clknet_leaf_69_clk),
    .D(net707),
    .Q(\mem[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4463_ (.CLK(clknet_leaf_48_clk),
    .D(net1133),
    .Q(\mem[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4464_ (.CLK(clknet_leaf_71_clk),
    .D(net2057),
    .Q(\mem[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4465_ (.CLK(clknet_leaf_36_clk),
    .D(net1965),
    .Q(\mem[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4466_ (.CLK(clknet_leaf_64_clk),
    .D(net1055),
    .Q(\mem[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4467_ (.CLK(clknet_leaf_47_clk),
    .D(net1907),
    .Q(\mem[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4468_ (.CLK(clknet_leaf_62_clk),
    .D(net1801),
    .Q(\mem[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4469_ (.CLK(clknet_leaf_34_clk),
    .D(net1397),
    .Q(\mem[4][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4470_ (.CLK(clknet_leaf_45_clk),
    .D(net1591),
    .Q(\mem[4][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4471_ (.CLK(clknet_leaf_60_clk),
    .D(net1489),
    .Q(\mem[4][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4472_ (.CLK(clknet_leaf_48_clk),
    .D(net1549),
    .Q(\mem[4][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4473_ (.CLK(clknet_leaf_44_clk),
    .D(net1351),
    .Q(\mem[4][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4474_ (.CLK(clknet_leaf_63_clk),
    .D(net1909),
    .Q(\mem[4][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4475_ (.CLK(clknet_leaf_66_clk),
    .D(net2005),
    .Q(\mem[4][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4476_ (.CLK(clknet_leaf_68_clk),
    .D(net891),
    .Q(\mem[4][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4477_ (.CLK(clknet_leaf_71_clk),
    .D(net2193),
    .Q(\mem[4][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4478_ (.CLK(clknet_leaf_71_clk),
    .D(net2083),
    .Q(\mem[4][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4479_ (.CLK(clknet_leaf_56_clk),
    .D(net1697),
    .Q(\mem[4][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4480_ (.CLK(clknet_leaf_44_clk),
    .D(net1039),
    .Q(\mem[4][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4481_ (.CLK(clknet_leaf_78_clk),
    .D(net1981),
    .Q(\mem[4][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4482_ (.CLK(clknet_leaf_76_clk),
    .D(net1939),
    .Q(\mem[4][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4483_ (.CLK(clknet_leaf_78_clk),
    .D(net1493),
    .Q(\mem[4][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4484_ (.CLK(clknet_leaf_53_clk),
    .D(net717),
    .Q(\mem[4][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4485_ (.CLK(clknet_leaf_22_clk),
    .D(net415),
    .Q(\mem[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4486_ (.CLK(clknet_leaf_29_clk),
    .D(net377),
    .Q(\mem[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4487_ (.CLK(clknet_leaf_0_clk),
    .D(net2053),
    .Q(\mem[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4488_ (.CLK(clknet_leaf_16_clk),
    .D(net1243),
    .Q(\mem[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4489_ (.CLK(clknet_leaf_22_clk),
    .D(net475),
    .Q(\mem[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4490_ (.CLK(clknet_leaf_22_clk),
    .D(net569),
    .Q(\mem[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4491_ (.CLK(clknet_leaf_20_clk),
    .D(net1849),
    .Q(\mem[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4492_ (.CLK(clknet_leaf_1_clk),
    .D(net2207),
    .Q(\mem[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4493_ (.CLK(clknet_leaf_9_clk),
    .D(net2251),
    .Q(\mem[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4494_ (.CLK(clknet_leaf_89_clk),
    .D(net2169),
    .Q(\mem[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4495_ (.CLK(clknet_leaf_5_clk),
    .D(net2289),
    .Q(\mem[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4496_ (.CLK(clknet_leaf_84_clk),
    .D(net2203),
    .Q(\mem[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4497_ (.CLK(clknet_leaf_16_clk),
    .D(net1049),
    .Q(\mem[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4498_ (.CLK(clknet_leaf_10_clk),
    .D(net2097),
    .Q(\mem[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4499_ (.CLK(clknet_leaf_19_clk),
    .D(net765),
    .Q(\mem[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4500_ (.CLK(clknet_leaf_5_clk),
    .D(net1533),
    .Q(\mem[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4501_ (.CLK(clknet_leaf_14_clk),
    .D(net1679),
    .Q(\mem[16][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4502_ (.CLK(clknet_leaf_31_clk),
    .D(net1341),
    .Q(\mem[16][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4503_ (.CLK(clknet_leaf_81_clk),
    .D(net1969),
    .Q(\mem[16][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4504_ (.CLK(clknet_leaf_31_clk),
    .D(net905),
    .Q(\mem[16][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4505_ (.CLK(clknet_leaf_20_clk),
    .D(net2119),
    .Q(\mem[16][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4506_ (.CLK(clknet_leaf_9_clk),
    .D(net2019),
    .Q(\mem[16][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4507_ (.CLK(clknet_leaf_84_clk),
    .D(net1709),
    .Q(\mem[16][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4508_ (.CLK(clknet_leaf_82_clk),
    .D(net1345),
    .Q(\mem[16][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4509_ (.CLK(clknet_leaf_0_clk),
    .D(net1897),
    .Q(\mem[16][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4510_ (.CLK(clknet_leaf_84_clk),
    .D(net1947),
    .Q(\mem[16][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4511_ (.CLK(clknet_leaf_2_clk),
    .D(net1367),
    .Q(\mem[16][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4512_ (.CLK(clknet_leaf_19_clk),
    .D(net1349),
    .Q(\mem[16][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4513_ (.CLK(clknet_leaf_7_clk),
    .D(net1585),
    .Q(\mem[16][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4514_ (.CLK(clknet_leaf_1_clk),
    .D(net1699),
    .Q(\mem[16][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4515_ (.CLK(clknet_leaf_1_clk),
    .D(net1467),
    .Q(\mem[16][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4516_ (.CLK(clknet_leaf_11_clk),
    .D(net1805),
    .Q(\mem[16][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4517_ (.CLK(clknet_leaf_23_clk),
    .D(net493),
    .Q(\mem[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4518_ (.CLK(clknet_leaf_24_clk),
    .D(net457),
    .Q(\mem[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4519_ (.CLK(clknet_leaf_93_clk),
    .D(net825),
    .Q(\mem[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4520_ (.CLK(clknet_leaf_16_clk),
    .D(net1597),
    .Q(\mem[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4521_ (.CLK(clknet_leaf_24_clk),
    .D(net521),
    .Q(\mem[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4522_ (.CLK(clknet_leaf_24_clk),
    .D(net1267),
    .Q(\mem[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4523_ (.CLK(clknet_leaf_19_clk),
    .D(net1053),
    .Q(\mem[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4524_ (.CLK(clknet_leaf_2_clk),
    .D(net915),
    .Q(\mem[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4525_ (.CLK(clknet_leaf_9_clk),
    .D(net2259),
    .Q(\mem[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4526_ (.CLK(clknet_leaf_89_clk),
    .D(net2319),
    .Q(\mem[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4527_ (.CLK(clknet_leaf_15_clk),
    .D(net1567),
    .Q(\mem[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4528_ (.CLK(clknet_leaf_83_clk),
    .D(net1859),
    .Q(\mem[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4529_ (.CLK(clknet_leaf_16_clk),
    .D(net1187),
    .Q(\mem[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4530_ (.CLK(clknet_leaf_9_clk),
    .D(net2209),
    .Q(\mem[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4531_ (.CLK(clknet_leaf_18_clk),
    .D(net1343),
    .Q(\mem[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4532_ (.CLK(clknet_leaf_4_clk),
    .D(net949),
    .Q(\mem[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4533_ (.CLK(clknet_leaf_17_clk),
    .D(net925),
    .Q(\mem[20][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4534_ (.CLK(clknet_leaf_31_clk),
    .D(net1427),
    .Q(\mem[20][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4535_ (.CLK(clknet_leaf_9_clk),
    .D(net2269),
    .Q(\mem[20][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4536_ (.CLK(clknet_leaf_12_clk),
    .D(net887),
    .Q(\mem[20][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4537_ (.CLK(clknet_leaf_20_clk),
    .D(net2017),
    .Q(\mem[20][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4538_ (.CLK(clknet_leaf_7_clk),
    .D(net1433),
    .Q(\mem[20][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4539_ (.CLK(clknet_leaf_84_clk),
    .D(net2025),
    .Q(\mem[20][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4540_ (.CLK(clknet_leaf_83_clk),
    .D(net1869),
    .Q(\mem[20][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4541_ (.CLK(clknet_leaf_0_clk),
    .D(net2323),
    .Q(\mem[20][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4542_ (.CLK(clknet_leaf_82_clk),
    .D(net847),
    .Q(\mem[20][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4543_ (.CLK(clknet_leaf_3_clk),
    .D(net955),
    .Q(\mem[20][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4544_ (.CLK(clknet_leaf_19_clk),
    .D(net1949),
    .Q(\mem[20][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4545_ (.CLK(clknet_leaf_4_clk),
    .D(net1163),
    .Q(\mem[20][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4546_ (.CLK(clknet_leaf_1_clk),
    .D(net1309),
    .Q(\mem[20][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4547_ (.CLK(clknet_leaf_2_clk),
    .D(net657),
    .Q(\mem[20][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4548_ (.CLK(clknet_leaf_15_clk),
    .D(net659),
    .Q(\mem[20][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4549_ (.CLK(clknet_leaf_41_clk),
    .D(net545),
    .Q(\mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4550_ (.CLK(clknet_leaf_41_clk),
    .D(net439),
    .Q(\mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4551_ (.CLK(clknet_leaf_74_clk),
    .D(net997),
    .Q(\mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4552_ (.CLK(clknet_leaf_34_clk),
    .D(net865),
    .Q(\mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4553_ (.CLK(clknet_leaf_26_clk),
    .D(net553),
    .Q(\mem[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4554_ (.CLK(clknet_leaf_26_clk),
    .D(net519),
    .Q(\mem[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4555_ (.CLK(clknet_leaf_46_clk),
    .D(net1563),
    .Q(\mem[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4556_ (.CLK(clknet_leaf_66_clk),
    .D(net779),
    .Q(\mem[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4557_ (.CLK(clknet_leaf_56_clk),
    .D(net1765),
    .Q(\mem[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4558_ (.CLK(clknet_leaf_66_clk),
    .D(net1047),
    .Q(\mem[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4559_ (.CLK(clknet_leaf_49_clk),
    .D(net1329),
    .Q(\mem[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4560_ (.CLK(clknet_leaf_71_clk),
    .D(net2011),
    .Q(\mem[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4561_ (.CLK(clknet_leaf_32_clk),
    .D(net1425),
    .Q(\mem[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4562_ (.CLK(clknet_leaf_59_clk),
    .D(net1605),
    .Q(\mem[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4563_ (.CLK(clknet_leaf_51_clk),
    .D(net977),
    .Q(\mem[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4564_ (.CLK(clknet_leaf_61_clk),
    .D(net1379),
    .Q(\mem[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4565_ (.CLK(clknet_leaf_35_clk),
    .D(net721),
    .Q(\mem[10][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4566_ (.CLK(clknet_leaf_45_clk),
    .D(net1105),
    .Q(\mem[10][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4567_ (.CLK(clknet_leaf_58_clk),
    .D(net1289),
    .Q(\mem[10][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4568_ (.CLK(clknet_leaf_50_clk),
    .D(net1171),
    .Q(\mem[10][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4569_ (.CLK(clknet_leaf_44_clk),
    .D(net1705),
    .Q(\mem[10][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4570_ (.CLK(clknet_leaf_61_clk),
    .D(net1085),
    .Q(\mem[10][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4571_ (.CLK(clknet_leaf_59_clk),
    .D(net1669),
    .Q(\mem[10][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4572_ (.CLK(clknet_leaf_65_clk),
    .D(net1791),
    .Q(\mem[10][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4573_ (.CLK(clknet_leaf_76_clk),
    .D(net1339),
    .Q(\mem[10][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4574_ (.CLK(clknet_leaf_76_clk),
    .D(net2141),
    .Q(\mem[10][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4575_ (.CLK(clknet_leaf_80_clk),
    .D(net1145),
    .Q(\mem[10][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4576_ (.CLK(clknet_leaf_38_clk),
    .D(net945),
    .Q(\mem[10][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4577_ (.CLK(clknet_leaf_80_clk),
    .D(net669),
    .Q(\mem[10][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4578_ (.CLK(clknet_leaf_74_clk),
    .D(net1061),
    .Q(\mem[10][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4579_ (.CLK(clknet_leaf_75_clk),
    .D(net1083),
    .Q(\mem[10][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4580_ (.CLK(clknet_leaf_54_clk),
    .D(net1231),
    .Q(\mem[10][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4581_ (.CLK(clknet_leaf_42_clk),
    .D(net547),
    .Q(\mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4582_ (.CLK(clknet_leaf_41_clk),
    .D(net473),
    .Q(\mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4583_ (.CLK(clknet_leaf_73_clk),
    .D(net1929),
    .Q(\mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4584_ (.CLK(clknet_leaf_55_clk),
    .D(net833),
    .Q(\mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4585_ (.CLK(clknet_leaf_41_clk),
    .D(net489),
    .Q(\mem[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4586_ (.CLK(clknet_leaf_42_clk),
    .D(net441),
    .Q(\mem[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4587_ (.CLK(clknet_leaf_51_clk),
    .D(net1635),
    .Q(\mem[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4588_ (.CLK(clknet_leaf_71_clk),
    .D(net2261),
    .Q(\mem[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4589_ (.CLK(clknet_leaf_57_clk),
    .D(net1201),
    .Q(\mem[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4590_ (.CLK(clknet_leaf_70_clk),
    .D(net1777),
    .Q(\mem[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4591_ (.CLK(clknet_leaf_50_clk),
    .D(net1087),
    .Q(\mem[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4592_ (.CLK(clknet_leaf_72_clk),
    .D(net1783),
    .Q(\mem[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4593_ (.CLK(clknet_leaf_35_clk),
    .D(net1203),
    .Q(\mem[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4594_ (.CLK(clknet_leaf_59_clk),
    .D(net1109),
    .Q(\mem[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4595_ (.CLK(clknet_leaf_51_clk),
    .D(net1529),
    .Q(\mem[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4596_ (.CLK(clknet_leaf_60_clk),
    .D(net703),
    .Q(\mem[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4597_ (.CLK(clknet_leaf_35_clk),
    .D(net995),
    .Q(\mem[14][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4598_ (.CLK(clknet_leaf_46_clk),
    .D(net1253),
    .Q(\mem[14][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4599_ (.CLK(clknet_leaf_77_clk),
    .D(net965),
    .Q(\mem[14][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4600_ (.CLK(clknet_leaf_50_clk),
    .D(net621),
    .Q(\mem[14][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4601_ (.CLK(clknet_leaf_52_clk),
    .D(net1517),
    .Q(\mem[14][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4602_ (.CLK(clknet_leaf_60_clk),
    .D(net1715),
    .Q(\mem[14][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4603_ (.CLK(clknet_leaf_70_clk),
    .D(net1497),
    .Q(\mem[14][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4604_ (.CLK(clknet_leaf_70_clk),
    .D(net1575),
    .Q(\mem[14][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4605_ (.CLK(clknet_leaf_72_clk),
    .D(net1919),
    .Q(\mem[14][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4606_ (.CLK(clknet_leaf_72_clk),
    .D(net2103),
    .Q(\mem[14][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4607_ (.CLK(clknet_leaf_80_clk),
    .D(net725),
    .Q(\mem[14][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4608_ (.CLK(clknet_leaf_37_clk),
    .D(net1023),
    .Q(\mem[14][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4609_ (.CLK(clknet_leaf_79_clk),
    .D(net629),
    .Q(\mem[14][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4610_ (.CLK(clknet_leaf_73_clk),
    .D(net813),
    .Q(\mem[14][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4611_ (.CLK(clknet_leaf_73_clk),
    .D(net705),
    .Q(\mem[14][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4612_ (.CLK(clknet_leaf_52_clk),
    .D(net1843),
    .Q(\mem[14][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4613_ (.CLK(clknet_leaf_42_clk),
    .D(net429),
    .Q(\mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4614_ (.CLK(clknet_leaf_41_clk),
    .D(net399),
    .Q(\mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4615_ (.CLK(clknet_leaf_73_clk),
    .D(net1075),
    .Q(\mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4616_ (.CLK(clknet_leaf_55_clk),
    .D(net797),
    .Q(\mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4617_ (.CLK(clknet_leaf_42_clk),
    .D(net419),
    .Q(\mem[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4618_ (.CLK(clknet_leaf_42_clk),
    .D(net393),
    .Q(\mem[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4619_ (.CLK(clknet_leaf_46_clk),
    .D(net1671),
    .Q(\mem[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4620_ (.CLK(clknet_leaf_71_clk),
    .D(net1785),
    .Q(\mem[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4621_ (.CLK(clknet_leaf_54_clk),
    .D(net1045),
    .Q(\mem[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4622_ (.CLK(clknet_leaf_70_clk),
    .D(net1593),
    .Q(\mem[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4623_ (.CLK(clknet_leaf_50_clk),
    .D(net763),
    .Q(\mem[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4624_ (.CLK(clknet_leaf_70_clk),
    .D(net1245),
    .Q(\mem[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4625_ (.CLK(clknet_leaf_36_clk),
    .D(net689),
    .Q(\mem[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4626_ (.CLK(clknet_leaf_59_clk),
    .D(net839),
    .Q(\mem[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4627_ (.CLK(clknet_leaf_51_clk),
    .D(net1399),
    .Q(\mem[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4628_ (.CLK(clknet_leaf_61_clk),
    .D(net775),
    .Q(\mem[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4629_ (.CLK(clknet_leaf_35_clk),
    .D(net1063),
    .Q(\mem[13][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4630_ (.CLK(clknet_leaf_46_clk),
    .D(net815),
    .Q(\mem[13][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4631_ (.CLK(clknet_leaf_58_clk),
    .D(net1113),
    .Q(\mem[13][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4632_ (.CLK(clknet_leaf_50_clk),
    .D(net1127),
    .Q(\mem[13][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4633_ (.CLK(clknet_leaf_52_clk),
    .D(net1629),
    .Q(\mem[13][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4634_ (.CLK(clknet_leaf_60_clk),
    .D(net1255),
    .Q(\mem[13][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4635_ (.CLK(clknet_leaf_70_clk),
    .D(net1125),
    .Q(\mem[13][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4636_ (.CLK(clknet_leaf_69_clk),
    .D(net963),
    .Q(\mem[13][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4637_ (.CLK(clknet_leaf_72_clk),
    .D(net2021),
    .Q(\mem[13][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4638_ (.CLK(clknet_leaf_72_clk),
    .D(net1893),
    .Q(\mem[13][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4639_ (.CLK(clknet_leaf_56_clk),
    .D(net1301),
    .Q(\mem[13][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4640_ (.CLK(clknet_leaf_37_clk),
    .D(net981),
    .Q(\mem[13][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4641_ (.CLK(clknet_leaf_80_clk),
    .D(net931),
    .Q(\mem[13][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4642_ (.CLK(clknet_leaf_73_clk),
    .D(net791),
    .Q(\mem[13][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4643_ (.CLK(clknet_leaf_72_clk),
    .D(net1761),
    .Q(\mem[13][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4644_ (.CLK(clknet_leaf_53_clk),
    .D(net863),
    .Q(\mem[13][31] ));
 sky130_fd_sc_hd__dfxtp_1 _4645_ (.CLK(clknet_leaf_43_clk),
    .D(net539),
    .Q(\mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _4646_ (.CLK(clknet_leaf_44_clk),
    .D(net571),
    .Q(\mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _4647_ (.CLK(clknet_leaf_74_clk),
    .D(net1819),
    .Q(\mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _4648_ (.CLK(clknet_leaf_55_clk),
    .D(net1093),
    .Q(\mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _4649_ (.CLK(clknet_leaf_43_clk),
    .D(net549),
    .Q(\mem[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _4650_ (.CLK(clknet_leaf_43_clk),
    .D(net601),
    .Q(\mem[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _4651_ (.CLK(clknet_leaf_45_clk),
    .D(net1185),
    .Q(\mem[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _4652_ (.CLK(clknet_leaf_67_clk),
    .D(net2105),
    .Q(\mem[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _4653_ (.CLK(clknet_leaf_54_clk),
    .D(net1335),
    .Q(\mem[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _4654_ (.CLK(clknet_leaf_69_clk),
    .D(net871),
    .Q(\mem[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _4655_ (.CLK(clknet_leaf_48_clk),
    .D(net1481),
    .Q(\mem[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _4656_ (.CLK(clknet_leaf_71_clk),
    .D(net2223),
    .Q(\mem[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _4657_ (.CLK(clknet_leaf_36_clk),
    .D(net841),
    .Q(\mem[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _4658_ (.CLK(clknet_leaf_65_clk),
    .D(net1421),
    .Q(\mem[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _4659_ (.CLK(clknet_leaf_47_clk),
    .D(net1511),
    .Q(\mem[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _4660_ (.CLK(clknet_leaf_62_clk),
    .D(net2125),
    .Q(\mem[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _4661_ (.CLK(clknet_leaf_34_clk),
    .D(net743),
    .Q(\mem[5][16] ));
 sky130_fd_sc_hd__dfxtp_1 _4662_ (.CLK(clknet_leaf_45_clk),
    .D(net1209),
    .Q(\mem[5][17] ));
 sky130_fd_sc_hd__dfxtp_1 _4663_ (.CLK(clknet_leaf_58_clk),
    .D(net1403),
    .Q(\mem[5][18] ));
 sky130_fd_sc_hd__dfxtp_1 _4664_ (.CLK(clknet_leaf_48_clk),
    .D(net1281),
    .Q(\mem[5][19] ));
 sky130_fd_sc_hd__dfxtp_1 _4665_ (.CLK(clknet_leaf_44_clk),
    .D(net1413),
    .Q(\mem[5][20] ));
 sky130_fd_sc_hd__dfxtp_1 _4666_ (.CLK(clknet_leaf_62_clk),
    .D(net1755),
    .Q(\mem[5][21] ));
 sky130_fd_sc_hd__dfxtp_1 _4667_ (.CLK(clknet_leaf_66_clk),
    .D(net731),
    .Q(\mem[5][22] ));
 sky130_fd_sc_hd__dfxtp_1 _4668_ (.CLK(clknet_leaf_68_clk),
    .D(net507),
    .Q(\mem[5][23] ));
 sky130_fd_sc_hd__dfxtp_1 _4669_ (.CLK(clknet_leaf_71_clk),
    .D(net2411),
    .Q(\mem[5][24] ));
 sky130_fd_sc_hd__dfxtp_1 _4670_ (.CLK(clknet_leaf_72_clk),
    .D(net1729),
    .Q(\mem[5][25] ));
 sky130_fd_sc_hd__dfxtp_1 _4671_ (.CLK(clknet_leaf_56_clk),
    .D(net1837),
    .Q(\mem[5][26] ));
 sky130_fd_sc_hd__dfxtp_1 _4672_ (.CLK(clknet_leaf_44_clk),
    .D(net2229),
    .Q(\mem[5][27] ));
 sky130_fd_sc_hd__dfxtp_1 _4673_ (.CLK(clknet_leaf_79_clk),
    .D(net595),
    .Q(\mem[5][28] ));
 sky130_fd_sc_hd__dfxtp_1 _4674_ (.CLK(clknet_leaf_74_clk),
    .D(net811),
    .Q(\mem[5][29] ));
 sky130_fd_sc_hd__dfxtp_1 _4675_ (.CLK(clknet_leaf_78_clk),
    .D(net855),
    .Q(\mem[5][30] ));
 sky130_fd_sc_hd__dfxtp_1 _4676_ (.CLK(clknet_leaf_51_clk),
    .D(net2363),
    .Q(\mem[5][31] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__buf_6 fanout100 (.A(_1784_),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_8 fanout101 (.A(_1784_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_8 fanout102 (.A(_1780_),
    .X(net102));
 sky130_fd_sc_hd__buf_4 fanout103 (.A(_1780_),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_8 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_8 fanout105 (.A(_1776_),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(_1772_),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(_1772_),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_8 fanout108 (.A(net109),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_8 fanout109 (.A(_1768_),
    .X(net109));
 sky130_fd_sc_hd__buf_6 fanout110 (.A(net111),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 fanout111 (.A(_1764_),
    .X(net111));
 sky130_fd_sc_hd__buf_6 fanout112 (.A(_1760_),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(_1760_),
    .X(net113));
 sky130_fd_sc_hd__buf_6 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_8 fanout115 (.A(_1756_),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(_1752_),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(_1752_),
    .X(net117));
 sky130_fd_sc_hd__buf_6 fanout118 (.A(_1748_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_8 fanout119 (.A(_1748_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_8 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_8 fanout121 (.A(_1744_),
    .X(net121));
 sky130_fd_sc_hd__buf_6 fanout122 (.A(_1739_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(_1739_),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(_1735_),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_8 fanout125 (.A(_1735_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(_1730_),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_8 fanout128 (.A(_1726_),
    .X(net128));
 sky130_fd_sc_hd__buf_4 fanout129 (.A(_1726_),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_8 fanout131 (.A(_1722_),
    .X(net131));
 sky130_fd_sc_hd__buf_6 fanout132 (.A(_1718_),
    .X(net132));
 sky130_fd_sc_hd__buf_4 fanout133 (.A(_1718_),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 fanout134 (.A(net135),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_8 fanout135 (.A(_1714_),
    .X(net135));
 sky130_fd_sc_hd__buf_6 fanout136 (.A(_1709_),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(_1709_),
    .X(net137));
 sky130_fd_sc_hd__buf_6 fanout138 (.A(_1705_),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(_1705_),
    .X(net139));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(_1701_),
    .X(net140));
 sky130_fd_sc_hd__buf_4 fanout141 (.A(_1701_),
    .X(net141));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(_1697_),
    .X(net142));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(_1697_),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(_1690_),
    .X(net144));
 sky130_fd_sc_hd__buf_4 fanout145 (.A(_1690_),
    .X(net145));
 sky130_fd_sc_hd__buf_6 fanout146 (.A(_1684_),
    .X(net146));
 sky130_fd_sc_hd__buf_4 fanout147 (.A(_1684_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_8 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_8 fanout149 (.A(_1679_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_8 fanout150 (.A(_1673_),
    .X(net150));
 sky130_fd_sc_hd__buf_4 fanout151 (.A(_1673_),
    .X(net151));
 sky130_fd_sc_hd__buf_6 fanout152 (.A(_1806_),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_8 fanout153 (.A(_1806_),
    .X(net153));
 sky130_fd_sc_hd__buf_6 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(_1802_),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_8 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__buf_8 fanout157 (.A(_1798_),
    .X(net157));
 sky130_fd_sc_hd__buf_6 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_6 fanout159 (.A(_1794_),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_8 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_8 fanout161 (.A(_1790_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_8 fanout163 (.A(_1786_),
    .X(net163));
 sky130_fd_sc_hd__buf_6 fanout164 (.A(_1782_),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_8 fanout165 (.A(_1782_),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_8 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_6 fanout167 (.A(_1778_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_8 fanout169 (.A(_1774_),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_8 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_8 fanout171 (.A(_1770_),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_8 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_6 fanout173 (.A(_1766_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_8 fanout175 (.A(_1762_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__buf_6 fanout177 (.A(_1758_),
    .X(net177));
 sky130_fd_sc_hd__buf_6 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_6 fanout179 (.A(_1754_),
    .X(net179));
 sky130_fd_sc_hd__buf_6 fanout180 (.A(_1750_),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_8 fanout181 (.A(_1750_),
    .X(net181));
 sky130_fd_sc_hd__buf_8 fanout182 (.A(_1746_),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(_1746_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__buf_6 fanout185 (.A(_1742_),
    .X(net185));
 sky130_fd_sc_hd__buf_6 fanout186 (.A(_1737_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_8 fanout187 (.A(_1737_),
    .X(net187));
 sky130_fd_sc_hd__buf_6 fanout188 (.A(_1733_),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(_1733_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_8 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(_1728_),
    .X(net191));
 sky130_fd_sc_hd__buf_6 fanout192 (.A(_1724_),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_8 fanout193 (.A(_1724_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(_1720_),
    .X(net195));
 sky130_fd_sc_hd__buf_6 fanout196 (.A(_1716_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_8 fanout197 (.A(_1716_),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_8 fanout199 (.A(_1712_),
    .X(net199));
 sky130_fd_sc_hd__buf_6 fanout200 (.A(_1707_),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(_1707_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_6 fanout203 (.A(_1703_),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_8 fanout204 (.A(_1699_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(_1699_),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_8 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_6 fanout207 (.A(_1695_),
    .X(net207));
 sky130_fd_sc_hd__buf_6 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__buf_6 fanout209 (.A(_1688_),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_8 fanout210 (.A(_1682_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(_1682_),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__buf_6 fanout213 (.A(_1677_),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_8 fanout215 (.A(_1671_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 fanout216 (.A(_1669_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_4 fanout217 (.A(_1669_),
    .X(net217));
 sky130_fd_sc_hd__buf_12 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_12 fanout219 (.A(_1026_),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(net222),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_8 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(_1025_),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(_1025_),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_4 fanout224 (.A(_1025_),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net9),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net9),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_8 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_8 fanout228 (.A(net8),
    .X(net228));
 sky130_fd_sc_hd__buf_8 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_16 fanout230 (.A(net6),
    .X(net230));
 sky130_fd_sc_hd__buf_8 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_8 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(net6),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_8 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_6 fanout235 (.A(net240),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(net237),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_8 fanout237 (.A(net240),
    .X(net237));
 sky130_fd_sc_hd__buf_8 fanout238 (.A(net240),
    .X(net238));
 sky130_fd_sc_hd__buf_8 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_8 fanout240 (.A(net5),
    .X(net240));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net4),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net4),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_8 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_8 fanout244 (.A(net4),
    .X(net244));
 sky130_fd_sc_hd__buf_8 fanout245 (.A(net248),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net248),
    .X(net246));
 sky130_fd_sc_hd__buf_8 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__buf_8 fanout248 (.A(net4),
    .X(net248));
 sky130_fd_sc_hd__buf_4 fanout249 (.A(net39),
    .X(net249));
 sky130_fd_sc_hd__buf_4 fanout250 (.A(net39),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net38),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(net38),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(net37),
    .X(net253));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(net37),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net36),
    .X(net255));
 sky130_fd_sc_hd__buf_4 fanout256 (.A(net36),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_8 fanout257 (.A(net35),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net35),
    .X(net258));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_8 fanout260 (.A(net34),
    .X(net260));
 sky130_fd_sc_hd__buf_4 fanout261 (.A(net263),
    .X(net261));
 sky130_fd_sc_hd__buf_2 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_4 fanout263 (.A(net33),
    .X(net263));
 sky130_fd_sc_hd__buf_4 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_8 fanout265 (.A(net32),
    .X(net265));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(net31),
    .X(net266));
 sky130_fd_sc_hd__buf_4 fanout267 (.A(net31),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(net30),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(net30),
    .X(net269));
 sky130_fd_sc_hd__buf_4 fanout270 (.A(net273),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net273),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(net285),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net285),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(net285),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net285),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net285),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(net280),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(net285),
    .X(net280));
 sky130_fd_sc_hd__buf_4 fanout281 (.A(net285),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 fanout282 (.A(net285),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(net285),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_4 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(net3),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_8 fanout286 (.A(net290),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_8 fanout287 (.A(net290),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_8 fanout288 (.A(net289),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_8 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net3),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_8 fanout291 (.A(net294),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_8 fanout292 (.A(net294),
    .X(net292));
 sky130_fd_sc_hd__buf_2 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_4 fanout294 (.A(net3),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_8 fanout295 (.A(net296),
    .X(net295));
 sky130_fd_sc_hd__buf_4 fanout296 (.A(net3),
    .X(net296));
 sky130_fd_sc_hd__buf_4 fanout297 (.A(net29),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(net29),
    .X(net298));
 sky130_fd_sc_hd__buf_4 fanout299 (.A(net28),
    .X(net299));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(net28),
    .X(net300));
 sky130_fd_sc_hd__buf_4 fanout301 (.A(net27),
    .X(net301));
 sky130_fd_sc_hd__buf_4 fanout302 (.A(net27),
    .X(net302));
 sky130_fd_sc_hd__buf_4 fanout303 (.A(net304),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 fanout305 (.A(net26),
    .X(net305));
 sky130_fd_sc_hd__buf_4 fanout306 (.A(net25),
    .X(net306));
 sky130_fd_sc_hd__buf_4 fanout307 (.A(net25),
    .X(net307));
 sky130_fd_sc_hd__buf_4 fanout308 (.A(net24),
    .X(net308));
 sky130_fd_sc_hd__buf_4 fanout309 (.A(net24),
    .X(net309));
 sky130_fd_sc_hd__buf_4 fanout310 (.A(net23),
    .X(net310));
 sky130_fd_sc_hd__buf_4 fanout311 (.A(net23),
    .X(net311));
 sky130_fd_sc_hd__buf_4 fanout312 (.A(net22),
    .X(net312));
 sky130_fd_sc_hd__buf_4 fanout313 (.A(net22),
    .X(net313));
 sky130_fd_sc_hd__buf_4 fanout314 (.A(net21),
    .X(net314));
 sky130_fd_sc_hd__buf_4 fanout315 (.A(net21),
    .X(net315));
 sky130_fd_sc_hd__buf_4 fanout316 (.A(net20),
    .X(net316));
 sky130_fd_sc_hd__buf_4 fanout317 (.A(net20),
    .X(net317));
 sky130_fd_sc_hd__buf_6 fanout318 (.A(net321),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_8 fanout319 (.A(net321),
    .X(net319));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(net333),
    .X(net321));
 sky130_fd_sc_hd__buf_6 fanout322 (.A(net333),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(net333),
    .X(net323));
 sky130_fd_sc_hd__buf_6 fanout324 (.A(net333),
    .X(net324));
 sky130_fd_sc_hd__buf_4 fanout325 (.A(net333),
    .X(net325));
 sky130_fd_sc_hd__buf_6 fanout326 (.A(net328),
    .X(net326));
 sky130_fd_sc_hd__buf_4 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__buf_4 fanout328 (.A(net333),
    .X(net328));
 sky130_fd_sc_hd__buf_6 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_8 fanout330 (.A(net333),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_8 fanout331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_8 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(net2),
    .X(net333));
 sky130_fd_sc_hd__buf_6 fanout334 (.A(net338),
    .X(net334));
 sky130_fd_sc_hd__buf_6 fanout335 (.A(net338),
    .X(net335));
 sky130_fd_sc_hd__buf_6 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_8 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_6 fanout338 (.A(net2),
    .X(net338));
 sky130_fd_sc_hd__buf_6 fanout339 (.A(net342),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_8 fanout340 (.A(net342),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 fanout342 (.A(net2),
    .X(net342));
 sky130_fd_sc_hd__buf_8 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__buf_4 fanout344 (.A(net2),
    .X(net344));
 sky130_fd_sc_hd__buf_4 fanout345 (.A(net19),
    .X(net345));
 sky130_fd_sc_hd__buf_4 fanout346 (.A(net19),
    .X(net346));
 sky130_fd_sc_hd__buf_4 fanout347 (.A(net18),
    .X(net347));
 sky130_fd_sc_hd__buf_4 fanout348 (.A(net18),
    .X(net348));
 sky130_fd_sc_hd__buf_4 fanout349 (.A(net17),
    .X(net349));
 sky130_fd_sc_hd__buf_4 fanout350 (.A(net17),
    .X(net350));
 sky130_fd_sc_hd__buf_4 fanout351 (.A(net16),
    .X(net351));
 sky130_fd_sc_hd__buf_4 fanout352 (.A(net16),
    .X(net352));
 sky130_fd_sc_hd__buf_4 fanout353 (.A(net15),
    .X(net353));
 sky130_fd_sc_hd__buf_4 fanout354 (.A(net15),
    .X(net354));
 sky130_fd_sc_hd__buf_4 fanout355 (.A(net14),
    .X(net355));
 sky130_fd_sc_hd__buf_4 fanout356 (.A(net14),
    .X(net356));
 sky130_fd_sc_hd__buf_4 fanout357 (.A(net13),
    .X(net357));
 sky130_fd_sc_hd__buf_4 fanout358 (.A(net13),
    .X(net358));
 sky130_fd_sc_hd__buf_4 fanout359 (.A(net12),
    .X(net359));
 sky130_fd_sc_hd__buf_4 fanout360 (.A(net12),
    .X(net360));
 sky130_fd_sc_hd__buf_4 fanout361 (.A(net11),
    .X(net361));
 sky130_fd_sc_hd__buf_4 fanout362 (.A(net11),
    .X(net362));
 sky130_fd_sc_hd__buf_4 fanout363 (.A(net10),
    .X(net363));
 sky130_fd_sc_hd__buf_4 fanout364 (.A(net10),
    .X(net364));
 sky130_fd_sc_hd__buf_4 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_4 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__buf_4 fanout367 (.A(net1),
    .X(net367));
 sky130_fd_sc_hd__buf_4 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_4 fanout369 (.A(net1),
    .X(net369));
 sky130_fd_sc_hd__buf_8 fanout88 (.A(_1808_),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_8 fanout89 (.A(_1808_),
    .X(net89));
 sky130_fd_sc_hd__buf_6 fanout90 (.A(_1804_),
    .X(net90));
 sky130_fd_sc_hd__buf_4 fanout91 (.A(_1804_),
    .X(net91));
 sky130_fd_sc_hd__buf_6 fanout92 (.A(_1800_),
    .X(net92));
 sky130_fd_sc_hd__buf_4 fanout93 (.A(_1800_),
    .X(net93));
 sky130_fd_sc_hd__buf_6 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_8 fanout95 (.A(_1796_),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_8 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_8 fanout97 (.A(_1792_),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_8 fanout98 (.A(net99),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_8 fanout99 (.A(_1788_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\mem[0][4] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_0285_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_0611_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(_0256_),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\mem[28][12] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(_0842_),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\mem[1][22] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(_0307_),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\mem[9][17] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(_0110_),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\mem[30][20] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(_0626_),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\mem[10][15] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\mem[12][4] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(_0428_),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\mem[12][30] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(_0155_),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\mem[28][6] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(_0836_),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\mem[27][11] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(_0777_),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\mem[29][12] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(_1002_),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\mem[12][9] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_0129_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(_0134_),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\mem[3][25] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(_0823_),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\mem[24][14] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(_0684_),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\mem[25][12] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(_0746_),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\mem[4][16] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(_0333_),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\mem[13][14] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\mem[14][1] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(_0491_),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\mem[1][3] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(_0288_),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\mem[5][18] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(_0527_),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\mem[7][27] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(_0056_),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\mem[6][3] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(_0961_),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\mem[27][20] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_0446_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(_0786_),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\mem[15][24] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(_0662_),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\mem[5][20] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(_0529_),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\mem[25][9] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(_0743_),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\mem[7][28] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(_0057_),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\mem[23][18] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\mem[16][4] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(_0175_),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\mem[5][13] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(_0522_),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\mem[6][15] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(_0973_),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\mem[10][12] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(_0425_),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\mem[20][17] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(_0398_),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\mem[21][6] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_0353_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(_0547_),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\mem[1][30] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(_0315_),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\mem[20][21] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(_0402_),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\mem[7][21] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(_0050_),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\mem[1][31] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(_0316_),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\mem[17][26] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\mem[21][0] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(_0952_),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\mem[9][21] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(_0114_),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\mem[2][23] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(_0885_),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\mem[12][2] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(_0127_),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\mem[17][28] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(_0954_),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\mem[30][21] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_0541_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(_0627_),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\mem[21][14] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(_0555_),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\mem[0][16] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(_0269_),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\mem[30][11] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(_0617_),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\mem[11][16] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(_0205_),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\mem[29][26] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\mem[17][1] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(_1016_),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\mem[22][7] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(_0581_),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\mem[12][27] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(_0152_),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\mem[28][19] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(_0849_),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\mem[16][30] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(_0379_),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\mem[3][18] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\mem[27][1] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_0927_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(_0816_),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\mem[7][17] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(_0046_),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\mem[23][14] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(_0171_),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\mem[17][17] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(_0943_),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\mem[2][17] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(_0879_),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\mem[29][30] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\mem[15][0] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(_1020_),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\mem[5][10] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(_0519_),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\mem[9][14] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(_0107_),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\mem[6][23] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(_0981_),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\mem[3][13] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(_0811_),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\mem[4][18] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_0638_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(_0335_),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\mem[2][20] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(_0882_),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\mem[4][30] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(_0347_),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\mem[0][11] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(_0264_),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\mem[14][22] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(_0467_),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\mem[22][17] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\mem[19][0] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(_0591_),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\mem[2][27] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(_0889_),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\mem[21][30] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(_0571_),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\mem[24][8] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(_0678_),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\mem[12][21] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(_0146_),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\mem[12][11] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_0894_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(_0136_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\mem[5][14] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(_0523_),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\mem[28][23] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(_0853_),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\mem[18][11] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(_0232_),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\mem[14][20] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(_0465_),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\mem[15][29] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\mem[24][4] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(_0667_),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\mem[23][26] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(_0183_),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\mem[26][23] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(_0084_),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\mem[22][27] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(_0601_),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\mem[28][10] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(_0840_),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\mem[14][14] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(_0674_),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(_0459_),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\mem[2][6] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(_0868_),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\mem[16][15] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(_0364_),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\mem[19][28] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(_0922_),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\mem[28][24] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(_0854_),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\mem[0][6] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\mem[8][1] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(_0259_),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\mem[25][20] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(_0754_),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\mem[7][6] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(_0035_),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\mem[27][21] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(_0787_),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\mem[7][2] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(_0031_),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\mem[4][19] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_1023_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(_0336_),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\mem[31][22] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(_0724_),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\mem[17][11] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(_0937_),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\mem[8][12] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(_0009_),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\mem[28][30] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(_0860_),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\mem[21][25] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\mem[14][4] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(_0566_),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\mem[30][30] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(_0636_),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\mem[10][6] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(_0419_),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\mem[26][24] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(_0085_),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\mem[20][10] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(_0391_),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\mem[24][2] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_0767_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_0449_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(_0672_),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\mem[19][6] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(_0900_),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\mem[26][7] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(_0068_),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\mem[14][23] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(_0468_),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\mem[23][28] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(_0185_),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\mem[27][22] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\mem[31][5] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(_0788_),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\mem[8][20] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(_0017_),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\mem[22][31] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(_0605_),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\mem[16][28] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(_0377_),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\mem[11][12] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(_0201_),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\mem[18][30] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_0707_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(_0251_),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\mem[4][17] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(_0334_),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\mem[13][9] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(_0486_),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\mem[31][6] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(_0708_),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\mem[20][3] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(_0384_),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\mem[22][18] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\mem[20][0] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(_0592_),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\mem[28][11] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(_0841_),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\mem[22][15] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(_0589_),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\mem[10][13] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(_0426_),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\mem[11][22] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(_0211_),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\mem[1][7] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_0381_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(_0292_),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\mem[29][11] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(_1001_),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\mem[19][17] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(_0911_),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\mem[3][30] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(_0828_),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\mem[19][10] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(_0904_),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\mem[15][16] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\mem[9][0] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(_0654_),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\mem[11][7] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(_0196_),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\mem[6][30] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(_0988_),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\mem[2][18] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(_0880_),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\mem[22][9] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(_0583_),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\mem[13][20] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_0093_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(_0497_),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\mem[12][10] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(_0135_),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\mem[0][19] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(_0272_),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\mem[14][6] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(_0451_),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\mem[18][19] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(_0240_),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\mem[21][11] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\mem[24][1] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(_0552_),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\mem[0][10] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(_0263_),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\mem[24][24] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(_0694_),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\mem[3][8] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(_0806_),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\mem[15][7] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(_0645_),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\mem[27][25] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_0671_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(_0791_),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\mem[7][19] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(_0048_),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\mem[30][9] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(_0615_),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\mem[15][9] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(_0647_),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\mem[31][7] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(_0709_),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\mem[3][6] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\mem[18][0] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(_0804_),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\mem[21][12] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(_0553_),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\mem[3][19] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(_0817_),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\mem[21][19] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(_0560_),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\mem[26][13] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(_0074_),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\mem[10][22] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\mem[0][0] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_0221_),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(_0435_),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\mem[13][6] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(_0483_),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\mem[29][10] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(_1000_),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\mem[24][19] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(_0689_),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\mem[29][25] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(_1015_),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\mem[16][16] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\mem[8][4] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(_0365_),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\mem[17][12] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(_0938_),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\mem[30][27] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(_0633_),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\mem[6][11] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(_0969_),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\mem[23][25] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(_0182_),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\mem[7][18] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_0001_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(_0047_),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\mem[30][18] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(_0624_),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\mem[31][25] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(_0727_),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\mem[3][7] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(_0805_),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\mem[4][26] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(_0343_),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\mem[16][29] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\mem[19][1] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(_0378_),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\mem[7][29] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(_0058_),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\mem[31][19] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(_0721_),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\mem[10][20] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(_0433_),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\mem[0][12] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(_0265_),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\mem[16][22] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_0895_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(_0371_),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\mem[24][26] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(_0696_),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\mem[1][28] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(_0313_),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\mem[14][21] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(_0466_),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\mem[19][30] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(_0924_),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\mem[26][22] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\mem[1][1] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(_0083_),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\mem[2][31] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(_0893_),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\mem[23][23] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(_0180_),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\mem[27][17] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(_0783_),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\mem[2][30] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(_0892_),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\mem[5][25] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_0286_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(_0534_),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\mem[4][6] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(_0323_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\mem[9][22] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(_0115_),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\mem[4][7] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(_0324_),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\mem[19][29] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(_0923_),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\mem[7][9] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\mem[5][23] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(_0038_),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\mem[4][0] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(_0317_),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\mem[22][12] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(_0586_),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\mem[2][10] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(_0872_),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\mem[22][22] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(_0596_),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\mem[26][16] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_0532_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(_0077_),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\mem[6][10] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(_0968_),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\mem[3][17] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(_0815_),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\mem[5][21] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(_0530_),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\mem[26][11] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(_0072_),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\mem[18][20] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\mem[29][0] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(_0241_),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\mem[13][30] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(_0507_),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\mem[26][0] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(_0061_),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\mem[10][8] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(_0421_),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\mem[18][27] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(_0248_),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\mem[0][17] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0253_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_0990_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(_0270_),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\mem[11][18] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(_0207_),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\mem[30][22] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(_0628_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\mem[31][21] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(_0723_),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\mem[14][9] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(_0454_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\mem[31][23] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\mem[2][0] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(_0725_),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\mem[1][19] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(_0304_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\mem[14][11] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(_0456_),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\mem[13][7] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(_0484_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\mem[1][24] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(_0309_),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\mem[29][27] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_0862_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(_1017_),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\mem[10][23] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(_0436_),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(\mem[8][27] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(_0024_),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\mem[23][11] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(_0168_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\mem[30][16] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(_0622_),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\mem[1][26] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\mem[4][1] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(_0311_),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\mem[4][15] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(_0332_),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\mem[22][26] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(_0600_),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\mem[16][31] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(_0380_),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\mem[4][2] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(_0319_),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\mem[17][22] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_0318_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(_0948_),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\mem[7][25] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(_0054_),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(\mem[19][21] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(_0915_),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\mem[17][29] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(_0955_),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\mem[18][22] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(_0243_),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\mem[5][2] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\mem[18][5] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(_0511_),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\mem[29][23] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(_1013_),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\mem[18][2] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(_0223_),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\mem[31][10] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(_0712_),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\mem[26][18] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(_0079_),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\mem[18][9] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_0226_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(_0230_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\mem[0][24] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(_0277_),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\mem[2][14] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(_0876_),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\mem[8][10] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(_0007_),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\mem[5][26] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(_0535_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(\mem[26][31] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\mem[6][4] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(_0092_),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\mem[3][2] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(_0800_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\mem[14][31] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(_0476_),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\mem[11][29] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(_0218_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\mem[12][16] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(_0141_),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\mem[16][6] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_0962_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(_0355_),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\mem[28][16] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(_0846_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\mem[27][8] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(_0774_),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\mem[9][26] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(_0119_),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\mem[7][24] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(_0053_),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\mem[20][11] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\mem[10][5] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(_0392_),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\mem[24][13] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(_0683_),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\mem[29][16] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(_1006_),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\mem[25][24] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(_0758_),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\mem[21][18] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(_0559_),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(\mem[20][23] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\mem[8][5] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(_0418_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(_0404_),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\mem[11][30] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(_0219_),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(\mem[22][29] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(_0603_),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\mem[22][3] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(_0577_),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(\mem[8][18] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(_0015_),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\mem[17][6] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\mem[20][4] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(_0932_),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\mem[29][2] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(_0992_),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\mem[19][8] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(_0902_),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\mem[28][27] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(_0857_),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\mem[1][6] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(_0291_),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\mem[26][14] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_0385_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(_0075_),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(\mem[8][26] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(_0023_),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\mem[13][25] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(_0502_),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\mem[2][22] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(_0884_),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\mem[16][24] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(_0373_),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\mem[3][27] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\mem[8][0] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(_0825_),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\mem[26][26] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(_0087_),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\mem[2][25] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(_0887_),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(\mem[2][7] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(_0869_),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\mem[4][14] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(_0331_),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(\mem[4][21] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_1022_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(_0338_),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(\mem[3][28] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(_0826_),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\mem[7][20] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(_0049_),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\mem[11][11] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(_0200_),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\mem[8][23] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(_0020_),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(\mem[14][24] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\mem[7][4] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(_0469_),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\mem[31][31] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(_0733_),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\mem[11][2] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(_0191_),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\mem[0][8] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(_0261_),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\mem[17][16] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(_0942_),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\mem[14][2] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_0033_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(_0447_),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\mem[22][14] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(_0588_),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\mem[29][29] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(_1019_),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\mem[17][14] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(_0940_),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\mem[25][29] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(_0763_),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\mem[4][29] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\mem[17][4] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(_0346_),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\mem[28][26] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(_0856_),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\mem[25][18] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(_0752_),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\mem[26][20] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(_0081_),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\mem[16][25] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(_0374_),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\mem[20][27] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_0930_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(_0408_),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\mem[24][11] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(_0681_),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\mem[3][23] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(_0821_),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(\mem[22][20] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(_0594_),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\mem[7][13] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(_0042_),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\mem[29][7] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\mem[21][5] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(_0997_),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\mem[6][6] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(_0964_),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\mem[19][16] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(_0910_),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\mem[4][12] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(_0329_),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\mem[17][30] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(_0956_),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\mem[16][18] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_0002_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_0546_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(_0367_),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\mem[30][13] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(_0619_),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\mem[24][29] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(_0699_),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\mem[27][3] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(_0769_),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(\mem[18][28] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(_0249_),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\mem[9][11] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\mem[23][5] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(_0104_),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\mem[4][28] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(_0345_),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\mem[29][17] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(_1007_),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(\mem[28][14] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(_0844_),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\mem[31][29] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(_0731_),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\mem[11][19] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_0162_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(_0208_),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\mem[8][6] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(_0003_),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\mem[27][18] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(_0784_),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\mem[31][11] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(_0713_),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(\mem[3][20] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(_0818_),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(\mem[9][18] ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\mem[27][0] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(_0111_),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\mem[30][24] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(_0630_),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\mem[24][9] ),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(_0679_),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\mem[4][22] ),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(_0339_),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(\mem[21][22] ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(_0563_),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\mem[26][9] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_0766_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(_0070_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(\mem[10][11] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(_0424_),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\mem[28][13] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(_0843_),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\mem[27][14] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(_0780_),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\mem[20][20] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(_0401_),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(\mem[16][21] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\mem[24][5] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(_0370_),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\mem[13][24] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(_0501_),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\mem[15][15] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(_0653_),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\mem[20][22] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(_0403_),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\mem[18][26] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(_0247_),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\mem[6][22] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_0675_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(_0980_),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\mem[0][28] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(_0281_),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\mem[31][9] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(_0711_),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\mem[28][20] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(_0850_),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\mem[25][28] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(_0762_),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\mem[17][9] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\mem[7][5] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(_0935_),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\mem[28][25] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(_0855_),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\mem[25][27] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(_0761_),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\mem[12][7] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(_0132_),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\mem[6][20] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(_0978_),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\mem[12][8] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_0034_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(_0133_),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\mem[24][12] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(_0682_),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\mem[16][2] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(_0351_),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(\mem[25][8] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(_0742_),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\mem[4][11] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(_0328_),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\mem[11][10] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\mem[5][0] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(_0199_),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\mem[30][28] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(_0634_),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\mem[8][25] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(_0022_),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\mem[1][17] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(_0302_),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\mem[12][29] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(_0154_),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\mem[28][22] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\mem[9][4] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_0509_),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(_0852_),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\mem[2][26] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(_0888_),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\mem[17][19] ),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(_0945_),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\mem[7][26] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(_0055_),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\mem[29][19] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(_1009_),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\mem[30][3] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\mem[12][1] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(_0609_),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\mem[1][23] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(_0308_),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\mem[4][25] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(_0342_),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\mem[3][24] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(_0822_),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\mem[21][15] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(_0556_),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\mem[27][24] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_0126_),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(_0790_),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\mem[17][10] ),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(_0936_),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\mem[18][13] ),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(_0234_),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\mem[22][19] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(_0593_),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\mem[16][13] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(_0362_),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\mem[28][7] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\mem[24][0] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(_0837_),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\mem[31][26] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(_0728_),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\mem[14][25] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(_0470_),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(\mem[5][7] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(_0516_),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\mem[24][25] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(_0695_),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\mem[25][13] ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_0670_),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(_0747_),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(\mem[22][25] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(_0599_),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\mem[3][14] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(_0812_),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(\mem[28][9] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(_0839_),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(\mem[21][24] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(_0565_),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\mem[16][20] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\mem[10][0] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(_0369_),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\mem[3][22] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(_0820_),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\mem[19][22] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(_0916_),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\mem[5][15] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(_0524_),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\mem[31][12] ),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(_0714_),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(\mem[18][14] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_0413_),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(_0235_),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\mem[17][24] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(_0950_),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(\mem[0][29] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(_0282_),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\mem[23][29] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(_0186_),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\mem[15][18] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(_0656_),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(\mem[30][12] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\mem[14][0] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(_0618_),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\mem[10][25] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(_0438_),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\mem[29][9] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(_0999_),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\mem[6][29] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(_0987_),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\mem[0][25] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(_0278_),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\mem[12][18] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_0445_),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(_0143_),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\mem[31][18] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(_0720_),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\mem[27][31] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(_0797_),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\mem[17][2] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(_0928_),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\mem[12][24] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(_0149_),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\mem[29][18] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\mem[5][4] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(_1008_),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\mem[31][28] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(_0730_),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\mem[3][31] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(_0829_),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(\mem[18][10] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(_0231_),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\mem[25][16] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(_0750_),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\mem[16][9] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_0097_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_0513_),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(_0358_),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\mem[6][26] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(_0984_),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(\mem[12][6] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(_0131_),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\mem[18][25] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(_0246_),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\mem[1][14] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(_0299_),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\mem[11][17] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\mem[2][5] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(_0206_),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\mem[22][13] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(_0587_),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\mem[8][8] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(_0005_),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\mem[17][18] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(_0944_),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(\mem[31][24] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(_0726_),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(\mem[17][15] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(_0867_),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(_0941_),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(\mem[9][20] ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(_0113_),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\mem[4][24] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(_0341_),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\mem[8][29] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(_0026_),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(\mem[8][16] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(_0013_),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(\mem[22][28] ),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\mem[10][4] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(_0602_),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(\mem[19][23] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(_0917_),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(\mem[16][11] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(_0360_),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(\mem[24][3] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(_0673_),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\mem[16][7] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(_0356_),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\mem[20][13] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_0417_),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(_0394_),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\mem[0][22] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(_0275_),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\mem[28][29] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(_0859_),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(\mem[29][28] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(_1018_),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(\mem[19][18] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(_0912_),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\mem[25][3] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\mem[12][5] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(_0737_),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(\mem[21][16] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(_0557_),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(\mem[5][11] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(_0520_),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(\mem[25][14] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(_0748_),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(\mem[29][3] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(_0993_),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(\mem[5][27] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_0130_),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(_0536_),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(\mem[0][14] ),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(_0267_),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(\mem[27][26] ),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(_0792_),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(\mem[19][14] ),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(_0908_),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(\mem[17][3] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(_0929_),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(\mem[29][20] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\mem[7][0] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(_1010_),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(\mem[26][3] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(_0064_),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(\mem[23][8] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(_0165_),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(\mem[26][25] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(_0086_),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(\mem[1][2] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(_0287_),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(\mem[22][21] ),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_0029_),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(_0595_),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\mem[16][8] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(_0357_),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(\mem[31][17] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(_0719_),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(\mem[15][14] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(_0652_),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(\mem[2][19] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(_0881_),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(\mem[20][8] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\mem[28][0] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(_0389_),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(\mem[14][7] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(_0452_),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(\mem[8][13] ),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(_0010_),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(\mem[28][18] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(_0848_),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(\mem[7][14] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(_0043_),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(\mem[20][18] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\mem[21][1] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_0830_),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(_0399_),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(\mem[28][21] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(_0851_),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(\mem[12][25] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(_0150_),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(\mem[17][20] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(_0946_),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(\mem[7][22] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(_0051_),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(\mem[30][15] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\mem[28][5] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(_0621_),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(\mem[24][18] ),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(_0688_),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(\mem[6][14] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(_0972_),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(\mem[18][29] ),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(_0250_),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(\mem[15][22] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(_0660_),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(\mem[16][10] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_0835_),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(_0359_),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(\mem[7][11] ),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(_0040_),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(\mem[17][7] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(_0933_),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(\mem[19][7] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(_0901_),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(\mem[23][20] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(_0177_),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(\mem[28][15] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\mem[0][5] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(_0845_),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(\mem[29][21] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(_1011_),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(\mem[19][3] ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(_0897_),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(\mem[22][8] ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(_0582_),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(\mem[19][19] ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(_0913_),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(\mem[31][8] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_0258_),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(_0710_),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(\mem[8][7] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(_0004_),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(\mem[6][24] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(_0982_),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(\mem[29][6] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(_0996_),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(\mem[18][12] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(_0233_),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(\mem[20][9] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\mem[28][4] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(_0390_),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(\mem[24][15] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(_0685_),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(\mem[20][24] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(_0405_),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(\mem[15][11] ),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(_0649_),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(\mem[21][20] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(_0561_),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(\mem[31][15] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_0834_),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(_0717_),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(\mem[27][13] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(_0779_),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(\mem[29][15] ),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(_1005_),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(\mem[29][24] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(_1014_),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(\mem[11][23] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(_0212_),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(\mem[19][31] ),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\mem[22][0] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(_0925_),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(\mem[23][13] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(_0170_),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(\mem[31][13] ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(_0715_),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(\mem[8][24] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(_0021_),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(\mem[18][31] ),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(_0252_),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(\mem[29][13] ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_0574_),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(_1003_),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(\mem[31][20] ),
    .X(net2350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(_0722_),
    .X(net2351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(\mem[30][8] ),
    .X(net2352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(_0614_),
    .X(net2353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(\mem[26][8] ),
    .X(net2354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(_0069_),
    .X(net2355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(\mem[28][8] ),
    .X(net2356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(_0838_),
    .X(net2357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(\mem[6][18] ),
    .X(net2358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\mem[16][5] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(_0976_),
    .X(net2359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(\mem[29][14] ),
    .X(net2360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(_1004_),
    .X(net2361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(\mem[5][31] ),
    .X(net2362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(_0540_),
    .X(net2363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(\mem[29][31] ),
    .X(net2364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(_1021_),
    .X(net2365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(\mem[6][25] ),
    .X(net2366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(_0983_),
    .X(net2367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(\mem[19][15] ),
    .X(net2368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0257_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_0542_),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(_0354_),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(_0909_),
    .X(net2369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(\mem[31][14] ),
    .X(net2370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(_0716_),
    .X(net2371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(\mem[17][31] ),
    .X(net2372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(_0957_),
    .X(net2373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(\mem[8][11] ),
    .X(net2374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(_0008_),
    .X(net2375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(\mem[19][13] ),
    .X(net2376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(_0907_),
    .X(net2377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(\mem[19][9] ),
    .X(net2378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\mem[5][1] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(_0903_),
    .X(net2379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(\mem[31][3] ),
    .X(net2380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(_0705_),
    .X(net2381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(\mem[19][25] ),
    .X(net2382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(_0919_),
    .X(net2383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(\mem[18][8] ),
    .X(net2384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(_0229_),
    .X(net2385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(\mem[31][30] ),
    .X(net2386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(_0732_),
    .X(net2387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(\mem[18][24] ),
    .X(net2388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_0510_),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(_0245_),
    .X(net2389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(\mem[17][25] ),
    .X(net2390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(_0951_),
    .X(net2391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(\mem[19][11] ),
    .X(net2392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(_0905_),
    .X(net2393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(\mem[21][8] ),
    .X(net2394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(_0549_),
    .X(net2395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(\mem[21][13] ),
    .X(net2396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(_0554_),
    .X(net2397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(\mem[17][13] ),
    .X(net2398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\mem[19][4] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(_0939_),
    .X(net2399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(\mem[17][8] ),
    .X(net2400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(_0934_),
    .X(net2401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(\mem[19][20] ),
    .X(net2402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(_0914_),
    .X(net2403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(\mem[31][2] ),
    .X(net2404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(_0704_),
    .X(net2405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(\mem[28][3] ),
    .X(net2406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(_0833_),
    .X(net2407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(\mem[23][17] ),
    .X(net2408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_0898_),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(_0174_),
    .X(net2409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(\mem[5][24] ),
    .X(net2410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(_0533_),
    .X(net2411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(\mem[19][2] ),
    .X(net2412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(_0896_),
    .X(net2413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(\mem[17][21] ),
    .X(net2414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(_0947_),
    .X(net2415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(\mem[29][8] ),
    .X(net2416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(_0998_),
    .X(net2417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\mem[12][0] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_0125_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\mem[27][5] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_0771_),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\mem[31][4] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\mem[2][1] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_0706_),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\mem[6][1] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_0959_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\mem[29][4] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_0994_),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\mem[1][9] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_0294_),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\mem[22][4] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_0578_),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\mem[24][20] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0863_),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_0690_),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\mem[2][4] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_0866_),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\mem[11][27] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_0216_),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\mem[5][28] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_0537_),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\mem[4][4] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_0321_),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\mem[26][4] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\mem[13][5] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_0065_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\mem[5][5] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_0514_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\mem[17][5] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_0931_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\mem[6][5] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_0963_),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\mem[7][1] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_0030_),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\mem[12][28] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_0482_),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_0153_),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\mem[30][31] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_0637_),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\mem[2][9] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_0871_),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\mem[21][10] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(_0551_),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\mem[6][12] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_0970_),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\mem[21][2] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\mem[1][5] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_0543_),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\mem[14][19] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_0464_),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\mem[24][30] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_0700_),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\mem[27][10] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_0776_),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\mem[15][5] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_0643_),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\mem[14][28] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_0290_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_0473_),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\mem[15][27] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_0665_),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\mem[27][27] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_0793_),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\mem[2][2] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_0864_),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\mem[31][1] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_0703_),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\mem[25][22] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\mem[25][1] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_0756_),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\mem[24][23] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_0693_),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\mem[23][2] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_0159_),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\mem[0][2] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_0255_),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\mem[22][24] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_0598_),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\mem[11][3] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0735_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_0192_),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\mem[24][6] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_0676_),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\mem[26][5] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_0066_),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\mem[2][12] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_0874_),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\mem[20][30] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_0411_),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\mem[20][31] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\mem[13][1] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_0412_),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\mem[7][31] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_0060_),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\mem[27][30] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(_0796_),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\mem[7][7] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(_0036_),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\mem[27][29] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(_0795_),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\mem[10][28] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\mem[3][1] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_0478_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_0441_),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\mem[12][31] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(_0156_),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\mem[11][13] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_0202_),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\mem[6][16] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_0974_),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\mem[9][24] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(_0117_),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\mem[21][27] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\mem[26][1] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_0568_),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\mem[30][23] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(_0629_),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\mem[8][3] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(_0000_),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\mem[6][7] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(_0965_),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\mem[25][19] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(_0753_),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\mem[13][12] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_0062_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_0489_),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\mem[28][2] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(_0832_),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\mem[3][3] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(_0801_),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\mem[12][15] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(_0140_),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\mem[4][5] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(_0322_),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\mem[18][17] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\mem[25][5] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_0238_),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\mem[25][21] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(_0755_),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\mem[14][15] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(_0460_),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\mem[14][30] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(_0475_),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\mem[4][9] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(_0326_),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\mem[30][2] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_0739_),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(_0608_),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\mem[26][12] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(_0073_),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\mem[7][12] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(_0041_),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\mem[27][16] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(_0782_),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\mem[4][31] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(_0348_),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\mem[23][31] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\mem[27][4] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(_0188_),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\mem[10][16] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_0429_),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\mem[3][16] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(_0814_),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\mem[14][26] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(_0471_),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\mem[29][5] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(_0995_),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\mem[2][8] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_0770_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(_0870_),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\mem[5][22] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(_0531_),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\mem[30][6] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(_0612_),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\mem[23][6] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(_0163_),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\mem[7][3] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(_0032_),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\mem[6][28] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\mem[11][5] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(_0986_),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\mem[6][27] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(_0985_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\mem[5][16] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(_0525_),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\mem[15][13] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(_0651_),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\mem[6][8] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(_0966_),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\mem[9][15] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_0194_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(_0108_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\mem[23][9] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(_0166_),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\mem[30][26] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(_0632_),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\mem[9][28] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(_0121_),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\mem[9][10] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(_0103_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\mem[3][9] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\mem[23][1] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(_0807_),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\mem[9][7] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(_0100_),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\mem[13][10] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(_0487_),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\mem[16][14] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(_0363_),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\mem[21][17] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(_0558_),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\mem[0][1] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_0799_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_0158_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(_0254_),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\mem[3][21] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(_0819_),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\mem[1][29] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(_0314_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\mem[13][15] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(_0492_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\mem[1][18] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(_0303_),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\mem[10][7] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\mem[3][0] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0420_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\mem[9][5] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(_0098_),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\mem[8][9] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(_0006_),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\mem[1][13] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(_0298_),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\mem[6][31] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(_0989_),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\mem[9][30] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_0798_),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(_0123_),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\mem[13][29] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(_0506_),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\mem[28][28] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(_0858_),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\mem[25][2] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(_0736_),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\mem[13][3] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(_0480_),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\mem[18][6] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\mem[25][4] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(_0227_),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\mem[23][19] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(_0176_),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\mem[2][21] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(_0883_),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\mem[24][27] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(_0697_),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\mem[27][6] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(_0772_),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\mem[23][7] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_0738_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(_0164_),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\mem[5][29] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(_0538_),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\mem[14][29] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(_0474_),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\mem[13][17] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(_0494_),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\mem[23][16] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(_0173_),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\mem[29][22] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\mem[16][0] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(_1012_),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\mem[2][16] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(_0878_),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\mem[18][18] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(_0239_),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\mem[20][2] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(_0383_),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\mem[18][21] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(_0242_),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\mem[15][23] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_0349_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(_0661_),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\mem[0][13] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(_0266_),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\mem[14][3] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(_0448_),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\mem[9][27] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(_0120_),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\mem[26][10] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(_0071_),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\mem[13][13] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\mem[30][4] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(_0490_),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\mem[5][12] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(_0521_),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\mem[21][29] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(_0570_),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\mem[9][12] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(_0105_),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\mem[20][25] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(_0406_),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\mem[23][3] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_0610_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(_0160_),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\mem[15][20] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(_0658_),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\mem[22][6] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(_0580_),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\mem[5][30] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(_0539_),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\mem[22][2] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(_0576_),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\mem[21][26] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\mem[13][4] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(_0567_),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\mem[3][10] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(_0808_),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\mem[13][31] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(_0508_),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\mem[10][3] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(_0416_),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\mem[19][27] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(_0921_),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\mem[3][11] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\mem[9][1] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_0481_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(_0809_),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\mem[5][9] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(_0518_),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\mem[23][30] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(_0187_),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\mem[21][3] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(_0544_),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\mem[8][19] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(_0016_),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\mem[12][19] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\mem[15][1] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(_0144_),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\mem[6][0] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(_0958_),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\mem[24][10] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(_0680_),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\mem[11][0] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(_0189_),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\mem[20][19] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(_0400_),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\mem[23][24] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_0639_),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(_0181_),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\mem[4][23] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(_0340_),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\mem[27][15] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(_0781_),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\mem[8][30] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(_0027_),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\mem[22][5] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(_0579_),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\mem[17][27] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\mem[15][4] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(_0953_),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\mem[22][30] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(_0604_),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\mem[1][16] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(_0301_),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\mem[16][19] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(_0368_),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\mem[11][24] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(_0213_),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\mem[11][15] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_0642_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(_0204_),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\mem[26][21] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(_0082_),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\mem[21][28] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(_0569_),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\mem[20][7] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(_0388_),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\mem[27][2] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(_0768_),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\mem[15][17] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\mem[25][0] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(_0655_),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\mem[7][30] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(_0059_),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\mem[0][30] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(_0283_),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\mem[20][16] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(_0397_),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\mem[1][20] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(_0305_),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\mem[25][17] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_0734_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(_0751_),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\mem[13][28] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(_0505_),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\mem[26][27] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(_0088_),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\mem[0][23] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(_0276_),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\mem[26][19] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(_0080_),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\mem[21][21] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\mem[11][1] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(_0562_),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\mem[12][17] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(_0142_),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\mem[11][14] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(_0203_),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\mem[10][27] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(_0440_),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\mem[12][3] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(_0128_),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\mem[20][15] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_0190_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(_0396_),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\mem[8][17] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(_0014_),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\mem[11][20] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(_0209_),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\mem[20][26] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(_0407_),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\mem[25][6] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(_0740_),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\mem[2][28] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\mem[13][0] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(_0890_),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\mem[9][9] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(_0102_),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\mem[13][23] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(_0500_),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\mem[14][18] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(_0463_),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\mem[23][10] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(_0167_),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\mem[30][29] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0094_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_0477_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(_0635_),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\mem[6][2] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(_0960_),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\mem[19][24] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(_0918_),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\mem[0][21] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(_0274_),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\mem[10][14] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(_0427_),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\mem[0][15] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\mem[23][0] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(_0268_),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\mem[13][27] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(_0504_),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\mem[24][21] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(_0691_),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\mem[21][23] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(_0564_),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\mem[2][3] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(_0865_),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\mem[1][27] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(_0157_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(_0312_),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\mem[11][6] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(_0195_),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\mem[15][30] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(_0668_),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\mem[14][16] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(_0461_),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\mem[10][2] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(_0415_),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\mem[1][10] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\mem[18][1] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(_0295_),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\mem[15][31] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(_0669_),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\mem[8][15] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(_0012_),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\mem[26][15] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(_0076_),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\mem[0][9] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(_0262_),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\mem[6][9] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(_0222_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(_0967_),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\mem[25][25] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(_0759_),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\mem[3][15] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_0813_),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\mem[0][26] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(_0279_),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\mem[2][29] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(_0891_),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\mem[12][14] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\mem[18][4] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(_0139_),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\mem[30][17] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(_0623_),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\mem[14][27] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(_0472_),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\mem[27][19] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(_0785_),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\mem[7][8] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(_0037_),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\mem[1][15] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_0225_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(_0300_),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\mem[8][14] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(_0011_),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\mem[9][25] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(_0118_),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\mem[0][31] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(_0284_),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\mem[12][12] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(_0137_),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\mem[4][27] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\mem[1][4] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(_0344_),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\mem[0][7] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(_0260_),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\mem[30][19] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(_0625_),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\mem[13][8] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(_0485_),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\mem[10][9] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(_0422_),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\mem[16][12] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_0289_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(_0361_),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\mem[19][26] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(_0920_),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\mem[20][6] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(_0387_),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\mem[4][13] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(_0330_),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\mem[23][27] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(_0184_),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\mem[7][10] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\mem[10][1] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(_0039_),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\mem[10][29] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(_0442_),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\mem[13][16] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(_0493_),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\mem[9][23] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(_0116_),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\mem[9][19] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(_0112_),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\mem[6][19] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\mem[16][1] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(_0414_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(_0977_),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\mem[19][12] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(_0906_),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\mem[21][31] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(_0572_),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\mem[13][2] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(_0479_),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\mem[17][0] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(_0926_),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\mem[25][23] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\mem[14][5] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(_0757_),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\mem[25][15] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(_0749_),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\mem[10][30] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(_0443_),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\mem[10][21] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(_0434_),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\mem[14][10] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(_0455_),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\mem[26][2] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_0450_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(_0063_),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\mem[25][11] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(_0745_),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\mem[5][3] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(_0512_),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\mem[11][28] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(_0217_),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\mem[11][21] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(_0210_),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\mem[26][6] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\mem[22][1] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(_0067_),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\mem[3][12] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(_0810_),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\mem[26][28] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(_0089_),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\mem[10][17] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(_0430_),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\mem[11][25] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(_0214_),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\mem[14][13] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_0575_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(_0458_),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\mem[3][26] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(_0824_),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\mem[13][18] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(_0495_),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\mem[2][13] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(_0875_),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\mem[24][16] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(_0686_),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\mem[15][12] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\mem[30][0] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(_0650_),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\mem[26][30] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(_0091_),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\mem[11][8] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(_0197_),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\mem[13][22] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(_0499_),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\mem[13][19] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(_0496_),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\mem[30][25] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_0606_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(_0631_),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\mem[25][26] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(_0760_),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\mem[4][10] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(_0327_),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\mem[22][11] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(_0585_),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\mem[12][26] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(_0151_),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\mem[28][17] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\mem[31][0] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(_0847_),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\mem[15][8] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(_0646_),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\mem[11][31] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(_0220_),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\mem[10][26] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(_0439_),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\mem[9][6] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(_0099_),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\mem[27][23] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_0702_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(_0789_),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\mem[26][17] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(_0078_),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\mem[25][31] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(_0765_),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\mem[8][21] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(_0018_),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\mem[7][15] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(_0044_),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\mem[25][7] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\mem[21][4] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(_0741_),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\mem[1][12] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(_0297_),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\mem[20][28] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(_0409_),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\mem[18][23] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(_0244_),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\mem[18][7] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(_0228_),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\mem[3][29] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_0350_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_0545_),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(_0827_),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\mem[10][19] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(_0432_),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\mem[11][26] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(_0215_),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\mem[6][17] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(_0975_),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\mem[1][8] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(_0293_),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\mem[15][2] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\mem[23][4] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(_0640_),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\mem[22][10] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(_0584_),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\mem[9][3] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(_0096_),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\mem[5][6] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(_0515_),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\mem[20][12] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(_0393_),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\mem[1][21] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_0161_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(_0306_),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\mem[4][8] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(_0325_),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\mem[9][29] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(_0122_),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\mem[8][22] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(_0019_),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\mem[12][23] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(_0148_),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\mem[1][11] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\mem[30][1] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(_0296_),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\mem[14][8] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(_0453_),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\mem[14][12] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(_0457_),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\mem[23][15] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(_0172_),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\mem[9][16] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(_0109_),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\mem[5][17] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_0607_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(_0526_),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\mem[9][8] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(_0101_),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\mem[27][28] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(_0794_),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\mem[27][7] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(_0773_),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\mem[0][18] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(_0271_),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\mem[26][29] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\mem[19][5] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(_0090_),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\mem[6][21] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(_0979_),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\mem[22][23] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(_0597_),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\mem[25][10] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(_0744_),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\mem[9][13] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(_0106_),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\mem[4][3] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_0899_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(_0320_),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\mem[10][31] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(_0444_),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\mem[0][20] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(_0273_),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\mem[15][10] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(_0648_),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\mem[12][13] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(_0138_),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\mem[18][15] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\mem[20][1] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(_0236_),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\mem[2][15] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(_0877_),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\mem[16][3] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(_0352_),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\mem[13][11] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(_0488_),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\mem[24][7] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(_0677_),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\mem[23][22] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_0382_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(_0179_),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\mem[12][20] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(_0145_),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\mem[14][17] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(_0462_),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\mem[13][21] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(_0498_),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\mem[22][16] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(_0590_),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\mem[7][23] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\mem[3][5] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(_0052_),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\mem[23][21] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(_0178_),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\mem[28][31] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(_0861_),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\mem[0][27] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(_0280_),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\mem[20][5] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(_0386_),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\mem[24][17] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\mem[1][0] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_0803_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(_0687_),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\mem[27][12] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(_0778_),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\mem[15][21] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(_0659_),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\mem[24][28] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(_0698_),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\mem[18][16] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(_0237_),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\mem[15][25] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\mem[3][4] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(_0663_),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\mem[5][19] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(_0528_),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\mem[9][2] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(_0095_),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\mem[21][9] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(_0550_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\mem[24][22] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(_0692_),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\mem[10][18] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_0802_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(_0431_),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\mem[6][13] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(_0971_),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\mem[15][28] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(_0666_),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\mem[8][31] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(_0028_),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\mem[30][10] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(_0616_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\mem[31][27] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\mem[11][4] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(_0729_),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\mem[13][26] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(_0503_),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\mem[30][14] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(_0620_),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\mem[18][3] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(_0224_),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\mem[31][16] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(_0718_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\mem[20][29] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_0193_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(_0410_),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\mem[15][19] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(_0657_),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\mem[9][31] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(_0124_),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\mem[11][9] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(_0198_),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\mem[24][31] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(_0701_),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\mem[23][12] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\mem[28][1] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(_0169_),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\mem[8][28] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(_0025_),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\mem[7][16] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(_0045_),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\mem[15][26] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(_0664_),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\mem[12][22] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(_0147_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\mem[10][10] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_0831_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(_0423_),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\mem[21][7] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(_0548_),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\mem[30][7] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(_0613_),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\mem[5][8] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(_0517_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\mem[2][24] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(_0886_),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\mem[10][24] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\mem[29][1] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(_0437_),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\mem[16][17] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(_0366_),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\mem[20][14] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(_0395_),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\mem[16][23] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(_0372_),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\mem[17][23] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(_0949_),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\mem[16][27] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_0991_),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(_0376_),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\mem[4][20] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(_0337_),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\mem[15][6] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(_0644_),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\mem[2][11] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(_0873_),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\mem[8][2] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(_1024_),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\mem[1][25] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\mem[30][5] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(_0310_),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\mem[25][30] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(_0764_),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\mem[15][3] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(_0641_),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\mem[27][9] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(_0775_),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\mem[16][26] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(_0375_),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\mem[0][3] ),
    .X(net1368));
 sky130_fd_sc_hd__buf_2 input1 (.A(rst),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_4 input10 (.A(wb_dat_i[11]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 input11 (.A(wb_dat_i[12]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input12 (.A(wb_dat_i[13]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 input13 (.A(wb_dat_i[14]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(wb_dat_i[15]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(wb_dat_i[16]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(wb_dat_i[17]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(wb_dat_i[18]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 input18 (.A(wb_dat_i[19]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(wb_dat_i[1]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input2 (.A(wb_adr_i[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(wb_dat_i[20]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(wb_dat_i[21]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(wb_dat_i[22]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(wb_dat_i[23]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(wb_dat_i[24]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(wb_dat_i[25]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(wb_dat_i[26]),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(wb_dat_i[27]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(wb_dat_i[28]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(wb_dat_i[29]),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input3 (.A(wb_adr_i[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(wb_dat_i[2]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 input31 (.A(wb_dat_i[30]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(wb_dat_i[31]),
    .X(net32));
 sky130_fd_sc_hd__buf_2 input33 (.A(wb_dat_i[3]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(wb_dat_i[4]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(wb_dat_i[5]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 input36 (.A(wb_dat_i[6]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 input37 (.A(wb_dat_i[7]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 input38 (.A(wb_dat_i[8]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(wb_dat_i[9]),
    .X(net39));
 sky130_fd_sc_hd__buf_4 input4 (.A(wb_adr_i[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_8 input40 (.A(wb_stb_i),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(wb_we_i),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(wb_adr_i[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_8 input6 (.A(wb_adr_i[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(wb_cyc_i),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(wb_dat_i[0]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(wb_dat_i[10]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output42 (.A(net42),
    .X(wb_ack_o));
 sky130_fd_sc_hd__buf_12 output43 (.A(net87),
    .X(wb_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output44 (.A(net84),
    .X(wb_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output45 (.A(net45),
    .X(wb_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output46 (.A(net46),
    .X(wb_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output47 (.A(net47),
    .X(wb_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output48 (.A(net83),
    .X(wb_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output49 (.A(net82),
    .X(wb_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output50 (.A(net50),
    .X(wb_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output51 (.A(net51),
    .X(wb_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output52 (.A(net81),
    .X(wb_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output53 (.A(net80),
    .X(wb_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output54 (.A(net86),
    .X(wb_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output55 (.A(net55),
    .X(wb_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output56 (.A(net79),
    .X(wb_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output57 (.A(net78),
    .X(wb_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output58 (.A(net58),
    .X(wb_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output59 (.A(net59),
    .X(wb_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output60 (.A(net77),
    .X(wb_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output61 (.A(net76),
    .X(wb_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .X(wb_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output63 (.A(net75),
    .X(wb_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output64 (.A(net64),
    .X(wb_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output65 (.A(net65),
    .X(wb_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output66 (.A(net66),
    .X(wb_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output67 (.A(net67),
    .X(wb_dat_o[31]));
 sky130_fd_sc_hd__buf_12 output68 (.A(net68),
    .X(wb_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output69 (.A(net69),
    .X(wb_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output70 (.A(net70),
    .X(wb_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output71 (.A(net71),
    .X(wb_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output72 (.A(net85),
    .X(wb_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output73 (.A(net73),
    .X(wb_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output74 (.A(net74),
    .X(wb_dat_o[9]));
 sky130_fd_sc_hd__buf_2 wire75 (.A(net63),
    .X(net75));
 sky130_fd_sc_hd__buf_2 wire76 (.A(net61),
    .X(net76));
 sky130_fd_sc_hd__buf_4 wire77 (.A(net60),
    .X(net77));
 sky130_fd_sc_hd__buf_4 wire78 (.A(net57),
    .X(net78));
 sky130_fd_sc_hd__buf_2 wire79 (.A(net56),
    .X(net79));
 sky130_fd_sc_hd__buf_2 wire80 (.A(net53),
    .X(net80));
 sky130_fd_sc_hd__buf_2 wire81 (.A(net52),
    .X(net81));
 sky130_fd_sc_hd__buf_2 wire82 (.A(net49),
    .X(net82));
 sky130_fd_sc_hd__buf_2 wire83 (.A(net48),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 wire84 (.A(net44),
    .X(net84));
 sky130_fd_sc_hd__buf_2 wire85 (.A(net72),
    .X(net85));
 sky130_fd_sc_hd__buf_4 wire86 (.A(net54),
    .X(net86));
 sky130_fd_sc_hd__buf_2 wire87 (.A(net43),
    .X(net87));
endmodule

